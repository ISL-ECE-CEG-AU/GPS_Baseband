magic
tech sky130A
magscale 1 2
timestamp 1638096800
<< locali >>
rect 544761 661759 544795 666417
rect 204211 650369 204637 650403
rect 214975 650369 215401 650403
rect 229511 650369 229937 650403
rect 230489 645507 230523 646085
rect 66211 644453 66637 644487
rect 221599 644249 222117 644283
rect 193137 643263 193171 643637
rect 198013 643569 198289 643603
rect 199059 643569 199301 643603
rect 66177 643195 66211 643229
rect 66177 643161 66637 643195
rect 198013 643127 198047 643569
rect 196909 640203 196943 642821
rect 206201 642311 206235 642345
rect 206201 642277 206569 642311
rect 201359 642141 201601 642175
rect 209789 641087 209823 643161
rect 221599 642277 222117 642311
rect 193137 639591 193171 639965
rect 221565 639557 222117 639591
rect 221565 639251 221599 639557
rect 443653 639183 443687 640305
rect 193137 635783 193171 636157
rect 193137 632111 193171 632485
rect 219909 631975 219943 634661
rect 220277 631975 220311 634661
rect 193137 628507 193171 628949
rect 545773 613411 545807 617865
rect 125643 606373 126161 606407
rect 298143 310369 298385 310403
rect 36737 309791 36771 310097
rect 39129 309927 39163 310097
rect 41337 309179 41371 310097
rect 46397 309247 46431 310097
rect 48789 309315 48823 310097
rect 55965 309383 55999 310165
rect 60657 309451 60691 310233
rect 63233 309519 63267 310233
rect 70317 309587 70351 310301
rect 298293 310131 298327 310301
rect 298661 309995 298695 310505
rect 269681 309859 269715 309961
rect 296177 309723 296211 309961
rect 112453 31535 112487 33813
rect 188353 31535 188387 31637
rect 127541 30583 127575 31365
rect 127633 30991 127667 31229
rect 127633 30651 127667 30821
rect 137293 30583 137327 30957
rect 145205 30651 145239 30889
rect 166273 30787 166307 31229
rect 195897 30855 195931 30957
rect 238769 30583 238803 31433
rect 270141 30617 270601 30651
rect 269439 30549 269773 30583
rect 239505 30379 239539 30549
rect 270141 30515 270175 30617
rect 248245 30379 248279 30481
rect 283239 9333 283389 9367
rect 286885 9299 286919 9469
rect 286827 9265 286919 9299
rect 300627 8993 300961 9027
rect 268209 4267 268243 4641
rect 268301 4335 268335 4641
rect 268393 4403 268427 4709
rect 268485 4199 268519 4505
rect 268577 4335 268611 4981
rect 268669 4267 268703 5049
rect 277317 4675 277351 4913
rect 277593 4879 277627 5185
rect 277869 4539 277903 5253
rect 277961 4743 277995 5049
rect 278053 4539 278087 5117
rect 278145 4607 278179 4845
rect 278237 4607 278271 4981
rect 278329 4675 278363 5321
rect 278513 4743 278547 5389
rect 291761 5321 291945 5355
rect 291761 5015 291795 5321
rect 301421 4743 301455 4913
rect 301605 4811 301639 4981
rect 301697 4743 301731 4777
rect 301421 4709 301731 4743
rect 26249 3655 26283 3893
rect 26341 3587 26375 3961
rect 81173 3791 81207 3961
rect 64429 3519 64463 3621
rect 71605 3315 71639 3757
rect 88901 3689 89269 3723
rect 71789 3315 71823 3485
rect 71881 3111 71915 3485
rect 87521 3315 87555 3621
rect 88901 3519 88935 3689
rect 90465 3315 90499 3485
rect 87521 3281 88073 3315
rect 90407 3281 90499 3315
rect 103529 3179 103563 4165
rect 108313 3791 108347 4029
rect 108405 3995 108439 4165
rect 368857 4165 369075 4199
rect 111717 3995 111751 4097
rect 109417 3383 109451 3893
rect 111809 3791 111843 3961
rect 103989 3281 104265 3315
rect 106875 3281 107117 3315
rect 103989 3247 104023 3281
rect 113005 3247 113039 3825
rect 113097 3247 113131 4165
rect 368857 4131 368891 4165
rect 117881 4029 118157 4063
rect 117881 3995 117915 4029
rect 114569 3519 114603 3757
rect 118065 3247 118099 3825
rect 121193 3519 121227 4029
rect 127541 3791 127575 3893
rect 127449 3451 127483 3757
rect 127725 3519 127759 4029
rect 132049 3519 132083 3689
rect 127817 3451 127851 3485
rect 127449 3417 127851 3451
rect 97583 2873 97733 2907
rect 103253 2703 103287 3077
rect 103379 2873 103471 2907
rect 103437 2839 103471 2873
rect 103529 2703 103563 2873
rect 105001 2771 105035 2941
rect 178049 2839 178083 3281
rect 178141 2839 178175 3077
rect 194241 3043 194275 3281
rect 186271 2941 186513 2975
rect 194333 2907 194367 3009
rect 195161 2907 195195 3213
rect 195437 3179 195471 3213
rect 195287 3145 195471 3179
rect 196909 2907 196943 4097
rect 200129 3723 200163 3961
rect 200589 3383 200623 3621
rect 205005 3315 205039 3893
rect 320649 2771 320683 3077
rect 320741 2975 320775 3077
rect 320833 2839 320867 2941
rect 333161 2771 333195 3009
rect 344201 2839 344235 3145
rect 344661 2907 344695 3213
rect 349077 3043 349111 3281
rect 349813 3043 349847 3213
rect 349721 2975 349755 3009
rect 349905 2975 349939 3213
rect 349721 2941 349939 2975
rect 355885 2907 355919 3349
rect 368949 3247 368983 4097
rect 369041 3451 369075 4165
rect 382933 4165 383611 4199
rect 369041 3417 369351 3451
rect 369133 3043 369167 3145
rect 369225 3043 369259 3349
rect 369317 3247 369351 3417
rect 373089 3383 373123 4097
rect 382933 3995 382967 4165
rect 383577 4131 383611 4165
rect 383427 4029 383669 4063
rect 382875 3961 382967 3995
rect 369317 3213 369501 3247
rect 583401 3111 583435 6137
rect 344753 2839 344787 2873
rect 334023 2805 334173 2839
rect 344201 2805 344787 2839
rect 355735 2805 355977 2839
rect 358863 2805 359013 2839
<< viali >>
rect 544761 666417 544795 666451
rect 544761 661725 544795 661759
rect 204177 650369 204211 650403
rect 204637 650369 204671 650403
rect 214941 650369 214975 650403
rect 215401 650369 215435 650403
rect 229477 650369 229511 650403
rect 229937 650369 229971 650403
rect 230489 646085 230523 646119
rect 230489 645473 230523 645507
rect 204122 645405 204156 645439
rect 66177 644453 66211 644487
rect 66637 644453 66671 644487
rect 221565 644249 221599 644283
rect 222117 644249 222151 644283
rect 193137 643637 193171 643671
rect 66177 643229 66211 643263
rect 193137 643229 193171 643263
rect 198289 643569 198323 643603
rect 199025 643569 199059 643603
rect 199301 643569 199335 643603
rect 66637 643161 66671 643195
rect 198013 643093 198047 643127
rect 209789 643161 209823 643195
rect 196909 642821 196943 642855
rect 206201 642345 206235 642379
rect 206569 642277 206603 642311
rect 201325 642141 201359 642175
rect 201601 642141 201635 642175
rect 221565 642277 221599 642311
rect 222117 642277 222151 642311
rect 209789 641053 209823 641087
rect 196909 640169 196943 640203
rect 443653 640305 443687 640339
rect 193137 639965 193171 639999
rect 193137 639557 193171 639591
rect 222117 639557 222151 639591
rect 221565 639217 221599 639251
rect 443653 639149 443687 639183
rect 193137 636157 193171 636191
rect 193137 635749 193171 635783
rect 219909 634661 219943 634695
rect 193137 632485 193171 632519
rect 193137 632077 193171 632111
rect 219909 631941 219943 631975
rect 220277 634661 220311 634695
rect 220277 631941 220311 631975
rect 193137 628949 193171 628983
rect 193137 628473 193171 628507
rect 545773 617865 545807 617899
rect 545773 613377 545807 613411
rect 125609 606373 125643 606407
rect 126161 606373 126195 606407
rect 298661 310505 298695 310539
rect 298109 310369 298143 310403
rect 298385 310369 298419 310403
rect 70317 310301 70351 310335
rect 60657 310233 60691 310267
rect 55965 310165 55999 310199
rect 36737 310097 36771 310131
rect 39129 310097 39163 310131
rect 39129 309893 39163 309927
rect 41337 310097 41371 310131
rect 36737 309757 36771 309791
rect 46397 310097 46431 310131
rect 48789 310097 48823 310131
rect 63233 310233 63267 310267
rect 298293 310301 298327 310335
rect 298293 310097 298327 310131
rect 269681 309961 269715 309995
rect 269681 309825 269715 309859
rect 296177 309961 296211 309995
rect 298661 309961 298695 309995
rect 296177 309689 296211 309723
rect 70317 309553 70351 309587
rect 63233 309485 63267 309519
rect 60657 309417 60691 309451
rect 55965 309349 55999 309383
rect 48789 309281 48823 309315
rect 46397 309213 46431 309247
rect 41337 309145 41371 309179
rect 112453 33813 112487 33847
rect 112453 31501 112487 31535
rect 188353 31637 188387 31671
rect 188353 31501 188387 31535
rect 238769 31433 238803 31467
rect 127541 31365 127575 31399
rect 127633 31229 127667 31263
rect 166273 31229 166307 31263
rect 127633 30957 127667 30991
rect 137293 30957 137327 30991
rect 127633 30821 127667 30855
rect 127633 30617 127667 30651
rect 127541 30549 127575 30583
rect 145205 30889 145239 30923
rect 195897 30957 195931 30991
rect 195897 30821 195931 30855
rect 166273 30753 166307 30787
rect 145205 30617 145239 30651
rect 137293 30549 137327 30583
rect 270601 30617 270635 30651
rect 238769 30549 238803 30583
rect 239505 30549 239539 30583
rect 269405 30549 269439 30583
rect 269773 30549 269807 30583
rect 239505 30345 239539 30379
rect 248245 30481 248279 30515
rect 270141 30481 270175 30515
rect 248245 30345 248279 30379
rect 286885 9469 286919 9503
rect 283205 9333 283239 9367
rect 283389 9333 283423 9367
rect 286793 9265 286827 9299
rect 300593 8993 300627 9027
rect 300961 8993 300995 9027
rect 583401 6137 583435 6171
rect 278513 5389 278547 5423
rect 278329 5321 278363 5355
rect 277869 5253 277903 5287
rect 277593 5185 277627 5219
rect 268669 5049 268703 5083
rect 268577 4981 268611 5015
rect 268393 4709 268427 4743
rect 268209 4641 268243 4675
rect 268301 4641 268335 4675
rect 268393 4369 268427 4403
rect 268485 4505 268519 4539
rect 268301 4301 268335 4335
rect 268209 4233 268243 4267
rect 268577 4301 268611 4335
rect 277317 4913 277351 4947
rect 277593 4845 277627 4879
rect 277317 4641 277351 4675
rect 278053 5117 278087 5151
rect 277961 5049 277995 5083
rect 277961 4709 277995 4743
rect 277869 4505 277903 4539
rect 278237 4981 278271 5015
rect 278145 4845 278179 4879
rect 278145 4573 278179 4607
rect 291945 5321 291979 5355
rect 291761 4981 291795 5015
rect 301605 4981 301639 5015
rect 278513 4709 278547 4743
rect 301421 4913 301455 4947
rect 301605 4777 301639 4811
rect 301697 4777 301731 4811
rect 278329 4641 278363 4675
rect 278237 4573 278271 4607
rect 278053 4505 278087 4539
rect 268669 4233 268703 4267
rect 103529 4165 103563 4199
rect 26341 3961 26375 3995
rect 26249 3893 26283 3927
rect 26249 3621 26283 3655
rect 81173 3961 81207 3995
rect 71605 3757 71639 3791
rect 81173 3757 81207 3791
rect 26341 3553 26375 3587
rect 64429 3621 64463 3655
rect 64429 3485 64463 3519
rect 89269 3689 89303 3723
rect 87521 3621 87555 3655
rect 71605 3281 71639 3315
rect 71789 3485 71823 3519
rect 71789 3281 71823 3315
rect 71881 3485 71915 3519
rect 88901 3485 88935 3519
rect 90465 3485 90499 3519
rect 88073 3281 88107 3315
rect 90373 3281 90407 3315
rect 108405 4165 108439 4199
rect 108313 4029 108347 4063
rect 113097 4165 113131 4199
rect 268485 4165 268519 4199
rect 108405 3961 108439 3995
rect 111717 4097 111751 4131
rect 111717 3961 111751 3995
rect 111809 3961 111843 3995
rect 108313 3757 108347 3791
rect 109417 3893 109451 3927
rect 111809 3757 111843 3791
rect 113005 3825 113039 3859
rect 109417 3349 109451 3383
rect 104265 3281 104299 3315
rect 106841 3281 106875 3315
rect 107117 3281 107151 3315
rect 103989 3213 104023 3247
rect 113005 3213 113039 3247
rect 196909 4097 196943 4131
rect 368857 4097 368891 4131
rect 368949 4097 368983 4131
rect 118157 4029 118191 4063
rect 121193 4029 121227 4063
rect 117881 3961 117915 3995
rect 118065 3825 118099 3859
rect 114569 3757 114603 3791
rect 114569 3485 114603 3519
rect 113097 3213 113131 3247
rect 127725 4029 127759 4063
rect 127541 3893 127575 3927
rect 121193 3485 121227 3519
rect 127449 3757 127483 3791
rect 127541 3757 127575 3791
rect 132049 3689 132083 3723
rect 127725 3485 127759 3519
rect 127817 3485 127851 3519
rect 132049 3485 132083 3519
rect 118065 3213 118099 3247
rect 178049 3281 178083 3315
rect 103529 3145 103563 3179
rect 71881 3077 71915 3111
rect 103253 3077 103287 3111
rect 97549 2873 97583 2907
rect 97733 2873 97767 2907
rect 105001 2941 105035 2975
rect 103345 2873 103379 2907
rect 103437 2805 103471 2839
rect 103529 2873 103563 2907
rect 103253 2669 103287 2703
rect 194241 3281 194275 3315
rect 178049 2805 178083 2839
rect 178141 3077 178175 3111
rect 195161 3213 195195 3247
rect 194241 3009 194275 3043
rect 194333 3009 194367 3043
rect 186237 2941 186271 2975
rect 186513 2941 186547 2975
rect 194333 2873 194367 2907
rect 195437 3213 195471 3247
rect 195253 3145 195287 3179
rect 195161 2873 195195 2907
rect 200129 3961 200163 3995
rect 200129 3689 200163 3723
rect 205005 3893 205039 3927
rect 200589 3621 200623 3655
rect 200589 3349 200623 3383
rect 355885 3349 355919 3383
rect 205005 3281 205039 3315
rect 349077 3281 349111 3315
rect 344661 3213 344695 3247
rect 344201 3145 344235 3179
rect 196909 2873 196943 2907
rect 320649 3077 320683 3111
rect 178141 2805 178175 2839
rect 105001 2737 105035 2771
rect 320741 3077 320775 3111
rect 333161 3009 333195 3043
rect 320741 2941 320775 2975
rect 320833 2941 320867 2975
rect 320833 2805 320867 2839
rect 320649 2737 320683 2771
rect 349813 3213 349847 3247
rect 349077 3009 349111 3043
rect 349721 3009 349755 3043
rect 349813 3009 349847 3043
rect 349905 3213 349939 3247
rect 373089 4097 373123 4131
rect 368949 3213 368983 3247
rect 369225 3349 369259 3383
rect 369133 3145 369167 3179
rect 369133 3009 369167 3043
rect 383577 4097 383611 4131
rect 383393 4029 383427 4063
rect 383669 4029 383703 4063
rect 382841 3961 382875 3995
rect 373089 3349 373123 3383
rect 369501 3213 369535 3247
rect 583401 3077 583435 3111
rect 369225 3009 369259 3043
rect 344661 2873 344695 2907
rect 344753 2873 344787 2907
rect 355885 2873 355919 2907
rect 333989 2805 334023 2839
rect 334173 2805 334207 2839
rect 355701 2805 355735 2839
rect 355977 2805 356011 2839
rect 358829 2805 358863 2839
rect 359013 2805 359047 2839
rect 333161 2737 333195 2771
rect 103529 2669 103563 2703
<< metal1 >>
rect 166902 700952 166908 701004
rect 166960 700992 166966 701004
rect 300118 700992 300124 701004
rect 166960 700964 300124 700992
rect 166960 700952 166966 700964
rect 300118 700952 300124 700964
rect 300176 700952 300182 701004
rect 24302 700884 24308 700936
rect 24360 700924 24366 700936
rect 185118 700924 185124 700936
rect 24360 700896 185124 700924
rect 24360 700884 24366 700896
rect 185118 700884 185124 700896
rect 185176 700884 185182 700936
rect 162762 700816 162768 700868
rect 162820 700856 162826 700868
rect 332502 700856 332508 700868
rect 162820 700828 332508 700856
rect 162820 700816 162826 700828
rect 332502 700816 332508 700828
rect 332560 700816 332566 700868
rect 164142 700748 164148 700800
rect 164200 700788 164206 700800
rect 348786 700788 348792 700800
rect 164200 700760 348792 700788
rect 164200 700748 164206 700760
rect 348786 700748 348792 700760
rect 348844 700748 348850 700800
rect 40494 700680 40500 700732
rect 40552 700720 40558 700732
rect 235994 700720 236000 700732
rect 40552 700692 236000 700720
rect 40552 700680 40558 700692
rect 235994 700680 236000 700692
rect 236052 700680 236058 700732
rect 154482 700612 154488 700664
rect 154540 700652 154546 700664
rect 397454 700652 397460 700664
rect 154540 700624 397460 700652
rect 154540 700612 154546 700624
rect 397454 700612 397460 700624
rect 397512 700612 397518 700664
rect 157242 700544 157248 700596
rect 157300 700584 157306 700596
rect 413646 700584 413652 700596
rect 157300 700556 413652 700584
rect 157300 700544 157306 700556
rect 413646 700544 413652 700556
rect 413704 700544 413710 700596
rect 147582 700476 147588 700528
rect 147640 700516 147646 700528
rect 462314 700516 462320 700528
rect 147640 700488 462320 700516
rect 147640 700476 147646 700488
rect 462314 700476 462320 700488
rect 462372 700476 462378 700528
rect 105446 700408 105452 700460
rect 105504 700448 105510 700460
rect 147306 700448 147312 700460
rect 105504 700420 147312 700448
rect 105504 700408 105510 700420
rect 147306 700408 147312 700420
rect 147364 700408 147370 700460
rect 150342 700408 150348 700460
rect 150400 700448 150406 700460
rect 478506 700448 478512 700460
rect 150400 700420 478512 700448
rect 150400 700408 150406 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 147122 700380 147128 700392
rect 73028 700352 147128 700380
rect 73028 700340 73034 700352
rect 147122 700340 147128 700352
rect 147180 700340 147186 700392
rect 147214 700340 147220 700392
rect 147272 700380 147278 700392
rect 494790 700380 494796 700392
rect 147272 700352 494796 700380
rect 147272 700340 147278 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 146938 700312 146944 700324
rect 89220 700284 146944 700312
rect 89220 700272 89226 700284
rect 146938 700272 146944 700284
rect 146996 700272 147002 700324
rect 147030 700272 147036 700324
rect 147088 700312 147094 700324
rect 527174 700312 527180 700324
rect 147088 700284 527180 700312
rect 147088 700272 147094 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 172422 700204 172428 700256
rect 172480 700244 172486 700256
rect 283834 700244 283840 700256
rect 172480 700216 283840 700244
rect 172480 700204 172486 700216
rect 283834 700204 283840 700216
rect 283892 700204 283898 700256
rect 169662 700136 169668 700188
rect 169720 700176 169726 700188
rect 267642 700176 267648 700188
rect 169720 700148 267648 700176
rect 169720 700136 169726 700148
rect 267642 700136 267648 700148
rect 267700 700136 267706 700188
rect 173802 700068 173808 700120
rect 173860 700108 173866 700120
rect 235166 700108 235172 700120
rect 173860 700080 235172 700108
rect 173860 700068 173866 700080
rect 235166 700068 235172 700080
rect 235224 700068 235230 700120
rect 137830 700000 137836 700052
rect 137888 700040 137894 700052
rect 182174 700040 182180 700052
rect 137888 700012 182180 700040
rect 137888 700000 137894 700012
rect 182174 700000 182180 700012
rect 182232 700000 182238 700052
rect 179322 699932 179328 699984
rect 179380 699972 179386 699984
rect 218974 699972 218980 699984
rect 179380 699944 218980 699972
rect 179380 699932 179386 699944
rect 218974 699932 218980 699944
rect 219032 699932 219038 699984
rect 154114 699864 154120 699916
rect 154172 699904 154178 699916
rect 180058 699904 180064 699916
rect 154172 699876 180064 699904
rect 154172 699864 154178 699876
rect 180058 699864 180064 699876
rect 180116 699864 180122 699916
rect 176562 699796 176568 699848
rect 176620 699836 176626 699848
rect 202782 699836 202788 699848
rect 176620 699808 202788 699836
rect 176620 699796 176626 699808
rect 202782 699796 202788 699808
rect 202840 699796 202846 699848
rect 170306 699728 170312 699780
rect 170364 699768 170370 699780
rect 180794 699768 180800 699780
rect 170364 699740 180800 699768
rect 170364 699728 170370 699740
rect 180794 699728 180800 699740
rect 180852 699728 180858 699780
rect 251450 699660 251456 699712
rect 251508 699700 251514 699712
rect 252462 699700 252468 699712
rect 251508 699672 252468 699700
rect 251508 699660 251514 699672
rect 252462 699660 252468 699672
rect 252520 699660 252526 699712
rect 381170 699660 381176 699712
rect 381228 699700 381234 699712
rect 382182 699700 382188 699712
rect 381228 699672 382188 699700
rect 381228 699660 381234 699672
rect 382182 699660 382188 699672
rect 382240 699660 382246 699712
rect 443730 688644 443736 688696
rect 443788 688684 443794 688696
rect 463326 688684 463332 688696
rect 443788 688656 463332 688684
rect 443788 688644 443794 688656
rect 463326 688644 463332 688656
rect 463384 688644 463390 688696
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 230474 683176 230480 683188
rect 3476 683148 230480 683176
rect 3476 683136 3482 683148
rect 230474 683136 230480 683148
rect 230532 683136 230538 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 193122 670732 193128 670744
rect 3568 670704 193128 670732
rect 3568 670692 3574 670704
rect 193122 670692 193128 670704
rect 193180 670692 193186 670744
rect 252462 666476 252468 666528
rect 252520 666516 252526 666528
rect 300762 666516 300768 666528
rect 252520 666488 300768 666516
rect 252520 666476 252526 666488
rect 300762 666476 300768 666488
rect 300820 666476 300826 666528
rect 542354 666408 542360 666460
rect 542412 666448 542418 666460
rect 544749 666451 544807 666457
rect 544749 666448 544761 666451
rect 542412 666420 544761 666448
rect 542412 666408 542418 666420
rect 544749 666417 544761 666420
rect 544795 666417 544807 666451
rect 544749 666411 544807 666417
rect 542354 661716 542360 661768
rect 542412 661756 542418 661768
rect 544749 661759 544807 661765
rect 544749 661756 544761 661759
rect 542412 661728 544761 661756
rect 542412 661716 542418 661728
rect 544749 661725 544761 661728
rect 544795 661725 544807 661759
rect 544749 661719 544807 661725
rect 235994 650604 236000 650616
rect 234186 650590 236000 650604
rect 234172 650576 236000 650590
rect 196986 650360 196992 650412
rect 197044 650400 197050 650412
rect 204165 650403 204223 650409
rect 204165 650400 204177 650403
rect 197044 650372 204177 650400
rect 197044 650360 197050 650372
rect 204165 650369 204177 650372
rect 204211 650369 204223 650403
rect 204165 650363 204223 650369
rect 204625 650403 204683 650409
rect 204625 650369 204637 650403
rect 204671 650400 204683 650403
rect 214929 650403 214987 650409
rect 214929 650400 214941 650403
rect 204671 650372 214941 650400
rect 204671 650369 204683 650372
rect 204625 650363 204683 650369
rect 214929 650369 214941 650372
rect 214975 650369 214987 650403
rect 214929 650363 214987 650369
rect 215389 650403 215447 650409
rect 215389 650369 215401 650403
rect 215435 650400 215447 650403
rect 229465 650403 229523 650409
rect 229465 650400 229477 650403
rect 215435 650372 229477 650400
rect 215435 650369 215447 650372
rect 215389 650363 215447 650369
rect 229465 650369 229477 650372
rect 229511 650369 229523 650403
rect 229465 650363 229523 650369
rect 229925 650403 229983 650409
rect 229925 650369 229937 650403
rect 229971 650400 229983 650403
rect 234172 650400 234200 650576
rect 235994 650564 236000 650576
rect 236052 650564 236058 650616
rect 229971 650372 234200 650400
rect 229971 650369 229983 650372
rect 229925 650363 229983 650369
rect 4798 650020 4804 650072
rect 4856 650060 4862 650072
rect 40126 650060 40132 650072
rect 4856 650032 40132 650060
rect 4856 650020 4862 650032
rect 40126 650020 40132 650032
rect 40184 650020 40190 650072
rect 230474 646116 230480 646128
rect 230435 646088 230480 646116
rect 230474 646076 230480 646088
rect 230532 646076 230538 646128
rect 230474 645504 230480 645516
rect 230435 645476 230480 645504
rect 230474 645464 230480 645476
rect 230532 645464 230538 645516
rect 202690 645396 202696 645448
rect 202748 645436 202754 645448
rect 204110 645439 204168 645445
rect 204110 645436 204122 645439
rect 202748 645408 204122 645436
rect 202748 645396 202754 645408
rect 204110 645405 204122 645408
rect 204156 645405 204168 645439
rect 204110 645399 204168 645405
rect 443822 644784 443828 644836
rect 443880 644784 443886 644836
rect 443730 644580 443736 644632
rect 443788 644620 443794 644632
rect 443840 644620 443868 644784
rect 443788 644592 443868 644620
rect 443788 644580 443794 644592
rect 3786 644444 3792 644496
rect 3844 644484 3850 644496
rect 66165 644487 66223 644493
rect 66165 644484 66177 644487
rect 3844 644456 66177 644484
rect 3844 644444 3850 644456
rect 66165 644453 66177 644456
rect 66211 644453 66223 644487
rect 66165 644447 66223 644453
rect 66625 644487 66683 644493
rect 66625 644453 66637 644487
rect 66671 644484 66683 644487
rect 104710 644484 104716 644496
rect 66671 644456 104716 644484
rect 66671 644453 66683 644456
rect 66625 644447 66683 644453
rect 104710 644444 104716 644456
rect 104768 644444 104774 644496
rect 429194 644348 429200 644360
rect 412606 644320 429200 644348
rect 98638 644240 98644 644292
rect 98696 644280 98702 644292
rect 104250 644280 104256 644292
rect 98696 644252 104256 644280
rect 98696 644240 98702 644252
rect 104250 644240 104256 644252
rect 104308 644240 104314 644292
rect 204530 644240 204536 644292
rect 204588 644280 204594 644292
rect 221553 644283 221611 644289
rect 221553 644280 221565 644283
rect 204588 644252 221565 644280
rect 204588 644240 204594 644252
rect 221553 644249 221565 644252
rect 221599 644249 221611 644283
rect 221553 644243 221611 644249
rect 222105 644283 222163 644289
rect 222105 644249 222117 644283
rect 222151 644280 222163 644283
rect 236178 644280 236184 644292
rect 222151 644252 236184 644280
rect 222151 644249 222163 644252
rect 222105 644243 222163 644249
rect 236178 644240 236184 644252
rect 236236 644240 236242 644292
rect 240686 644240 240692 644292
rect 240744 644280 240750 644292
rect 412606 644280 412634 644320
rect 429194 644308 429200 644320
rect 429252 644308 429258 644360
rect 240744 644252 412634 644280
rect 240744 644240 240750 644252
rect 193122 643668 193128 643680
rect 193083 643640 193128 643668
rect 193122 643628 193128 643640
rect 193180 643628 193186 643680
rect 199378 643628 199384 643680
rect 199436 643668 199442 643680
rect 199562 643668 199568 643680
rect 199436 643640 199568 643668
rect 199436 643628 199442 643640
rect 199562 643628 199568 643640
rect 199620 643628 199626 643680
rect 185118 643560 185124 643612
rect 185176 643560 185182 643612
rect 196618 643560 196624 643612
rect 196676 643600 196682 643612
rect 197998 643600 198004 643612
rect 196676 643572 198004 643600
rect 196676 643560 196682 643572
rect 197998 643560 198004 643572
rect 198056 643560 198062 643612
rect 198277 643603 198335 643609
rect 198277 643569 198289 643603
rect 198323 643600 198335 643603
rect 199013 643603 199071 643609
rect 199013 643600 199025 643603
rect 198323 643572 199025 643600
rect 198323 643569 198335 643572
rect 198277 643563 198335 643569
rect 199013 643569 199025 643572
rect 199059 643569 199071 643603
rect 199013 643563 199071 643569
rect 199289 643603 199347 643609
rect 199289 643569 199301 643603
rect 199335 643600 199347 643603
rect 204530 643600 204536 643612
rect 199335 643572 204536 643600
rect 199335 643569 199347 643572
rect 199289 643563 199347 643569
rect 204530 643560 204536 643572
rect 204588 643560 204594 643612
rect 185136 643340 185164 643560
rect 185118 643288 185124 643340
rect 185176 643288 185182 643340
rect 3602 643220 3608 643272
rect 3660 643260 3666 643272
rect 66165 643263 66223 643269
rect 66165 643260 66177 643263
rect 3660 643232 66177 643260
rect 3660 643220 3666 643232
rect 66165 643229 66177 643232
rect 66211 643229 66223 643263
rect 133782 643260 133788 643272
rect 66165 643223 66223 643229
rect 93826 643232 133788 643260
rect 66625 643195 66683 643201
rect 66625 643161 66637 643195
rect 66671 643192 66683 643195
rect 93826 643192 93854 643232
rect 133782 643220 133788 643232
rect 133840 643220 133846 643272
rect 193122 643260 193128 643272
rect 193083 643232 193128 643260
rect 193122 643220 193128 643232
rect 193180 643220 193186 643272
rect 66671 643164 93854 643192
rect 66671 643161 66683 643164
rect 66625 643155 66683 643161
rect 208394 643152 208400 643204
rect 208452 643192 208458 643204
rect 209777 643195 209835 643201
rect 209777 643192 209789 643195
rect 208452 643164 209789 643192
rect 208452 643152 208458 643164
rect 209777 643161 209789 643164
rect 209823 643192 209835 643195
rect 220170 643192 220176 643204
rect 209823 643164 220176 643192
rect 209823 643161 209835 643164
rect 209777 643155 209835 643161
rect 220170 643152 220176 643164
rect 220228 643152 220234 643204
rect 192202 643084 192208 643136
rect 192260 643124 192266 643136
rect 198001 643127 198059 643133
rect 198001 643124 198013 643127
rect 192260 643096 198013 643124
rect 192260 643084 192266 643096
rect 198001 643093 198013 643096
rect 198047 643093 198059 643127
rect 198001 643087 198059 643093
rect 206554 643084 206560 643136
rect 206612 643124 206618 643136
rect 209682 643124 209688 643136
rect 206612 643096 209688 643124
rect 206612 643084 206618 643096
rect 209682 643084 209688 643096
rect 209740 643124 209746 643136
rect 220078 643124 220084 643136
rect 209740 643096 220084 643124
rect 209740 643084 209746 643096
rect 220078 643084 220084 643096
rect 220136 643084 220142 643136
rect 160002 642880 160008 642932
rect 160060 642920 160066 642932
rect 190914 642920 190920 642932
rect 160060 642892 190920 642920
rect 160060 642880 160066 642892
rect 190914 642880 190920 642892
rect 190972 642880 190978 642932
rect 196897 642855 196955 642861
rect 196897 642821 196909 642855
rect 196943 642852 196955 642855
rect 196986 642852 196992 642864
rect 196943 642824 196992 642852
rect 196943 642821 196955 642824
rect 196897 642815 196955 642821
rect 196986 642812 196992 642824
rect 197044 642812 197050 642864
rect 201770 642444 201776 642456
rect 201696 642416 201776 642444
rect 201696 642240 201724 642416
rect 201770 642404 201776 642416
rect 201828 642404 201834 642456
rect 206189 642379 206247 642385
rect 206189 642376 206201 642379
rect 201880 642348 206201 642376
rect 201770 642240 201776 642252
rect 201696 642212 201776 642240
rect 201770 642200 201776 642212
rect 201828 642200 201834 642252
rect 192202 642132 192208 642184
rect 192260 642172 192266 642184
rect 201313 642175 201371 642181
rect 201313 642172 201325 642175
rect 192260 642144 201325 642172
rect 192260 642132 192266 642144
rect 201313 642141 201325 642144
rect 201359 642141 201371 642175
rect 201313 642135 201371 642141
rect 201589 642175 201647 642181
rect 201589 642141 201601 642175
rect 201635 642172 201647 642175
rect 201880 642172 201908 642348
rect 206189 642345 206201 642348
rect 206235 642345 206247 642379
rect 206189 642339 206247 642345
rect 206557 642311 206615 642317
rect 206557 642277 206569 642311
rect 206603 642308 206615 642311
rect 221553 642311 221611 642317
rect 221553 642308 221565 642311
rect 206603 642280 221565 642308
rect 206603 642277 206615 642280
rect 206557 642271 206615 642277
rect 221553 642277 221565 642280
rect 221599 642277 221611 642311
rect 221553 642271 221611 642277
rect 222105 642311 222163 642317
rect 222105 642277 222117 642311
rect 222151 642308 222163 642311
rect 236178 642308 236184 642320
rect 222151 642280 236184 642308
rect 222151 642277 222163 642280
rect 222105 642271 222163 642277
rect 236178 642268 236184 642280
rect 236236 642268 236242 642320
rect 241606 642268 241612 642320
rect 241664 642308 241670 642320
rect 364334 642308 364340 642320
rect 241664 642280 364340 642308
rect 241664 642268 241670 642280
rect 364334 642268 364340 642280
rect 364392 642268 364398 642320
rect 201635 642144 201908 642172
rect 201635 642141 201647 642144
rect 201589 642135 201647 642141
rect 580534 641696 580540 641708
rect 475672 641668 580540 641696
rect 209777 641087 209835 641093
rect 209777 641053 209789 641087
rect 209823 641053 209835 641087
rect 209777 641047 209835 641053
rect 209792 640866 209820 641047
rect 471790 640840 471796 640892
rect 471848 640880 471854 640892
rect 475672 640880 475700 641668
rect 580534 641656 580540 641668
rect 580592 641656 580598 641708
rect 471848 640852 475700 640880
rect 471848 640840 471854 640852
rect 443641 640339 443699 640345
rect 443641 640305 443653 640339
rect 443687 640336 443699 640339
rect 459554 640336 459560 640348
rect 443687 640308 459560 640336
rect 443687 640305 443699 640308
rect 443641 640299 443699 640305
rect 459554 640296 459560 640308
rect 459612 640296 459618 640348
rect 196894 640200 196900 640212
rect 196855 640172 196900 640200
rect 196894 640160 196900 640172
rect 196952 640160 196958 640212
rect 185118 639956 185124 640008
rect 185176 639956 185182 640008
rect 193122 639996 193128 640008
rect 193083 639968 193128 639996
rect 193122 639956 193128 639968
rect 193180 639956 193186 640008
rect 185136 639736 185164 639956
rect 185118 639684 185124 639736
rect 185176 639684 185182 639736
rect 443730 639616 443736 639668
rect 443788 639616 443794 639668
rect 193122 639588 193128 639600
rect 193083 639560 193128 639588
rect 193122 639548 193128 639560
rect 193180 639548 193186 639600
rect 222105 639591 222163 639597
rect 222105 639557 222117 639591
rect 222151 639588 222163 639591
rect 224862 639588 224868 639600
rect 222151 639560 224868 639588
rect 222151 639557 222163 639560
rect 222105 639551 222163 639557
rect 224862 639548 224868 639560
rect 224920 639588 224926 639600
rect 230474 639588 230480 639600
rect 224920 639560 230480 639588
rect 224920 639548 224926 639560
rect 230474 639548 230480 639560
rect 230532 639548 230538 639600
rect 202230 639208 202236 639260
rect 202288 639248 202294 639260
rect 221553 639251 221611 639257
rect 221553 639248 221565 639251
rect 202288 639220 221565 639248
rect 202288 639208 202294 639220
rect 221553 639217 221565 639220
rect 221599 639217 221611 639251
rect 221553 639211 221611 639217
rect 443748 639192 443776 639616
rect 443638 639180 443644 639192
rect 443599 639152 443644 639180
rect 443638 639140 443644 639152
rect 443696 639140 443702 639192
rect 443730 639140 443736 639192
rect 443788 639140 443794 639192
rect 193122 636188 193128 636200
rect 193083 636160 193128 636188
rect 193122 636148 193128 636160
rect 193180 636148 193186 636200
rect 185118 636080 185124 636132
rect 185176 636080 185182 636132
rect 185136 635860 185164 636080
rect 185118 635808 185124 635860
rect 185176 635808 185182 635860
rect 193122 635780 193128 635792
rect 193083 635752 193128 635780
rect 193122 635740 193128 635752
rect 193180 635740 193186 635792
rect 219897 634695 219955 634701
rect 219897 634661 219909 634695
rect 219943 634692 219955 634695
rect 220078 634692 220084 634704
rect 219943 634664 220084 634692
rect 219943 634661 219955 634664
rect 219897 634655 219955 634661
rect 220078 634652 220084 634664
rect 220136 634652 220142 634704
rect 220262 634692 220268 634704
rect 220223 634664 220268 634692
rect 220262 634652 220268 634664
rect 220320 634652 220326 634704
rect 193122 632516 193128 632528
rect 193083 632488 193128 632516
rect 193122 632476 193128 632488
rect 193180 632476 193186 632528
rect 185118 632408 185124 632460
rect 185176 632408 185182 632460
rect 185136 632188 185164 632408
rect 185118 632136 185124 632188
rect 185176 632136 185182 632188
rect 193122 632108 193128 632120
rect 193083 632080 193128 632108
rect 193122 632068 193128 632080
rect 193180 632068 193186 632120
rect 219894 631972 219900 631984
rect 219855 631944 219900 631972
rect 219894 631932 219900 631944
rect 219952 631932 219958 631984
rect 220265 631975 220323 631981
rect 220265 631941 220277 631975
rect 220311 631972 220323 631975
rect 220354 631972 220360 631984
rect 220311 631944 220360 631972
rect 220311 631941 220323 631944
rect 220265 631935 220323 631941
rect 220354 631932 220360 631944
rect 220412 631932 220418 631984
rect 193122 628980 193128 628992
rect 193083 628952 193128 628980
rect 193122 628940 193128 628952
rect 193180 628940 193186 628992
rect 185118 628872 185124 628924
rect 185176 628872 185182 628924
rect 185136 628652 185164 628872
rect 196894 628668 196900 628720
rect 196952 628668 196958 628720
rect 185118 628600 185124 628652
rect 185176 628600 185182 628652
rect 193122 628504 193128 628516
rect 193083 628476 193128 628504
rect 193122 628464 193128 628476
rect 193180 628464 193186 628516
rect 196912 628368 196940 628668
rect 196986 628368 196992 628380
rect 196912 628340 196992 628368
rect 196986 628328 196992 628340
rect 197044 628328 197050 628380
rect 542354 617856 542360 617908
rect 542412 617896 542418 617908
rect 545761 617899 545819 617905
rect 545761 617896 545773 617899
rect 542412 617868 545773 617896
rect 542412 617856 542418 617868
rect 545761 617865 545773 617868
rect 545807 617865 545819 617899
rect 545761 617859 545819 617865
rect 382182 615476 382188 615528
rect 382240 615516 382246 615528
rect 382240 615488 452778 615516
rect 382240 615476 382246 615488
rect 542354 613368 542360 613420
rect 542412 613408 542418 613420
rect 545761 613411 545819 613417
rect 545761 613408 545773 613411
rect 542412 613380 545773 613408
rect 542412 613368 542418 613380
rect 545761 613377 545773 613380
rect 545807 613377 545819 613411
rect 545761 613371 545819 613377
rect 114462 606364 114468 606416
rect 114520 606404 114526 606416
rect 118970 606404 118976 606416
rect 114520 606376 118976 606404
rect 114520 606364 114526 606376
rect 118970 606364 118976 606376
rect 119028 606364 119034 606416
rect 119982 606364 119988 606416
rect 120040 606404 120046 606416
rect 125597 606407 125655 606413
rect 125597 606404 125609 606407
rect 120040 606376 125609 606404
rect 120040 606364 120046 606376
rect 125597 606373 125609 606376
rect 125643 606373 125655 606407
rect 125597 606367 125655 606373
rect 126149 606407 126207 606413
rect 126149 606373 126161 606407
rect 126195 606404 126207 606407
rect 211154 606404 211160 606416
rect 126195 606376 211160 606404
rect 126195 606373 126207 606376
rect 126149 606367 126207 606373
rect 211154 606364 211160 606376
rect 211212 606364 211218 606416
rect 3142 593308 3148 593360
rect 3200 593348 3206 593360
rect 40034 593348 40040 593360
rect 3200 593320 40040 593348
rect 3200 593308 3206 593320
rect 40034 593308 40040 593320
rect 40092 593308 40098 593360
rect 167454 591268 167460 591320
rect 167512 591308 167518 591320
rect 580166 591308 580172 591320
rect 167512 591280 580172 591308
rect 167512 591268 167518 591280
rect 580166 591268 580172 591280
rect 580224 591268 580230 591320
rect 167454 579640 167460 579692
rect 167512 579680 167518 579692
rect 210418 579680 210424 579692
rect 167512 579652 210424 579680
rect 167512 579640 167518 579652
rect 210418 579640 210424 579652
rect 210476 579640 210482 579692
rect 167454 577464 167460 577516
rect 167512 577504 167518 577516
rect 580166 577504 580172 577516
rect 167512 577476 580172 577504
rect 167512 577464 167518 577476
rect 580166 577464 580172 577476
rect 580224 577464 580230 577516
rect 424962 570596 424968 570648
rect 425020 570636 425026 570648
rect 443730 570636 443736 570648
rect 425020 570608 443736 570636
rect 425020 570596 425026 570608
rect 443730 570596 443736 570608
rect 443788 570596 443794 570648
rect 410334 569916 410340 569968
rect 410392 569956 410398 569968
rect 424318 569956 424324 569968
rect 410392 569928 424324 569956
rect 410392 569916 410398 569928
rect 424318 569916 424324 569928
rect 424376 569956 424382 569968
rect 424962 569956 424968 569968
rect 424376 569928 424968 569956
rect 424376 569916 424382 569928
rect 424962 569916 424968 569928
rect 425020 569916 425026 569968
rect 404262 566856 404268 566908
rect 404320 566856 404326 566908
rect 404280 566488 404308 566856
rect 427814 566488 427820 566500
rect 404280 566460 427820 566488
rect 427814 566448 427820 566460
rect 427872 566448 427878 566500
rect 92382 558900 92388 558952
rect 92440 558940 92446 558952
rect 391842 558940 391848 558952
rect 92440 558912 391848 558940
rect 92440 558900 92446 558912
rect 391842 558900 391848 558912
rect 391900 558900 391906 558952
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 218054 553432 218060 553444
rect 3384 553404 218060 553432
rect 3384 553392 3390 553404
rect 218054 553392 218060 553404
rect 218112 553392 218118 553444
rect 99282 542376 99288 542428
rect 99340 542416 99346 542428
rect 391382 542416 391388 542428
rect 99340 542388 391388 542416
rect 99340 542376 99346 542388
rect 391382 542376 391388 542388
rect 391440 542416 391446 542428
rect 391750 542416 391756 542428
rect 391440 542388 391756 542416
rect 391440 542376 391446 542388
rect 391750 542376 391756 542388
rect 391808 542376 391814 542428
rect 3326 540880 3332 540932
rect 3384 540920 3390 540932
rect 40218 540920 40224 540932
rect 3384 540892 40224 540920
rect 3384 540880 3390 540892
rect 40218 540880 40224 540892
rect 40276 540880 40282 540932
rect 111702 536800 111708 536852
rect 111760 536840 111766 536852
rect 580166 536840 580172 536852
rect 111760 536812 580172 536840
rect 111760 536800 111766 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 417694 534012 417700 534064
rect 417752 534052 417758 534064
rect 580718 534052 580724 534064
rect 417752 534024 580724 534052
rect 417752 534012 417758 534024
rect 580718 534012 580724 534024
rect 580776 534012 580782 534064
rect 401594 533944 401600 533996
rect 401652 533984 401658 533996
rect 402054 533984 402060 533996
rect 401652 533956 402060 533984
rect 401652 533944 401658 533956
rect 402054 533944 402060 533956
rect 402112 533984 402118 533996
rect 542354 533984 542360 533996
rect 402112 533956 542360 533984
rect 402112 533944 402118 533956
rect 542354 533944 542360 533956
rect 542412 533944 542418 533996
rect 143442 533400 143448 533452
rect 143500 533440 143506 533452
rect 401594 533440 401600 533452
rect 143500 533412 401600 533440
rect 143500 533400 143506 533412
rect 401594 533400 401600 533412
rect 401652 533400 401658 533452
rect 115842 533332 115848 533384
rect 115900 533372 115906 533384
rect 417694 533372 417700 533384
rect 115900 533344 417700 533372
rect 115900 533332 115906 533344
rect 417694 533332 417700 533344
rect 417752 533332 417758 533384
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 223574 527184 223580 527196
rect 3384 527156 223580 527184
rect 3384 527144 3390 527156
rect 223574 527144 223580 527156
rect 223632 527144 223638 527196
rect 114462 524424 114468 524476
rect 114520 524464 114526 524476
rect 580166 524464 580172 524476
rect 114520 524436 580172 524464
rect 114520 524424 114526 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 108942 510620 108948 510672
rect 109000 510660 109006 510672
rect 580166 510660 580172 510672
rect 109000 510632 580172 510660
rect 109000 510620 109006 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 226334 501004 226340 501016
rect 3384 500976 226340 501004
rect 3384 500964 3390 500976
rect 226334 500964 226340 500976
rect 226392 500964 226398 501016
rect 3142 489812 3148 489864
rect 3200 489852 3206 489864
rect 40126 489852 40132 489864
rect 3200 489824 40132 489852
rect 3200 489812 3206 489824
rect 40126 489812 40132 489824
rect 40184 489812 40190 489864
rect 104802 484372 104808 484424
rect 104860 484412 104866 484424
rect 579614 484412 579620 484424
rect 104860 484384 579620 484412
rect 104860 484372 104866 484384
rect 579614 484372 579620 484384
rect 579672 484372 579678 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 230474 474756 230480 474768
rect 3108 474728 230480 474756
rect 3108 474716 3114 474728
rect 230474 474716 230480 474728
rect 230532 474716 230538 474768
rect 106182 470568 106188 470620
rect 106240 470608 106246 470620
rect 579982 470608 579988 470620
rect 106240 470580 579988 470608
rect 106240 470568 106246 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 200758 462380 200764 462392
rect 3384 462352 200764 462380
rect 3384 462340 3390 462352
rect 200758 462340 200764 462352
rect 200816 462340 200822 462392
rect 424318 458124 424324 458176
rect 424376 458164 424382 458176
rect 424962 458164 424968 458176
rect 424376 458136 424968 458164
rect 424376 458124 424382 458136
rect 424962 458124 424968 458136
rect 425020 458164 425026 458176
rect 580166 458164 580172 458176
rect 425020 458136 580172 458164
rect 425020 458124 425026 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 100754 457444 100760 457496
rect 100812 457484 100818 457496
rect 424962 457484 424968 457496
rect 100812 457456 424968 457484
rect 100812 457444 100818 457456
rect 424962 457444 424968 457456
rect 425020 457444 425026 457496
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 233234 448576 233240 448588
rect 3384 448548 233240 448576
rect 3384 448536 3390 448548
rect 233234 448536 233240 448548
rect 233292 448536 233298 448588
rect 3326 437384 3332 437436
rect 3384 437424 3390 437436
rect 40034 437424 40040 437436
rect 3384 437396 40040 437424
rect 3384 437384 3390 437396
rect 40034 437384 40040 437396
rect 40092 437384 40098 437436
rect 96522 430584 96528 430636
rect 96580 430624 96586 430636
rect 580166 430624 580172 430636
rect 96580 430596 580172 430624
rect 96580 430584 96586 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3142 422288 3148 422340
rect 3200 422328 3206 422340
rect 237374 422328 237380 422340
rect 3200 422300 237380 422328
rect 3200 422288 3206 422300
rect 237374 422288 237380 422300
rect 237432 422288 237438 422340
rect 391750 419432 391756 419484
rect 391808 419472 391814 419484
rect 579614 419472 579620 419484
rect 391808 419444 579620 419472
rect 391808 419432 391814 419444
rect 579614 419432 579620 419444
rect 579672 419432 579678 419484
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 217318 409884 217324 409896
rect 3384 409856 217324 409884
rect 3384 409844 3390 409856
rect 217318 409844 217324 409856
rect 217376 409844 217382 409896
rect 95142 404336 95148 404388
rect 95200 404376 95206 404388
rect 580166 404376 580172 404388
rect 95200 404348 580172 404376
rect 95200 404336 95206 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 240134 397508 240140 397520
rect 3384 397480 240140 397508
rect 3384 397468 3390 397480
rect 240134 397468 240140 397480
rect 240192 397468 240198 397520
rect 89622 378156 89628 378208
rect 89680 378196 89686 378208
rect 579614 378196 579620 378208
rect 89680 378168 579620 378196
rect 89680 378156 89686 378168
rect 579614 378156 579620 378168
rect 579672 378156 579678 378208
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 245654 371260 245660 371272
rect 3384 371232 245660 371260
rect 3384 371220 3390 371232
rect 245654 371220 245660 371232
rect 245712 371220 245718 371272
rect 391842 365644 391848 365696
rect 391900 365684 391906 365696
rect 580166 365684 580172 365696
rect 391900 365656 580172 365684
rect 391900 365644 391906 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 88242 351908 88248 351960
rect 88300 351948 88306 351960
rect 580166 351948 580172 351960
rect 88300 351920 580172 351948
rect 88300 351908 88306 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 247034 345080 247040 345092
rect 3384 345052 247040 345080
rect 3384 345040 3390 345052
rect 247034 345040 247040 345052
rect 247092 345040 247098 345092
rect 82538 324300 82544 324352
rect 82596 324340 82602 324352
rect 579982 324340 579988 324352
rect 82596 324312 579988 324340
rect 82596 324300 82602 324312
rect 579982 324300 579988 324312
rect 580040 324300 580046 324352
rect 3602 318792 3608 318844
rect 3660 318832 3666 318844
rect 252738 318832 252744 318844
rect 3660 318804 252744 318832
rect 3660 318792 3666 318804
rect 252738 318792 252744 318804
rect 252796 318792 252802 318844
rect 147122 314576 147128 314628
rect 147180 314616 147186 314628
rect 190454 314616 190460 314628
rect 147180 314588 190460 314616
rect 147180 314576 147186 314588
rect 190454 314576 190460 314588
rect 190512 314576 190518 314628
rect 8202 314508 8208 314560
rect 8260 314548 8266 314560
rect 197446 314548 197452 314560
rect 8260 314520 197452 314548
rect 8260 314508 8266 314520
rect 197446 314508 197452 314520
rect 197504 314508 197510 314560
rect 3418 314440 3424 314492
rect 3476 314480 3482 314492
rect 204622 314480 204628 314492
rect 3476 314452 204628 314480
rect 3476 314440 3482 314452
rect 204622 314440 204628 314452
rect 204680 314440 204686 314492
rect 3510 314372 3516 314424
rect 3568 314412 3574 314424
rect 209774 314412 209780 314424
rect 3568 314384 209780 314412
rect 3568 314372 3574 314384
rect 209774 314372 209780 314384
rect 209832 314372 209838 314424
rect 135070 314304 135076 314356
rect 135128 314344 135134 314356
rect 443638 314344 443644 314356
rect 135128 314316 443644 314344
rect 135128 314304 135134 314316
rect 443638 314304 443644 314316
rect 443696 314304 443702 314356
rect 137830 314236 137836 314288
rect 137888 314276 137894 314288
rect 558914 314276 558920 314288
rect 137888 314248 558920 314276
rect 137888 314236 137894 314248
rect 558914 314236 558920 314248
rect 558972 314236 558978 314288
rect 133046 314168 133052 314220
rect 133104 314208 133110 314220
rect 580258 314208 580264 314220
rect 133104 314180 580264 314208
rect 133104 314168 133110 314180
rect 580258 314168 580264 314180
rect 580316 314168 580322 314220
rect 130654 314100 130660 314152
rect 130712 314140 130718 314152
rect 580350 314140 580356 314152
rect 130712 314112 580356 314140
rect 130712 314100 130718 314112
rect 580350 314100 580356 314112
rect 580408 314100 580414 314152
rect 128262 314032 128268 314084
rect 128320 314072 128326 314084
rect 580534 314072 580540 314084
rect 128320 314044 580540 314072
rect 128320 314032 128326 314044
rect 580534 314032 580540 314044
rect 580592 314032 580598 314084
rect 125502 313964 125508 314016
rect 125560 314004 125566 314016
rect 580442 314004 580448 314016
rect 125560 313976 580448 314004
rect 125560 313964 125566 313976
rect 580442 313964 580448 313976
rect 580500 313964 580506 314016
rect 123386 313896 123392 313948
rect 123444 313936 123450 313948
rect 580626 313936 580632 313948
rect 123444 313908 580632 313936
rect 123444 313896 123450 313908
rect 580626 313896 580632 313908
rect 580684 313896 580690 313948
rect 147306 313828 147312 313880
rect 147364 313868 147370 313880
rect 187786 313868 187792 313880
rect 147364 313840 187792 313868
rect 147364 313828 147370 313840
rect 187786 313828 187792 313840
rect 187844 313828 187850 313880
rect 220078 313352 220084 313404
rect 220136 313392 220142 313404
rect 228726 313392 228732 313404
rect 220136 313364 228732 313392
rect 220136 313352 220142 313364
rect 228726 313352 228732 313364
rect 228784 313352 228790 313404
rect 144730 313284 144736 313336
rect 144788 313324 144794 313336
rect 147214 313324 147220 313336
rect 144788 313296 147220 313324
rect 144788 313284 144794 313296
rect 147214 313284 147220 313296
rect 147272 313284 147278 313336
rect 195698 313284 195704 313336
rect 195756 313324 195762 313336
rect 196986 313324 196992 313336
rect 195756 313296 196992 313324
rect 195756 313284 195762 313296
rect 196986 313284 196992 313296
rect 197044 313284 197050 313336
rect 220170 313284 220176 313336
rect 220228 313324 220234 313336
rect 221550 313324 221556 313336
rect 220228 313296 221556 313324
rect 220228 313284 220234 313296
rect 221550 313284 221556 313296
rect 221608 313284 221614 313336
rect 185118 313216 185124 313268
rect 185176 313256 185182 313268
rect 185670 313256 185676 313268
rect 185176 313228 185676 313256
rect 185176 313216 185182 313228
rect 185670 313216 185676 313228
rect 185728 313216 185734 313268
rect 146938 313148 146944 313200
rect 146996 313188 147002 313200
rect 192570 313188 192576 313200
rect 146996 313160 151814 313188
rect 146996 313148 147002 313160
rect 140314 313080 140320 313132
rect 140372 313120 140378 313132
rect 147030 313120 147036 313132
rect 140372 313092 147036 313120
rect 140372 313080 140378 313092
rect 147030 313080 147036 313092
rect 147088 313080 147094 313132
rect 87322 313012 87328 313064
rect 87380 313052 87386 313064
rect 88242 313052 88248 313064
rect 87380 313024 88248 313052
rect 87380 313012 87386 313024
rect 88242 313012 88248 313024
rect 88300 313012 88306 313064
rect 94498 313012 94504 313064
rect 94556 313052 94562 313064
rect 95142 313052 95148 313064
rect 94556 313024 95148 313052
rect 94556 313012 94562 313024
rect 95142 313012 95148 313024
rect 95200 313012 95206 313064
rect 104158 313012 104164 313064
rect 104216 313052 104222 313064
rect 104802 313052 104808 313064
rect 104216 313024 104808 313052
rect 104216 313012 104222 313024
rect 104802 313012 104808 313024
rect 104860 313012 104866 313064
rect 113818 313012 113824 313064
rect 113876 313052 113882 313064
rect 114462 313052 114468 313064
rect 113876 313024 114468 313052
rect 113876 313012 113882 313024
rect 114462 313012 114468 313024
rect 114520 313012 114526 313064
rect 142706 313012 142712 313064
rect 142764 313052 142770 313064
rect 143442 313052 143448 313064
rect 142764 313024 143448 313052
rect 142764 313012 142770 313024
rect 143442 313012 143448 313024
rect 143500 313012 143506 313064
rect 149882 313012 149888 313064
rect 149940 313052 149946 313064
rect 150342 313052 150348 313064
rect 149940 313024 150348 313052
rect 149940 313012 149946 313024
rect 150342 313012 150348 313024
rect 150400 313012 150406 313064
rect 151786 313052 151814 313160
rect 185596 313160 192576 313188
rect 152274 313080 152280 313132
rect 152332 313120 152338 313132
rect 153102 313120 153108 313132
rect 152332 313092 153108 313120
rect 152332 313080 152338 313092
rect 153102 313080 153108 313092
rect 153160 313080 153166 313132
rect 159542 313080 159548 313132
rect 159600 313120 159606 313132
rect 160002 313120 160008 313132
rect 159600 313092 160008 313120
rect 159600 313080 159606 313092
rect 160002 313080 160008 313092
rect 160060 313080 160066 313132
rect 161934 313080 161940 313132
rect 161992 313120 161998 313132
rect 162762 313120 162768 313132
rect 161992 313092 162768 313120
rect 161992 313080 161998 313092
rect 162762 313080 162768 313092
rect 162820 313080 162826 313132
rect 169202 313080 169208 313132
rect 169260 313120 169266 313132
rect 169662 313120 169668 313132
rect 169260 313092 169668 313120
rect 169260 313080 169266 313092
rect 169662 313080 169668 313092
rect 169720 313080 169726 313132
rect 171594 313080 171600 313132
rect 171652 313120 171658 313132
rect 172422 313120 172428 313132
rect 171652 313092 172428 313120
rect 171652 313080 171658 313092
rect 172422 313080 172428 313092
rect 172480 313080 172486 313132
rect 178770 313080 178776 313132
rect 178828 313120 178834 313132
rect 179322 313120 179328 313132
rect 178828 313092 179328 313120
rect 178828 313080 178834 313092
rect 179322 313080 179328 313092
rect 179380 313080 179386 313132
rect 180058 313080 180064 313132
rect 180116 313120 180122 313132
rect 185394 313120 185400 313132
rect 180116 313092 185400 313120
rect 180116 313080 180122 313092
rect 185394 313080 185400 313092
rect 185452 313080 185458 313132
rect 185596 313052 185624 313160
rect 192570 313148 192576 313160
rect 192628 313148 192634 313200
rect 193122 313148 193128 313200
rect 193180 313188 193186 313200
rect 193180 313160 201724 313188
rect 193180 313148 193186 313160
rect 185670 313080 185676 313132
rect 185728 313120 185734 313132
rect 200114 313120 200120 313132
rect 185728 313092 200120 313120
rect 185728 313080 185734 313092
rect 200114 313080 200120 313092
rect 200172 313080 200178 313132
rect 201696 313120 201724 313160
rect 201770 313148 201776 313200
rect 201828 313188 201834 313200
rect 214282 313188 214288 313200
rect 201828 313160 214288 313188
rect 201828 313148 201834 313160
rect 214282 313148 214288 313160
rect 214340 313148 214346 313200
rect 207014 313120 207020 313132
rect 201696 313092 207020 313120
rect 207014 313080 207020 313092
rect 207072 313080 207078 313132
rect 210418 313080 210424 313132
rect 210476 313120 210482 313132
rect 216674 313120 216680 313132
rect 210476 313092 216680 313120
rect 210476 313080 210482 313092
rect 216674 313080 216680 313092
rect 216732 313080 216738 313132
rect 217318 313080 217324 313132
rect 217376 313120 217382 313132
rect 243170 313120 243176 313132
rect 217376 313092 243176 313120
rect 217376 313080 217382 313092
rect 243170 313080 243176 313092
rect 243228 313080 243234 313132
rect 151786 313024 185624 313052
rect 200758 313012 200764 313064
rect 200816 313052 200822 313064
rect 235994 313052 236000 313064
rect 200816 313024 236000 313052
rect 200816 313012 200822 313024
rect 235994 313012 236000 313024
rect 236052 313012 236058 313064
rect 77662 312944 77668 312996
rect 77720 312984 77726 312996
rect 304626 312984 304632 312996
rect 77720 312956 304632 312984
rect 77720 312944 77726 312956
rect 304626 312944 304632 312956
rect 304684 312944 304690 312996
rect 3878 312876 3884 312928
rect 3936 312916 3942 312928
rect 250438 312916 250444 312928
rect 3936 312888 250444 312916
rect 3936 312876 3942 312888
rect 250438 312876 250444 312888
rect 250496 312876 250502 312928
rect 6362 312808 6368 312860
rect 6420 312848 6426 312860
rect 257614 312848 257620 312860
rect 6420 312820 257620 312848
rect 6420 312808 6426 312820
rect 257614 312808 257620 312820
rect 257672 312808 257678 312860
rect 5442 312740 5448 312792
rect 5500 312780 5506 312792
rect 260006 312780 260012 312792
rect 5500 312752 260012 312780
rect 5500 312740 5506 312752
rect 260006 312740 260012 312752
rect 260064 312740 260070 312792
rect 5350 312672 5356 312724
rect 5408 312712 5414 312724
rect 267274 312712 267280 312724
rect 5408 312684 267280 312712
rect 5408 312672 5414 312684
rect 267274 312672 267280 312684
rect 267332 312672 267338 312724
rect 3326 312604 3332 312656
rect 3384 312644 3390 312656
rect 264974 312644 264980 312656
rect 3384 312616 264980 312644
rect 3384 312604 3390 312616
rect 264974 312604 264980 312616
rect 265032 312604 265038 312656
rect 3970 312536 3976 312588
rect 4028 312576 4034 312588
rect 272058 312576 272064 312588
rect 4028 312548 272064 312576
rect 4028 312536 4034 312548
rect 272058 312536 272064 312548
rect 272116 312536 272122 312588
rect 5258 312468 5264 312520
rect 5316 312508 5322 312520
rect 274634 312508 274640 312520
rect 5316 312480 274640 312508
rect 5316 312468 5322 312480
rect 274634 312468 274640 312480
rect 274692 312468 274698 312520
rect 3694 312400 3700 312452
rect 3752 312440 3758 312452
rect 276934 312440 276940 312452
rect 3752 312412 276940 312440
rect 3752 312400 3758 312412
rect 276934 312400 276940 312412
rect 276992 312400 276998 312452
rect 3786 312332 3792 312384
rect 3844 312372 3850 312384
rect 279326 312372 279332 312384
rect 3844 312344 279332 312372
rect 3844 312332 3850 312344
rect 279326 312332 279332 312344
rect 279384 312332 279390 312384
rect 5166 312264 5172 312316
rect 5224 312304 5230 312316
rect 281718 312304 281724 312316
rect 5224 312276 281724 312304
rect 5224 312264 5230 312276
rect 281718 312264 281724 312276
rect 281776 312264 281782 312316
rect 5074 312196 5080 312248
rect 5132 312236 5138 312248
rect 284294 312236 284300 312248
rect 5132 312208 284300 312236
rect 5132 312196 5138 312208
rect 284294 312196 284300 312208
rect 284352 312196 284358 312248
rect 6270 312128 6276 312180
rect 6328 312168 6334 312180
rect 286502 312168 286508 312180
rect 6328 312140 286508 312168
rect 6328 312128 6334 312140
rect 286502 312128 286508 312140
rect 286560 312128 286566 312180
rect 4982 312060 4988 312112
rect 5040 312100 5046 312112
rect 288894 312100 288900 312112
rect 5040 312072 288900 312100
rect 5040 312060 5046 312072
rect 288894 312060 288900 312072
rect 288952 312060 288958 312112
rect 6178 311992 6184 312044
rect 6236 312032 6242 312044
rect 291378 312032 291384 312044
rect 6236 312004 291384 312032
rect 6236 311992 6242 312004
rect 291378 311992 291384 312004
rect 291436 311992 291442 312044
rect 3602 311924 3608 311976
rect 3660 311964 3666 311976
rect 293954 311964 293960 311976
rect 3660 311936 293960 311964
rect 3660 311924 3666 311936
rect 293954 311924 293960 311936
rect 294012 311924 294018 311976
rect 84930 311856 84936 311908
rect 84988 311896 84994 311908
rect 580166 311896 580172 311908
rect 84988 311868 580172 311896
rect 84988 311856 84994 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 298649 310539 298707 310545
rect 298649 310536 298661 310539
rect 298112 310508 298661 310536
rect 79962 310428 79968 310480
rect 80020 310468 80026 310480
rect 298112 310468 298140 310508
rect 298649 310505 298661 310508
rect 298695 310505 298707 310539
rect 298649 310499 298707 310505
rect 304534 310468 304540 310480
rect 80020 310440 298140 310468
rect 298204 310440 304540 310468
rect 80020 310428 80026 310440
rect 75270 310360 75276 310412
rect 75328 310400 75334 310412
rect 298097 310403 298155 310409
rect 298097 310400 298109 310403
rect 75328 310372 298109 310400
rect 75328 310360 75334 310372
rect 298097 310369 298109 310372
rect 298143 310369 298155 310403
rect 298097 310363 298155 310369
rect 70302 310332 70308 310344
rect 70263 310304 70308 310332
rect 70302 310292 70308 310304
rect 70360 310292 70366 310344
rect 72878 310292 72884 310344
rect 72936 310332 72942 310344
rect 298204 310332 298232 310440
rect 304534 310428 304540 310440
rect 304592 310428 304598 310480
rect 298373 310403 298431 310409
rect 298373 310369 298385 310403
rect 298419 310400 298431 310403
rect 303522 310400 303528 310412
rect 298419 310372 303528 310400
rect 298419 310369 298431 310372
rect 298373 310363 298431 310369
rect 303522 310360 303528 310372
rect 303580 310360 303586 310412
rect 72936 310304 298232 310332
rect 298281 310335 298339 310341
rect 72936 310292 72942 310304
rect 298281 310301 298293 310335
rect 298327 310332 298339 310335
rect 304350 310332 304356 310344
rect 298327 310304 304356 310332
rect 298327 310301 298339 310304
rect 298281 310295 298339 310301
rect 304350 310292 304356 310304
rect 304408 310292 304414 310344
rect 60642 310264 60648 310276
rect 60603 310236 60648 310264
rect 60642 310224 60648 310236
rect 60700 310224 60706 310276
rect 63218 310264 63224 310276
rect 63179 310236 63224 310264
rect 63218 310224 63224 310236
rect 63276 310224 63282 310276
rect 65610 310224 65616 310276
rect 65668 310264 65674 310276
rect 303430 310264 303436 310276
rect 65668 310236 303436 310264
rect 65668 310224 65674 310236
rect 303430 310224 303436 310236
rect 303488 310224 303494 310276
rect 55950 310196 55956 310208
rect 55911 310168 55956 310196
rect 55950 310156 55956 310168
rect 56008 310156 56014 310208
rect 58434 310156 58440 310208
rect 58492 310196 58498 310208
rect 303246 310196 303252 310208
rect 58492 310168 303252 310196
rect 58492 310156 58498 310168
rect 303246 310156 303252 310168
rect 303304 310156 303310 310208
rect 36722 310128 36728 310140
rect 36683 310100 36728 310128
rect 36722 310088 36728 310100
rect 36780 310088 36786 310140
rect 39114 310128 39120 310140
rect 39075 310100 39120 310128
rect 39114 310088 39120 310100
rect 39172 310088 39178 310140
rect 41322 310128 41328 310140
rect 41283 310100 41328 310128
rect 41322 310088 41328 310100
rect 41380 310088 41386 310140
rect 46382 310128 46388 310140
rect 46343 310100 46388 310128
rect 46382 310088 46388 310100
rect 46440 310088 46446 310140
rect 48774 310128 48780 310140
rect 48735 310100 48780 310128
rect 48774 310088 48780 310100
rect 48832 310088 48838 310140
rect 53558 310088 53564 310140
rect 53616 310128 53622 310140
rect 298281 310131 298339 310137
rect 298281 310128 298293 310131
rect 53616 310100 298293 310128
rect 53616 310088 53622 310100
rect 298281 310097 298293 310100
rect 298327 310097 298339 310131
rect 304258 310128 304264 310140
rect 298281 310091 298339 310097
rect 298388 310100 304264 310128
rect 4706 310020 4712 310072
rect 4764 310060 4770 310072
rect 255314 310060 255320 310072
rect 4764 310032 255320 310060
rect 4764 310020 4770 310032
rect 255314 310020 255320 310032
rect 255372 310020 255378 310072
rect 4062 309952 4068 310004
rect 4120 309992 4126 310004
rect 262490 309992 262496 310004
rect 4120 309964 262496 309992
rect 4120 309952 4126 309964
rect 262490 309952 262496 309964
rect 262548 309952 262554 310004
rect 269666 309992 269672 310004
rect 269627 309964 269672 309992
rect 269666 309952 269672 309964
rect 269724 309952 269730 310004
rect 296162 309992 296168 310004
rect 296123 309964 296168 309992
rect 296162 309952 296168 309964
rect 296220 309952 296226 310004
rect 39117 309927 39175 309933
rect 39117 309893 39129 309927
rect 39163 309924 39175 309927
rect 298388 309924 298416 310100
rect 304258 310088 304264 310100
rect 304316 310088 304322 310140
rect 303062 310060 303068 310072
rect 39163 309896 298416 309924
rect 298480 310032 303068 310060
rect 39163 309893 39175 309896
rect 39117 309887 39175 309893
rect 3878 309816 3884 309868
rect 3936 309856 3942 309868
rect 269669 309859 269727 309865
rect 269669 309856 269681 309859
rect 3936 309828 269681 309856
rect 3936 309816 3942 309828
rect 269669 309825 269681 309828
rect 269715 309825 269727 309859
rect 269669 309819 269727 309825
rect 36725 309791 36783 309797
rect 36725 309757 36737 309791
rect 36771 309788 36783 309791
rect 298480 309788 298508 310032
rect 303062 310020 303068 310032
rect 303120 310020 303126 310072
rect 298554 309952 298560 310004
rect 298612 309952 298618 310004
rect 298649 309995 298707 310001
rect 298649 309961 298661 309995
rect 298695 309992 298707 309995
rect 304718 309992 304724 310004
rect 298695 309964 304724 309992
rect 298695 309961 298707 309964
rect 298649 309955 298707 309961
rect 304718 309952 304724 309964
rect 304776 309952 304782 310004
rect 36771 309760 298508 309788
rect 36771 309757 36783 309760
rect 36725 309751 36783 309757
rect 4890 309680 4896 309732
rect 4948 309720 4954 309732
rect 296165 309723 296223 309729
rect 296165 309720 296177 309723
rect 4948 309692 296177 309720
rect 4948 309680 4954 309692
rect 296165 309689 296177 309692
rect 296211 309689 296223 309723
rect 296165 309683 296223 309689
rect 3418 309612 3424 309664
rect 3476 309652 3482 309664
rect 298572 309652 298600 309952
rect 3476 309624 298600 309652
rect 3476 309612 3482 309624
rect 70305 309587 70363 309593
rect 70305 309553 70317 309587
rect 70351 309584 70363 309587
rect 580810 309584 580816 309596
rect 70351 309556 580816 309584
rect 70351 309553 70363 309556
rect 70305 309547 70363 309553
rect 580810 309544 580816 309556
rect 580868 309544 580874 309596
rect 63221 309519 63279 309525
rect 63221 309485 63233 309519
rect 63267 309516 63279 309519
rect 580626 309516 580632 309528
rect 63267 309488 580632 309516
rect 63267 309485 63279 309488
rect 63221 309479 63279 309485
rect 580626 309476 580632 309488
rect 580684 309476 580690 309528
rect 60645 309451 60703 309457
rect 60645 309417 60657 309451
rect 60691 309448 60703 309451
rect 580718 309448 580724 309460
rect 60691 309420 580724 309448
rect 60691 309417 60703 309420
rect 60645 309411 60703 309417
rect 580718 309408 580724 309420
rect 580776 309408 580782 309460
rect 55953 309383 56011 309389
rect 55953 309349 55965 309383
rect 55999 309380 56011 309383
rect 580534 309380 580540 309392
rect 55999 309352 580540 309380
rect 55999 309349 56011 309352
rect 55953 309343 56011 309349
rect 580534 309340 580540 309352
rect 580592 309340 580598 309392
rect 48777 309315 48835 309321
rect 48777 309281 48789 309315
rect 48823 309312 48835 309315
rect 580350 309312 580356 309324
rect 48823 309284 580356 309312
rect 48823 309281 48835 309284
rect 48777 309275 48835 309281
rect 580350 309272 580356 309284
rect 580408 309272 580414 309324
rect 46385 309247 46443 309253
rect 46385 309213 46397 309247
rect 46431 309244 46443 309247
rect 580442 309244 580448 309256
rect 46431 309216 580448 309244
rect 46431 309213 46443 309216
rect 46385 309207 46443 309213
rect 580442 309204 580448 309216
rect 580500 309204 580506 309256
rect 41325 309179 41383 309185
rect 41325 309145 41337 309179
rect 41371 309176 41383 309179
rect 580258 309176 580264 309188
rect 41371 309148 580264 309176
rect 41371 309145 41383 309148
rect 41325 309139 41383 309145
rect 580258 309136 580264 309148
rect 580316 309136 580322 309188
rect 2958 306212 2964 306264
rect 3016 306252 3022 306264
rect 6362 306252 6368 306264
rect 3016 306224 6368 306252
rect 3016 306212 3022 306224
rect 6362 306212 6368 306224
rect 6420 306212 6426 306264
rect 304718 299412 304724 299464
rect 304776 299452 304782 299464
rect 580166 299452 580172 299464
rect 304776 299424 580172 299452
rect 304776 299412 304782 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 2774 293224 2780 293276
rect 2832 293264 2838 293276
rect 4706 293264 4712 293276
rect 2832 293236 4712 293264
rect 2832 293224 2838 293236
rect 4706 293224 4712 293236
rect 4764 293224 4770 293276
rect 303522 273164 303528 273216
rect 303580 273204 303586 273216
rect 579982 273204 579988 273216
rect 303580 273176 579988 273204
rect 303580 273164 303586 273176
rect 579982 273164 579988 273176
rect 580040 273164 580046 273216
rect 2774 267180 2780 267232
rect 2832 267220 2838 267232
rect 5442 267220 5448 267232
rect 2832 267192 5448 267220
rect 2832 267180 2838 267192
rect 5442 267180 5448 267192
rect 5500 267180 5506 267232
rect 304626 259360 304632 259412
rect 304684 259400 304690 259412
rect 579798 259400 579804 259412
rect 304684 259372 579804 259400
rect 304684 259360 304690 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 304534 245556 304540 245608
rect 304592 245596 304598 245608
rect 580166 245596 580172 245608
rect 304592 245568 580172 245596
rect 304592 245556 304598 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 304442 233180 304448 233232
rect 304500 233220 304506 233232
rect 579982 233220 579988 233232
rect 304500 233192 579988 233220
rect 304500 233180 304506 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 2774 214956 2780 215008
rect 2832 214996 2838 215008
rect 5350 214996 5356 215008
rect 2832 214968 5356 214996
rect 2832 214956 2838 214968
rect 5350 214956 5356 214968
rect 5408 214956 5414 215008
rect 303430 206932 303436 206984
rect 303488 206972 303494 206984
rect 579614 206972 579620 206984
rect 303488 206944 579620 206972
rect 303488 206932 303494 206944
rect 579614 206932 579620 206944
rect 579672 206932 579678 206984
rect 303246 166948 303252 167000
rect 303304 166988 303310 167000
rect 580166 166988 580172 167000
rect 303304 166960 580172 166988
rect 303304 166948 303310 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 2774 163344 2780 163396
rect 2832 163384 2838 163396
rect 5258 163384 5264 163396
rect 2832 163356 5264 163384
rect 2832 163344 2838 163356
rect 5258 163344 5264 163356
rect 5316 163344 5322 163396
rect 304350 153144 304356 153196
rect 304408 153184 304414 153196
rect 580166 153184 580172 153196
rect 304408 153156 580172 153184
rect 304408 153144 304414 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 303338 126896 303344 126948
rect 303396 126936 303402 126948
rect 579614 126936 579620 126948
rect 303396 126908 579620 126936
rect 303396 126896 303402 126908
rect 579614 126896 579620 126908
rect 579672 126896 579678 126948
rect 2774 123836 2780 123888
rect 2832 123876 2838 123888
rect 4798 123876 4804 123888
rect 2832 123848 4804 123876
rect 2832 123836 2838 123848
rect 4798 123836 4804 123848
rect 4856 123836 4862 123888
rect 2774 110712 2780 110764
rect 2832 110752 2838 110764
rect 5166 110752 5172 110764
rect 2832 110724 5172 110752
rect 2832 110712 2838 110724
rect 5166 110712 5172 110724
rect 5224 110712 5230 110764
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 6270 97764 6276 97776
rect 2832 97736 6276 97764
rect 2832 97724 2838 97736
rect 6270 97724 6276 97736
rect 6328 97724 6334 97776
rect 303154 86912 303160 86964
rect 303212 86952 303218 86964
rect 580166 86952 580172 86964
rect 303212 86924 580172 86952
rect 303212 86912 303218 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 2774 85144 2780 85196
rect 2832 85184 2838 85196
rect 5074 85184 5080 85196
rect 2832 85156 5080 85184
rect 2832 85144 2838 85156
rect 5074 85144 5080 85156
rect 5132 85144 5138 85196
rect 304258 73108 304264 73160
rect 304316 73148 304322 73160
rect 579982 73148 579988 73160
rect 304316 73120 579988 73148
rect 304316 73108 304322 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 2774 71612 2780 71664
rect 2832 71652 2838 71664
rect 4982 71652 4988 71664
rect 2832 71624 4988 71652
rect 2832 71612 2838 71624
rect 4982 71612 4988 71624
rect 5040 71612 5046 71664
rect 303062 46860 303068 46912
rect 303120 46900 303126 46912
rect 580166 46900 580172 46912
rect 303120 46872 580172 46900
rect 303120 46860 303126 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3142 45500 3148 45552
rect 3200 45540 3206 45552
rect 6178 45540 6184 45552
rect 3200 45512 6184 45540
rect 3200 45500 3206 45512
rect 6178 45500 6184 45512
rect 6236 45500 6242 45552
rect 107332 33804 107338 33856
rect 107390 33844 107396 33856
rect 112441 33847 112499 33853
rect 112441 33844 112453 33847
rect 107390 33816 112453 33844
rect 107390 33804 107396 33816
rect 112441 33813 112453 33816
rect 112487 33813 112499 33847
rect 112441 33807 112499 33813
rect 302970 33056 302976 33108
rect 303028 33096 303034 33108
rect 580166 33096 580172 33108
rect 303028 33068 580172 33096
rect 303028 33056 303034 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 2774 32852 2780 32904
rect 2832 32892 2838 32904
rect 4890 32892 4896 32904
rect 2832 32864 4896 32892
rect 2832 32852 2838 32864
rect 4890 32852 4896 32864
rect 4948 32852 4954 32904
rect 250806 31764 250812 31816
rect 250864 31804 250870 31816
rect 251082 31804 251088 31816
rect 250864 31776 251088 31804
rect 250864 31764 250870 31776
rect 251082 31764 251088 31776
rect 251140 31764 251146 31816
rect 261938 31764 261944 31816
rect 261996 31804 262002 31816
rect 262122 31804 262128 31816
rect 261996 31776 262128 31804
rect 261996 31764 262002 31776
rect 262122 31764 262128 31776
rect 262180 31764 262186 31816
rect 264698 31764 264704 31816
rect 264756 31804 264762 31816
rect 264882 31804 264888 31816
rect 264756 31776 264888 31804
rect 264756 31764 264762 31776
rect 264882 31764 264888 31776
rect 264940 31764 264946 31816
rect 19242 31696 19248 31748
rect 19300 31736 19306 31748
rect 36262 31736 36268 31748
rect 19300 31708 36268 31736
rect 19300 31696 19306 31708
rect 36262 31696 36268 31708
rect 36320 31696 36326 31748
rect 41322 31696 41328 31748
rect 41380 31736 41386 31748
rect 46934 31736 46940 31748
rect 41380 31708 46940 31736
rect 41380 31696 41386 31708
rect 46934 31696 46940 31708
rect 46992 31696 46998 31748
rect 110966 31696 110972 31748
rect 111024 31736 111030 31748
rect 160738 31736 160744 31748
rect 111024 31708 160744 31736
rect 111024 31696 111030 31708
rect 160738 31696 160744 31708
rect 160796 31696 160802 31748
rect 188982 31696 188988 31748
rect 189040 31736 189046 31748
rect 330478 31736 330484 31748
rect 189040 31708 330484 31736
rect 189040 31696 189046 31708
rect 330478 31696 330484 31708
rect 330536 31696 330542 31748
rect 16482 31628 16488 31680
rect 16540 31668 16546 31680
rect 35158 31668 35164 31680
rect 16540 31640 35164 31668
rect 16540 31628 16546 31640
rect 35158 31628 35164 31640
rect 35216 31628 35222 31680
rect 44082 31628 44088 31680
rect 44140 31668 44146 31680
rect 47946 31668 47952 31680
rect 44140 31640 47952 31668
rect 44140 31628 44146 31640
rect 47946 31628 47952 31640
rect 48004 31628 48010 31680
rect 68830 31628 68836 31680
rect 68888 31668 68894 31680
rect 68888 31640 75040 31668
rect 68888 31628 68894 31640
rect 20530 31560 20536 31612
rect 20588 31600 20594 31612
rect 37366 31600 37372 31612
rect 20588 31572 37372 31600
rect 20588 31560 20594 31572
rect 37366 31560 37372 31572
rect 37424 31560 37430 31612
rect 42702 31560 42708 31612
rect 42760 31600 42766 31612
rect 47394 31600 47400 31612
rect 42760 31572 47400 31600
rect 42760 31560 42766 31572
rect 47394 31560 47400 31572
rect 47452 31560 47458 31612
rect 75012 31600 75040 31640
rect 83182 31628 83188 31680
rect 83240 31668 83246 31680
rect 90266 31668 90272 31680
rect 83240 31640 90272 31668
rect 83240 31628 83246 31640
rect 90266 31628 90272 31640
rect 90324 31628 90330 31680
rect 90358 31628 90364 31680
rect 90416 31668 90422 31680
rect 94498 31668 94504 31680
rect 90416 31640 94504 31668
rect 90416 31628 90422 31640
rect 94498 31628 94504 31640
rect 94556 31628 94562 31680
rect 105998 31628 106004 31680
rect 106056 31668 106062 31680
rect 156598 31668 156604 31680
rect 106056 31640 156604 31668
rect 106056 31628 106062 31640
rect 156598 31628 156604 31640
rect 156656 31628 156662 31680
rect 188341 31671 188399 31677
rect 188341 31637 188353 31671
rect 188387 31668 188399 31671
rect 200758 31668 200764 31680
rect 188387 31640 200764 31668
rect 188387 31637 188399 31640
rect 188341 31631 188399 31637
rect 200758 31628 200764 31640
rect 200816 31628 200822 31680
rect 215662 31628 215668 31680
rect 215720 31668 215726 31680
rect 358078 31668 358084 31680
rect 215720 31640 358084 31668
rect 215720 31628 215726 31640
rect 358078 31628 358084 31640
rect 358136 31628 358142 31680
rect 85758 31600 85764 31612
rect 75012 31572 85764 31600
rect 85758 31560 85764 31572
rect 85816 31560 85822 31612
rect 93670 31560 93676 31612
rect 93728 31600 93734 31612
rect 95878 31600 95884 31612
rect 93728 31572 95884 31600
rect 93728 31560 93734 31572
rect 95878 31560 95884 31572
rect 95936 31560 95942 31612
rect 104342 31560 104348 31612
rect 104400 31600 104406 31612
rect 155218 31600 155224 31612
rect 104400 31572 155224 31600
rect 104400 31560 104406 31572
rect 155218 31560 155224 31572
rect 155276 31560 155282 31612
rect 165522 31560 165528 31612
rect 165580 31600 165586 31612
rect 204898 31600 204904 31612
rect 165580 31572 188476 31600
rect 165580 31560 165586 31572
rect 15102 31492 15108 31544
rect 15160 31532 15166 31544
rect 34606 31532 34612 31544
rect 15160 31504 34612 31532
rect 15160 31492 15166 31504
rect 34606 31492 34612 31504
rect 34664 31492 34670 31544
rect 38562 31492 38568 31544
rect 38620 31532 38626 31544
rect 45738 31532 45744 31544
rect 38620 31504 45744 31532
rect 38620 31492 38626 31504
rect 45738 31492 45744 31504
rect 45796 31492 45802 31544
rect 72602 31492 72608 31544
rect 72660 31532 72666 31544
rect 87506 31532 87512 31544
rect 72660 31504 87512 31532
rect 72660 31492 72666 31504
rect 87506 31492 87512 31504
rect 87564 31492 87570 31544
rect 112441 31535 112499 31541
rect 112441 31501 112453 31535
rect 112487 31532 112499 31535
rect 157978 31532 157984 31544
rect 112487 31504 157984 31532
rect 112487 31501 112499 31504
rect 112441 31495 112499 31501
rect 157978 31492 157984 31504
rect 158036 31492 158042 31544
rect 162210 31492 162216 31544
rect 162268 31532 162274 31544
rect 188341 31535 188399 31541
rect 188341 31532 188353 31535
rect 162268 31504 188353 31532
rect 162268 31492 162274 31504
rect 188341 31501 188353 31504
rect 188387 31501 188399 31535
rect 188448 31532 188476 31572
rect 193186 31572 204904 31600
rect 193186 31532 193214 31572
rect 204898 31560 204904 31572
rect 204956 31560 204962 31612
rect 209038 31560 209044 31612
rect 209096 31600 209102 31612
rect 351178 31600 351184 31612
rect 209096 31572 351184 31600
rect 209096 31560 209102 31572
rect 351178 31560 351184 31572
rect 351236 31560 351242 31612
rect 188448 31504 193214 31532
rect 188341 31495 188399 31501
rect 205542 31492 205548 31544
rect 205600 31532 205606 31544
rect 348418 31532 348424 31544
rect 205600 31504 348424 31532
rect 205600 31492 205606 31504
rect 348418 31492 348424 31504
rect 348476 31492 348482 31544
rect 13722 31424 13728 31476
rect 13780 31464 13786 31476
rect 34054 31464 34060 31476
rect 13780 31436 34060 31464
rect 13780 31424 13786 31436
rect 34054 31424 34060 31436
rect 34112 31424 34118 31476
rect 86494 31424 86500 31476
rect 86552 31464 86558 31476
rect 101398 31464 101404 31476
rect 86552 31436 101404 31464
rect 86552 31424 86558 31436
rect 101398 31424 101404 31436
rect 101456 31424 101462 31476
rect 159358 31464 159364 31476
rect 115906 31436 159364 31464
rect 10962 31356 10968 31408
rect 11020 31396 11026 31408
rect 32398 31396 32404 31408
rect 11020 31368 32404 31396
rect 11020 31356 11026 31368
rect 32398 31356 32404 31368
rect 32456 31356 32462 31408
rect 70946 31356 70952 31408
rect 71004 31396 71010 31408
rect 88978 31396 88984 31408
rect 71004 31368 88984 31396
rect 71004 31356 71010 31368
rect 88978 31356 88984 31368
rect 89036 31356 89042 31408
rect 105538 31396 105544 31408
rect 93826 31368 105544 31396
rect 12342 31288 12348 31340
rect 12400 31328 12406 31340
rect 33134 31328 33140 31340
rect 12400 31300 33140 31328
rect 12400 31288 12406 31300
rect 33134 31288 33140 31300
rect 33192 31288 33198 31340
rect 34422 31288 34428 31340
rect 34480 31328 34486 31340
rect 43530 31328 43536 31340
rect 34480 31300 43536 31328
rect 34480 31288 34486 31300
rect 43530 31288 43536 31300
rect 43588 31288 43594 31340
rect 45462 31288 45468 31340
rect 45520 31328 45526 31340
rect 48498 31328 48504 31340
rect 45520 31300 48504 31328
rect 45520 31288 45526 31300
rect 48498 31288 48504 31300
rect 48556 31288 48562 31340
rect 84838 31288 84844 31340
rect 84896 31328 84902 31340
rect 93826 31328 93854 31368
rect 105538 31356 105544 31368
rect 105596 31356 105602 31408
rect 109310 31356 109316 31408
rect 109368 31396 109374 31408
rect 115906 31396 115934 31436
rect 159358 31424 159364 31436
rect 159416 31424 159422 31476
rect 166902 31424 166908 31476
rect 166960 31464 166966 31476
rect 209038 31464 209044 31476
rect 166960 31436 209044 31464
rect 166960 31424 166966 31436
rect 209038 31424 209044 31436
rect 209096 31424 209102 31476
rect 237926 31424 237932 31476
rect 237984 31464 237990 31476
rect 238662 31464 238668 31476
rect 237984 31436 238668 31464
rect 237984 31424 237990 31436
rect 238662 31424 238668 31436
rect 238720 31424 238726 31476
rect 238757 31467 238815 31473
rect 238757 31433 238769 31467
rect 238803 31464 238815 31467
rect 376018 31464 376024 31476
rect 238803 31436 376024 31464
rect 238803 31433 238815 31436
rect 238757 31427 238815 31433
rect 376018 31424 376024 31436
rect 376076 31424 376082 31476
rect 109368 31368 115934 31396
rect 127529 31399 127587 31405
rect 109368 31356 109374 31368
rect 127529 31365 127541 31399
rect 127575 31396 127587 31399
rect 170398 31396 170404 31408
rect 127575 31368 170404 31396
rect 127575 31365 127587 31368
rect 127529 31359 127587 31365
rect 170398 31356 170404 31368
rect 170456 31356 170462 31408
rect 219066 31356 219072 31408
rect 219124 31396 219130 31408
rect 362218 31396 362224 31408
rect 219124 31368 362224 31396
rect 219124 31356 219130 31368
rect 362218 31356 362224 31368
rect 362276 31356 362282 31408
rect 84896 31300 93854 31328
rect 84896 31288 84902 31300
rect 115842 31288 115848 31340
rect 115900 31328 115906 31340
rect 169018 31328 169024 31340
rect 115900 31300 169024 31328
rect 115900 31288 115906 31300
rect 169018 31288 169024 31300
rect 169076 31288 169082 31340
rect 198642 31288 198648 31340
rect 198700 31328 198706 31340
rect 341518 31328 341524 31340
rect 198700 31300 341524 31328
rect 198700 31288 198706 31300
rect 341518 31288 341524 31300
rect 341576 31288 341582 31340
rect 9582 31220 9588 31272
rect 9640 31260 9646 31272
rect 31846 31260 31852 31272
rect 9640 31232 31852 31260
rect 9640 31220 9646 31232
rect 31846 31220 31852 31232
rect 31904 31220 31910 31272
rect 35802 31220 35808 31272
rect 35860 31260 35866 31272
rect 44174 31260 44180 31272
rect 35860 31232 44180 31260
rect 35860 31220 35866 31232
rect 44174 31220 44180 31232
rect 44232 31220 44238 31272
rect 77018 31220 77024 31272
rect 77076 31260 77082 31272
rect 102318 31260 102324 31272
rect 77076 31232 102324 31260
rect 77076 31220 77082 31232
rect 102318 31220 102324 31232
rect 102376 31220 102382 31272
rect 127621 31263 127679 31269
rect 127621 31229 127633 31263
rect 127667 31260 127679 31263
rect 166261 31263 166319 31269
rect 166261 31260 166273 31263
rect 127667 31232 166273 31260
rect 127667 31229 127679 31232
rect 127621 31223 127679 31229
rect 166261 31229 166273 31232
rect 166307 31229 166319 31263
rect 166261 31223 166319 31229
rect 225690 31220 225696 31272
rect 225748 31260 225754 31272
rect 369118 31260 369124 31272
rect 225748 31232 369124 31260
rect 225748 31220 225754 31232
rect 369118 31220 369124 31232
rect 369176 31220 369182 31272
rect 6822 31152 6828 31204
rect 6880 31192 6886 31204
rect 30742 31192 30748 31204
rect 6880 31164 30748 31192
rect 6880 31152 6886 31164
rect 30742 31152 30748 31164
rect 30800 31152 30806 31204
rect 33042 31152 33048 31204
rect 33100 31192 33106 31204
rect 42978 31192 42984 31204
rect 33100 31164 42984 31192
rect 33100 31152 33106 31164
rect 42978 31152 42984 31164
rect 43036 31152 43042 31204
rect 45370 31152 45376 31204
rect 45428 31192 45434 31204
rect 49142 31192 49148 31204
rect 45428 31164 49148 31192
rect 45428 31152 45434 31164
rect 49142 31152 49148 31164
rect 49200 31152 49206 31204
rect 78582 31152 78588 31204
rect 78640 31192 78646 31204
rect 104158 31192 104164 31204
rect 78640 31164 104164 31192
rect 78640 31152 78646 31164
rect 104158 31152 104164 31164
rect 104216 31152 104222 31204
rect 114370 31152 114376 31204
rect 114428 31192 114434 31204
rect 167638 31192 167644 31204
rect 114428 31164 167644 31192
rect 114428 31152 114434 31164
rect 167638 31152 167644 31164
rect 167696 31152 167702 31204
rect 212350 31152 212356 31204
rect 212408 31192 212414 31204
rect 355318 31192 355324 31204
rect 212408 31164 355324 31192
rect 212408 31152 212414 31164
rect 355318 31152 355324 31164
rect 355376 31152 355382 31204
rect 5442 31084 5448 31136
rect 5500 31124 5506 31136
rect 30374 31124 30380 31136
rect 5500 31096 30380 31124
rect 5500 31084 5506 31096
rect 30374 31084 30380 31096
rect 30432 31084 30438 31136
rect 31662 31084 31668 31136
rect 31720 31124 31726 31136
rect 42426 31124 42432 31136
rect 31720 31096 42432 31124
rect 31720 31084 31726 31096
rect 42426 31084 42432 31096
rect 42484 31084 42490 31136
rect 82078 31084 82084 31136
rect 82136 31124 82142 31136
rect 108298 31124 108304 31136
rect 82136 31096 108304 31124
rect 82136 31084 82142 31096
rect 108298 31084 108304 31096
rect 108356 31084 108362 31136
rect 112622 31084 112628 31136
rect 112680 31124 112686 31136
rect 166258 31124 166264 31136
rect 112680 31096 166264 31124
rect 112680 31084 112686 31096
rect 166258 31084 166264 31096
rect 166316 31084 166322 31136
rect 168926 31084 168932 31136
rect 168984 31124 168990 31136
rect 213178 31124 213184 31136
rect 168984 31096 213184 31124
rect 168984 31084 168990 31096
rect 213178 31084 213184 31096
rect 213236 31084 213242 31136
rect 222010 31084 222016 31136
rect 222068 31124 222074 31136
rect 366358 31124 366364 31136
rect 222068 31096 366364 31124
rect 222068 31084 222074 31096
rect 366358 31084 366364 31096
rect 366416 31084 366422 31136
rect 4062 31016 4068 31068
rect 4120 31056 4126 31068
rect 29638 31056 29644 31068
rect 4120 31028 29644 31056
rect 4120 31016 4126 31028
rect 29638 31016 29644 31028
rect 29696 31016 29702 31068
rect 30282 31016 30288 31068
rect 30340 31056 30346 31068
rect 41874 31056 41880 31068
rect 30340 31028 41880 31056
rect 30340 31016 30346 31028
rect 41874 31016 41880 31028
rect 41932 31016 41938 31068
rect 67542 31016 67548 31068
rect 67600 31056 67606 31068
rect 82998 31056 83004 31068
rect 67600 31028 83004 31056
rect 67600 31016 67606 31028
rect 82998 31016 83004 31028
rect 83056 31016 83062 31068
rect 85390 31016 85396 31068
rect 85448 31056 85454 31068
rect 119338 31056 119344 31068
rect 85448 31028 119344 31056
rect 85448 31016 85454 31028
rect 119338 31016 119344 31028
rect 119396 31016 119402 31068
rect 120994 31016 121000 31068
rect 121052 31056 121058 31068
rect 175918 31056 175924 31068
rect 121052 31028 175924 31056
rect 121052 31016 121058 31028
rect 175918 31016 175924 31028
rect 175976 31016 175982 31068
rect 180518 31016 180524 31068
rect 180576 31056 180582 31068
rect 185486 31056 185492 31068
rect 180576 31028 185492 31056
rect 180576 31016 180582 31028
rect 185486 31016 185492 31028
rect 185544 31016 185550 31068
rect 228910 31016 228916 31068
rect 228968 31056 228974 31068
rect 373258 31056 373264 31068
rect 228968 31028 373264 31056
rect 228968 31016 228974 31028
rect 373258 31016 373264 31028
rect 373316 31016 373322 31068
rect 23382 30948 23388 31000
rect 23440 30988 23446 31000
rect 38654 30988 38660 31000
rect 23440 30960 38660 30988
rect 23440 30948 23446 30960
rect 38654 30948 38660 30960
rect 38712 30948 38718 31000
rect 39942 30948 39948 31000
rect 40000 30988 40006 31000
rect 46290 30988 46296 31000
rect 40000 30960 46296 30988
rect 40000 30948 40006 30960
rect 46290 30948 46296 30960
rect 46348 30948 46354 31000
rect 119246 30948 119252 31000
rect 119304 30988 119310 31000
rect 127621 30991 127679 30997
rect 127621 30988 127633 30991
rect 119304 30960 127633 30988
rect 119304 30948 119310 30960
rect 127621 30957 127633 30960
rect 127667 30957 127679 30991
rect 127621 30951 127679 30957
rect 137281 30991 137339 30997
rect 137281 30957 137293 30991
rect 137327 30988 137339 30991
rect 177390 30988 177396 31000
rect 137327 30960 177396 30988
rect 137327 30957 137339 30960
rect 137281 30951 137339 30957
rect 177390 30948 177396 30960
rect 177448 30948 177454 31000
rect 192294 30948 192300 31000
rect 192352 30988 192358 31000
rect 195885 30991 195943 30997
rect 195885 30988 195897 30991
rect 192352 30960 195897 30988
rect 192352 30948 192358 30960
rect 195885 30957 195897 30960
rect 195931 30957 195943 30991
rect 195885 30951 195943 30957
rect 202322 30948 202328 31000
rect 202380 30988 202386 31000
rect 344278 30988 344284 31000
rect 202380 30960 344284 30988
rect 202380 30948 202386 30960
rect 344278 30948 344284 30960
rect 344336 30948 344342 31000
rect 20622 30880 20628 30932
rect 20680 30920 20686 30932
rect 36814 30920 36820 30932
rect 20680 30892 36820 30920
rect 20680 30880 20686 30892
rect 36814 30880 36820 30892
rect 36872 30880 36878 30932
rect 92290 30880 92296 30932
rect 92348 30920 92354 30932
rect 135438 30920 135444 30932
rect 92348 30892 135444 30920
rect 92348 30880 92354 30892
rect 135438 30880 135444 30892
rect 135496 30880 135502 30932
rect 145193 30923 145251 30929
rect 145193 30889 145205 30923
rect 145239 30920 145251 30923
rect 179966 30920 179972 30932
rect 145239 30892 179972 30920
rect 145239 30889 145251 30892
rect 145193 30883 145251 30889
rect 179966 30880 179972 30892
rect 180024 30880 180030 30932
rect 195606 30880 195612 30932
rect 195664 30920 195670 30932
rect 337378 30920 337384 30932
rect 195664 30892 337384 30920
rect 195664 30880 195670 30892
rect 337378 30880 337384 30892
rect 337436 30880 337442 30932
rect 22002 30812 22008 30864
rect 22060 30852 22066 30864
rect 37918 30852 37924 30864
rect 22060 30824 37924 30852
rect 22060 30812 22066 30824
rect 37918 30812 37924 30824
rect 37976 30812 37982 30864
rect 90910 30812 90916 30864
rect 90968 30852 90974 30864
rect 127621 30855 127679 30861
rect 127621 30852 127633 30855
rect 90968 30824 127633 30852
rect 90968 30812 90974 30824
rect 127621 30821 127633 30824
rect 127667 30821 127679 30855
rect 127621 30815 127679 30821
rect 139946 30812 139952 30864
rect 140004 30852 140010 30864
rect 181438 30852 181444 30864
rect 140004 30824 181444 30852
rect 140004 30812 140010 30824
rect 181438 30812 181444 30824
rect 181496 30812 181502 30864
rect 188430 30812 188436 30864
rect 188488 30852 188494 30864
rect 188982 30852 188988 30864
rect 188488 30824 188988 30852
rect 188488 30812 188494 30824
rect 188982 30812 188988 30824
rect 189040 30812 189046 30864
rect 195054 30812 195060 30864
rect 195112 30852 195118 30864
rect 195790 30852 195796 30864
rect 195112 30824 195796 30852
rect 195112 30812 195118 30824
rect 195790 30812 195796 30824
rect 195848 30812 195854 30864
rect 195885 30855 195943 30861
rect 195885 30821 195897 30855
rect 195931 30852 195943 30855
rect 333238 30852 333244 30864
rect 195931 30824 333244 30852
rect 195931 30821 195943 30824
rect 195885 30815 195943 30821
rect 333238 30812 333244 30824
rect 333296 30812 333302 30864
rect 24762 30744 24768 30796
rect 24820 30784 24826 30796
rect 39114 30784 39120 30796
rect 24820 30756 39120 30784
rect 24820 30744 24826 30756
rect 39114 30744 39120 30756
rect 39172 30744 39178 30796
rect 102042 30744 102048 30796
rect 102100 30784 102106 30796
rect 166261 30787 166319 30793
rect 102100 30756 132494 30784
rect 102100 30744 102106 30756
rect 28810 30676 28816 30728
rect 28868 30716 28874 30728
rect 41414 30716 41420 30728
rect 28868 30688 41420 30716
rect 28868 30676 28874 30688
rect 41414 30676 41420 30688
rect 41472 30676 41478 30728
rect 89622 30676 89628 30728
rect 89680 30716 89686 30728
rect 129734 30716 129740 30728
rect 89680 30688 129740 30716
rect 89680 30676 89686 30688
rect 129734 30676 129740 30688
rect 129792 30676 129798 30728
rect 132466 30716 132494 30756
rect 166261 30753 166273 30787
rect 166307 30784 166319 30787
rect 173158 30784 173164 30796
rect 166307 30756 173164 30784
rect 166307 30753 166319 30756
rect 166261 30747 166319 30753
rect 173158 30744 173164 30756
rect 173216 30744 173222 30796
rect 185578 30744 185584 30796
rect 185636 30784 185642 30796
rect 323670 30784 323676 30796
rect 185636 30756 323676 30784
rect 185636 30744 185642 30756
rect 323670 30744 323676 30756
rect 323728 30744 323734 30796
rect 142798 30716 142804 30728
rect 132466 30688 142804 30716
rect 142798 30676 142804 30688
rect 142856 30676 142862 30728
rect 175182 30676 175188 30728
rect 175240 30716 175246 30728
rect 301498 30716 301504 30728
rect 175240 30688 301504 30716
rect 175240 30676 175246 30688
rect 301498 30676 301504 30688
rect 301556 30676 301562 30728
rect 27522 30608 27528 30660
rect 27580 30648 27586 30660
rect 40218 30648 40224 30660
rect 27580 30620 40224 30648
rect 27580 30608 27586 30620
rect 40218 30608 40224 30620
rect 40276 30608 40282 30660
rect 88150 30608 88156 30660
rect 88208 30648 88214 30660
rect 127158 30648 127164 30660
rect 88208 30620 127164 30648
rect 88208 30608 88214 30620
rect 127158 30608 127164 30620
rect 127216 30608 127222 30660
rect 127621 30651 127679 30657
rect 127621 30617 127633 30651
rect 127667 30648 127679 30651
rect 132494 30648 132500 30660
rect 127667 30620 132500 30648
rect 127667 30617 127679 30620
rect 127621 30611 127679 30617
rect 132494 30608 132500 30620
rect 132552 30608 132558 30660
rect 136542 30608 136548 30660
rect 136600 30648 136606 30660
rect 136600 30620 137876 30648
rect 136600 30608 136606 30620
rect 26142 30540 26148 30592
rect 26200 30580 26206 30592
rect 39666 30580 39672 30592
rect 26200 30552 39672 30580
rect 26200 30540 26206 30552
rect 39666 30540 39672 30552
rect 39724 30540 39730 30592
rect 117682 30540 117688 30592
rect 117740 30580 117746 30592
rect 127529 30583 127587 30589
rect 127529 30580 127541 30583
rect 117740 30552 127541 30580
rect 117740 30540 117746 30552
rect 127529 30549 127541 30552
rect 127575 30549 127587 30583
rect 127529 30543 127587 30549
rect 128262 30540 128268 30592
rect 128320 30580 128326 30592
rect 137281 30583 137339 30589
rect 137281 30580 137293 30583
rect 128320 30552 137293 30580
rect 128320 30540 128326 30552
rect 137281 30549 137293 30552
rect 137327 30549 137339 30583
rect 137848 30580 137876 30620
rect 137922 30608 137928 30660
rect 137980 30648 137986 30660
rect 145193 30651 145251 30657
rect 145193 30648 145205 30651
rect 137980 30620 145205 30648
rect 137980 30608 137986 30620
rect 145193 30617 145205 30620
rect 145239 30617 145251 30651
rect 177206 30648 177212 30660
rect 145193 30611 145251 30617
rect 151786 30620 177212 30648
rect 151786 30580 151814 30620
rect 177206 30608 177212 30620
rect 177264 30608 177270 30660
rect 178954 30608 178960 30660
rect 179012 30648 179018 30660
rect 179012 30620 269620 30648
rect 179012 30608 179018 30620
rect 137848 30552 151814 30580
rect 137281 30543 137339 30549
rect 181162 30540 181168 30592
rect 181220 30580 181226 30592
rect 182082 30580 182088 30592
rect 181220 30552 182088 30580
rect 181220 30540 181226 30552
rect 182082 30540 182088 30552
rect 182140 30540 182146 30592
rect 183922 30540 183928 30592
rect 183980 30580 183986 30592
rect 184842 30580 184848 30592
rect 183980 30552 184848 30580
rect 183980 30540 183986 30552
rect 184842 30540 184848 30552
rect 184900 30540 184906 30592
rect 187326 30540 187332 30592
rect 187384 30580 187390 30592
rect 187602 30580 187608 30592
rect 187384 30552 187608 30580
rect 187384 30540 187390 30552
rect 187602 30540 187608 30552
rect 187660 30540 187666 30592
rect 203426 30540 203432 30592
rect 203484 30580 203490 30592
rect 204070 30580 204076 30592
rect 203484 30552 204076 30580
rect 203484 30540 203490 30552
rect 204070 30540 204076 30552
rect 204128 30540 204134 30592
rect 210694 30540 210700 30592
rect 210752 30580 210758 30592
rect 211062 30580 211068 30592
rect 210752 30552 211068 30580
rect 210752 30540 210758 30552
rect 211062 30540 211068 30552
rect 211120 30540 211126 30592
rect 224034 30540 224040 30592
rect 224092 30580 224098 30592
rect 224862 30580 224868 30592
rect 224092 30552 224868 30580
rect 224092 30540 224098 30552
rect 224862 30540 224868 30552
rect 224920 30540 224926 30592
rect 227346 30540 227352 30592
rect 227404 30580 227410 30592
rect 227622 30580 227628 30592
rect 227404 30552 227628 30580
rect 227404 30540 227410 30552
rect 227622 30540 227628 30552
rect 227680 30540 227686 30592
rect 232406 30540 232412 30592
rect 232464 30580 232470 30592
rect 238757 30583 238815 30589
rect 238757 30580 238769 30583
rect 232464 30552 238769 30580
rect 232464 30540 232470 30552
rect 238757 30549 238769 30552
rect 238803 30549 238815 30583
rect 238757 30543 238815 30549
rect 239493 30583 239551 30589
rect 239493 30549 239505 30583
rect 239539 30580 239551 30583
rect 269393 30583 269451 30589
rect 269393 30580 269405 30583
rect 239539 30552 269405 30580
rect 239539 30549 239551 30552
rect 239493 30543 239551 30549
rect 269393 30549 269405 30552
rect 269439 30549 269451 30583
rect 269393 30543 269451 30549
rect 28902 30472 28908 30524
rect 28960 30512 28966 30524
rect 40770 30512 40776 30524
rect 28960 30484 40776 30512
rect 28960 30472 28966 30484
rect 40770 30472 40776 30484
rect 40828 30472 40834 30524
rect 49602 30472 49608 30524
rect 49660 30512 49666 30524
rect 51074 30512 51080 30524
rect 49660 30484 51080 30512
rect 49660 30472 49666 30484
rect 51074 30472 51080 30484
rect 51132 30472 51138 30524
rect 172238 30472 172244 30524
rect 172296 30512 172302 30524
rect 244918 30512 244924 30524
rect 172296 30484 244924 30512
rect 172296 30472 172302 30484
rect 244918 30472 244924 30484
rect 244976 30472 244982 30524
rect 248233 30515 248291 30521
rect 248233 30512 248245 30515
rect 245396 30484 248245 30512
rect 37090 30404 37096 30456
rect 37148 30444 37154 30456
rect 45186 30444 45192 30456
rect 37148 30416 45192 30444
rect 37148 30404 37154 30416
rect 45186 30404 45192 30416
rect 45244 30404 45250 30456
rect 46842 30404 46848 30456
rect 46900 30444 46906 30456
rect 49694 30444 49700 30456
rect 46900 30416 49700 30444
rect 46900 30404 46906 30416
rect 49694 30404 49700 30416
rect 49752 30404 49758 30456
rect 63126 30404 63132 30456
rect 63184 30444 63190 30456
rect 63402 30444 63408 30456
rect 63184 30416 63408 30444
rect 63184 30404 63190 30416
rect 63402 30404 63408 30416
rect 63460 30404 63466 30456
rect 65886 30404 65892 30456
rect 65944 30444 65950 30456
rect 66162 30444 66168 30456
rect 65944 30416 66168 30444
rect 65944 30404 65950 30416
rect 66162 30404 66168 30416
rect 66220 30404 66226 30456
rect 88702 30404 88708 30456
rect 88760 30444 88766 30456
rect 93118 30444 93124 30456
rect 88760 30416 93124 30444
rect 88760 30404 88766 30416
rect 93118 30404 93124 30416
rect 93176 30404 93182 30456
rect 97074 30404 97080 30456
rect 97132 30444 97138 30456
rect 97902 30444 97908 30456
rect 97132 30416 97908 30444
rect 97132 30404 97138 30416
rect 97902 30404 97908 30416
rect 97960 30404 97966 30456
rect 100294 30404 100300 30456
rect 100352 30444 100358 30456
rect 100662 30444 100668 30456
rect 100352 30416 100668 30444
rect 100352 30404 100358 30416
rect 100662 30404 100668 30416
rect 100720 30404 100726 30456
rect 123846 30404 123852 30456
rect 123904 30444 123910 30456
rect 124122 30444 124128 30456
rect 123904 30416 124128 30444
rect 123904 30404 123910 30416
rect 124122 30404 124128 30416
rect 124180 30404 124186 30456
rect 128814 30404 128820 30456
rect 128872 30444 128878 30456
rect 129642 30444 129648 30456
rect 128872 30416 129648 30444
rect 128872 30404 128878 30416
rect 129642 30404 129648 30416
rect 129700 30404 129706 30456
rect 132126 30404 132132 30456
rect 132184 30444 132190 30456
rect 132402 30444 132408 30456
rect 132184 30416 132408 30444
rect 132184 30404 132190 30416
rect 132402 30404 132408 30416
rect 132460 30404 132466 30456
rect 149422 30404 149428 30456
rect 149480 30444 149486 30456
rect 150342 30444 150348 30456
rect 149480 30416 150348 30444
rect 149480 30404 149486 30416
rect 150342 30404 150348 30416
rect 150400 30404 150406 30456
rect 152734 30404 152740 30456
rect 152792 30444 152798 30456
rect 153102 30444 153108 30456
rect 152792 30416 153108 30444
rect 152792 30404 152798 30416
rect 153102 30404 153108 30416
rect 153160 30404 153166 30456
rect 158346 30404 158352 30456
rect 158404 30444 158410 30456
rect 158622 30444 158628 30456
rect 158404 30416 158628 30444
rect 158404 30404 158410 30416
rect 158622 30404 158628 30416
rect 158680 30404 158686 30456
rect 161106 30404 161112 30456
rect 161164 30444 161170 30456
rect 161382 30444 161388 30456
rect 161164 30416 161388 30444
rect 161164 30404 161170 30416
rect 161382 30404 161388 30416
rect 161440 30404 161446 30456
rect 163314 30404 163320 30456
rect 163372 30444 163378 30456
rect 164142 30444 164148 30456
rect 163372 30416 164148 30444
rect 163372 30404 163378 30416
rect 164142 30404 164148 30416
rect 164200 30404 164206 30456
rect 170582 30404 170588 30456
rect 170640 30444 170646 30456
rect 242158 30444 242164 30456
rect 170640 30416 242164 30444
rect 170640 30404 170646 30416
rect 242158 30404 242164 30416
rect 242216 30404 242222 30456
rect 242434 30404 242440 30456
rect 242492 30444 242498 30456
rect 245396 30444 245424 30484
rect 248233 30481 248245 30484
rect 248279 30481 248291 30515
rect 248233 30475 248291 30481
rect 250162 30472 250168 30524
rect 250220 30512 250226 30524
rect 250990 30512 250996 30524
rect 250220 30484 250996 30512
rect 250220 30472 250226 30484
rect 250990 30472 250996 30484
rect 251048 30472 251054 30524
rect 251910 30472 251916 30524
rect 251968 30512 251974 30524
rect 252462 30512 252468 30524
rect 251968 30484 252468 30512
rect 251968 30472 251974 30484
rect 252462 30472 252468 30484
rect 252520 30472 252526 30524
rect 253014 30472 253020 30524
rect 253072 30512 253078 30524
rect 253566 30512 253572 30524
rect 253072 30484 253572 30512
rect 253072 30472 253078 30484
rect 253566 30472 253572 30484
rect 253624 30472 253630 30524
rect 254670 30472 254676 30524
rect 254728 30512 254734 30524
rect 255130 30512 255136 30524
rect 254728 30484 255136 30512
rect 254728 30472 254734 30484
rect 255130 30472 255136 30484
rect 255188 30472 255194 30524
rect 255774 30472 255780 30524
rect 255832 30512 255838 30524
rect 256510 30512 256516 30524
rect 255832 30484 256516 30512
rect 255832 30472 255838 30484
rect 256510 30472 256516 30484
rect 256568 30472 256574 30524
rect 257430 30472 257436 30524
rect 257488 30512 257494 30524
rect 257982 30512 257988 30524
rect 257488 30484 257988 30512
rect 257488 30472 257494 30484
rect 257982 30472 257988 30484
rect 258040 30472 258046 30524
rect 259086 30472 259092 30524
rect 259144 30512 259150 30524
rect 259270 30512 259276 30524
rect 259144 30484 259276 30512
rect 259144 30472 259150 30484
rect 259270 30472 259276 30484
rect 259328 30472 259334 30524
rect 260190 30472 260196 30524
rect 260248 30512 260254 30524
rect 260742 30512 260748 30524
rect 260248 30484 260748 30512
rect 260248 30472 260254 30484
rect 260742 30472 260748 30484
rect 260800 30472 260806 30524
rect 261386 30472 261392 30524
rect 261444 30512 261450 30524
rect 261938 30512 261944 30524
rect 261444 30484 261944 30512
rect 261444 30472 261450 30484
rect 261938 30472 261944 30484
rect 261996 30472 262002 30524
rect 263042 30472 263048 30524
rect 263100 30512 263106 30524
rect 263502 30512 263508 30524
rect 263100 30484 263508 30512
rect 263100 30472 263106 30484
rect 263502 30472 263508 30484
rect 263560 30472 263566 30524
rect 264146 30472 264152 30524
rect 264204 30512 264210 30524
rect 264698 30512 264704 30524
rect 264204 30484 264704 30512
rect 264204 30472 264210 30484
rect 264698 30472 264704 30484
rect 264756 30472 264762 30524
rect 266906 30472 266912 30524
rect 266964 30512 266970 30524
rect 267550 30512 267556 30524
rect 266964 30484 267556 30512
rect 266964 30472 266970 30484
rect 267550 30472 267556 30484
rect 267608 30472 267614 30524
rect 268562 30472 268568 30524
rect 268620 30512 268626 30524
rect 269022 30512 269028 30524
rect 268620 30484 269028 30512
rect 268620 30472 268626 30484
rect 269022 30472 269028 30484
rect 269080 30472 269086 30524
rect 269592 30512 269620 30620
rect 269666 30608 269672 30660
rect 269724 30648 269730 30660
rect 270494 30648 270500 30660
rect 269724 30620 270500 30648
rect 269724 30608 269730 30620
rect 270494 30608 270500 30620
rect 270552 30608 270558 30660
rect 270589 30651 270647 30657
rect 270589 30617 270601 30651
rect 270635 30648 270647 30651
rect 276290 30648 276296 30660
rect 270635 30620 276296 30648
rect 270635 30617 270647 30620
rect 270589 30611 270647 30617
rect 276290 30608 276296 30620
rect 276348 30608 276354 30660
rect 276382 30608 276388 30660
rect 276440 30648 276446 30660
rect 277302 30648 277308 30660
rect 276440 30620 277308 30648
rect 276440 30608 276446 30620
rect 277302 30608 277308 30620
rect 277360 30608 277366 30660
rect 279694 30608 279700 30660
rect 279752 30648 279758 30660
rect 280062 30648 280068 30660
rect 279752 30620 280068 30648
rect 279752 30608 279758 30620
rect 280062 30608 280068 30620
rect 280120 30608 280126 30660
rect 284754 30608 284760 30660
rect 284812 30648 284818 30660
rect 285582 30648 285588 30660
rect 284812 30620 285588 30648
rect 284812 30608 284818 30620
rect 285582 30608 285588 30620
rect 285640 30608 285646 30660
rect 288066 30608 288072 30660
rect 288124 30648 288130 30660
rect 288342 30648 288348 30660
rect 288124 30620 288348 30648
rect 288124 30608 288130 30620
rect 288342 30608 288348 30620
rect 288400 30608 288406 30660
rect 293126 30608 293132 30660
rect 293184 30648 293190 30660
rect 293954 30648 293960 30660
rect 293184 30620 293960 30648
rect 293184 30608 293190 30620
rect 293954 30608 293960 30620
rect 294012 30608 294018 30660
rect 301406 30608 301412 30660
rect 301464 30648 301470 30660
rect 308398 30648 308404 30660
rect 301464 30620 308404 30648
rect 301464 30608 301470 30620
rect 308398 30608 308404 30620
rect 308456 30608 308462 30660
rect 269761 30583 269819 30589
rect 269761 30549 269773 30583
rect 269807 30580 269819 30583
rect 309778 30580 309784 30592
rect 269807 30552 309784 30580
rect 269807 30549 269819 30552
rect 269761 30543 269819 30549
rect 309778 30540 309784 30552
rect 309836 30540 309842 30592
rect 270129 30515 270187 30521
rect 270129 30512 270141 30515
rect 269592 30484 270141 30512
rect 270129 30481 270141 30484
rect 270175 30481 270187 30515
rect 270129 30475 270187 30481
rect 270218 30472 270224 30524
rect 270276 30512 270282 30524
rect 270402 30512 270408 30524
rect 270276 30484 270408 30512
rect 270276 30472 270282 30484
rect 270402 30472 270408 30484
rect 270460 30472 270466 30524
rect 271322 30472 271328 30524
rect 271380 30512 271386 30524
rect 271782 30512 271788 30524
rect 271380 30484 271788 30512
rect 271380 30472 271386 30484
rect 271782 30472 271788 30484
rect 271840 30472 271846 30524
rect 272518 30472 272524 30524
rect 272576 30512 272582 30524
rect 273070 30512 273076 30524
rect 272576 30484 273076 30512
rect 272576 30472 272582 30484
rect 273070 30472 273076 30484
rect 273128 30472 273134 30524
rect 273622 30472 273628 30524
rect 273680 30512 273686 30524
rect 274450 30512 274456 30524
rect 273680 30484 274456 30512
rect 273680 30472 273686 30484
rect 274450 30472 274456 30484
rect 274508 30472 274514 30524
rect 275278 30472 275284 30524
rect 275336 30512 275342 30524
rect 275922 30512 275928 30524
rect 275336 30484 275928 30512
rect 275336 30472 275342 30484
rect 275922 30472 275928 30484
rect 275980 30472 275986 30524
rect 276934 30472 276940 30524
rect 276992 30512 276998 30524
rect 277210 30512 277216 30524
rect 276992 30484 277216 30512
rect 276992 30472 276998 30484
rect 277210 30472 277216 30484
rect 277268 30472 277274 30524
rect 278038 30472 278044 30524
rect 278096 30512 278102 30524
rect 278682 30512 278688 30524
rect 278096 30484 278688 30512
rect 278096 30472 278102 30484
rect 278682 30472 278688 30484
rect 278740 30472 278746 30524
rect 279142 30472 279148 30524
rect 279200 30512 279206 30524
rect 279878 30512 279884 30524
rect 279200 30484 279884 30512
rect 279200 30472 279206 30484
rect 279878 30472 279884 30484
rect 279936 30472 279942 30524
rect 280798 30472 280804 30524
rect 280856 30512 280862 30524
rect 281350 30512 281356 30524
rect 280856 30484 281356 30512
rect 280856 30472 280862 30484
rect 281350 30472 281356 30484
rect 281408 30472 281414 30524
rect 281902 30472 281908 30524
rect 281960 30512 281966 30524
rect 282730 30512 282736 30524
rect 281960 30484 282736 30512
rect 281960 30472 281966 30484
rect 282730 30472 282736 30484
rect 282788 30472 282794 30524
rect 283650 30472 283656 30524
rect 283708 30512 283714 30524
rect 284202 30512 284208 30524
rect 283708 30484 284208 30512
rect 283708 30472 283714 30484
rect 284202 30472 284208 30484
rect 284260 30472 284266 30524
rect 285306 30472 285312 30524
rect 285364 30512 285370 30524
rect 285490 30512 285496 30524
rect 285364 30484 285496 30512
rect 285364 30472 285370 30484
rect 285490 30472 285496 30484
rect 285548 30472 285554 30524
rect 286410 30472 286416 30524
rect 286468 30512 286474 30524
rect 286962 30512 286968 30524
rect 286468 30484 286968 30512
rect 286468 30472 286474 30484
rect 286962 30472 286968 30484
rect 287020 30472 287026 30524
rect 287514 30472 287520 30524
rect 287572 30512 287578 30524
rect 288158 30512 288164 30524
rect 287572 30484 288164 30512
rect 287572 30472 287578 30484
rect 288158 30472 288164 30484
rect 288216 30472 288222 30524
rect 289170 30472 289176 30524
rect 289228 30512 289234 30524
rect 289630 30512 289636 30524
rect 289228 30484 289636 30512
rect 289228 30472 289234 30484
rect 289630 30472 289636 30484
rect 289688 30472 289694 30524
rect 290274 30472 290280 30524
rect 290332 30512 290338 30524
rect 291010 30512 291016 30524
rect 290332 30484 291016 30512
rect 290332 30472 290338 30484
rect 291010 30472 291016 30484
rect 291068 30472 291074 30524
rect 291930 30472 291936 30524
rect 291988 30512 291994 30524
rect 292390 30512 292396 30524
rect 291988 30484 292396 30512
rect 291988 30472 291994 30484
rect 292390 30472 292396 30484
rect 292448 30472 292454 30524
rect 293678 30472 293684 30524
rect 293736 30512 293742 30524
rect 293862 30512 293868 30524
rect 293736 30484 293868 30512
rect 293736 30472 293742 30484
rect 293862 30472 293868 30484
rect 293920 30472 293926 30524
rect 294782 30472 294788 30524
rect 294840 30512 294846 30524
rect 295242 30512 295248 30524
rect 294840 30484 295248 30512
rect 294840 30472 294846 30484
rect 295242 30472 295248 30484
rect 295300 30472 295306 30524
rect 295886 30472 295892 30524
rect 295944 30512 295950 30524
rect 296438 30512 296444 30524
rect 295944 30484 296444 30512
rect 295944 30472 295950 30484
rect 296438 30472 296444 30484
rect 296496 30472 296502 30524
rect 298646 30472 298652 30524
rect 298704 30512 298710 30524
rect 299290 30512 299296 30524
rect 298704 30484 299296 30512
rect 298704 30472 298710 30484
rect 299290 30472 299296 30484
rect 299348 30472 299354 30524
rect 301958 30472 301964 30524
rect 302016 30512 302022 30524
rect 304258 30512 304264 30524
rect 302016 30484 304264 30512
rect 302016 30472 302022 30484
rect 304258 30472 304264 30484
rect 304316 30472 304322 30524
rect 242492 30416 245424 30444
rect 242492 30404 242498 30416
rect 245470 30404 245476 30456
rect 245528 30444 245534 30456
rect 315390 30444 315396 30456
rect 245528 30416 315396 30444
rect 245528 30404 245534 30416
rect 315390 30404 315396 30416
rect 315448 30404 315454 30456
rect 37182 30336 37188 30388
rect 37240 30376 37246 30388
rect 44634 30376 44640 30388
rect 37240 30348 44640 30376
rect 37240 30336 37246 30348
rect 44634 30336 44640 30348
rect 44692 30336 44698 30388
rect 48222 30336 48228 30388
rect 48280 30376 48286 30388
rect 50246 30376 50252 30388
rect 48280 30348 50252 30376
rect 48280 30336 48286 30348
rect 50246 30336 50252 30348
rect 50304 30336 50310 30388
rect 52454 30336 52460 30388
rect 52512 30376 52518 30388
rect 53006 30376 53012 30388
rect 52512 30348 53012 30376
rect 52512 30336 52518 30348
rect 53006 30336 53012 30348
rect 53064 30336 53070 30388
rect 54754 30336 54760 30388
rect 54812 30376 54818 30388
rect 55122 30376 55128 30388
rect 54812 30348 55128 30376
rect 54812 30336 54818 30348
rect 55122 30336 55128 30348
rect 55180 30336 55186 30388
rect 55858 30336 55864 30388
rect 55916 30376 55922 30388
rect 56410 30376 56416 30388
rect 55916 30348 56416 30376
rect 55916 30336 55922 30348
rect 56410 30336 56416 30348
rect 56468 30336 56474 30388
rect 56962 30336 56968 30388
rect 57020 30376 57026 30388
rect 57790 30376 57796 30388
rect 57020 30348 57796 30376
rect 57020 30336 57026 30348
rect 57790 30336 57796 30348
rect 57848 30336 57854 30388
rect 58618 30336 58624 30388
rect 58676 30376 58682 30388
rect 59170 30376 59176 30388
rect 58676 30348 59176 30376
rect 58676 30336 58682 30348
rect 59170 30336 59176 30348
rect 59228 30336 59234 30388
rect 59722 30336 59728 30388
rect 59780 30376 59786 30388
rect 60642 30376 60648 30388
rect 59780 30348 60648 30376
rect 59780 30336 59786 30348
rect 60642 30336 60648 30348
rect 60700 30336 60706 30388
rect 61470 30336 61476 30388
rect 61528 30376 61534 30388
rect 62022 30376 62028 30388
rect 61528 30348 62028 30376
rect 61528 30336 61534 30348
rect 62022 30336 62028 30348
rect 62080 30336 62086 30388
rect 62574 30336 62580 30388
rect 62632 30376 62638 30388
rect 63218 30376 63224 30388
rect 62632 30348 63224 30376
rect 62632 30336 62638 30348
rect 63218 30336 63224 30348
rect 63276 30336 63282 30388
rect 64230 30336 64236 30388
rect 64288 30376 64294 30388
rect 64690 30376 64696 30388
rect 64288 30348 64696 30376
rect 64288 30336 64294 30348
rect 64690 30336 64696 30348
rect 64748 30336 64754 30388
rect 65334 30336 65340 30388
rect 65392 30376 65398 30388
rect 65978 30376 65984 30388
rect 65392 30348 65984 30376
rect 65392 30336 65398 30348
rect 65978 30336 65984 30348
rect 66036 30336 66042 30388
rect 66990 30336 66996 30388
rect 67048 30376 67054 30388
rect 67542 30376 67548 30388
rect 67048 30348 67548 30376
rect 67048 30336 67054 30348
rect 67542 30336 67548 30348
rect 67600 30336 67606 30388
rect 68094 30336 68100 30388
rect 68152 30376 68158 30388
rect 68922 30376 68928 30388
rect 68152 30348 68928 30376
rect 68152 30336 68158 30348
rect 68922 30336 68928 30348
rect 68980 30336 68986 30388
rect 69750 30336 69756 30388
rect 69808 30376 69814 30388
rect 70302 30376 70308 30388
rect 69808 30348 70308 30376
rect 69808 30336 69814 30348
rect 70302 30336 70308 30348
rect 70360 30336 70366 30388
rect 71498 30336 71504 30388
rect 71556 30376 71562 30388
rect 71682 30376 71688 30388
rect 71556 30348 71688 30376
rect 71556 30336 71562 30348
rect 71682 30336 71688 30348
rect 71740 30336 71746 30388
rect 73706 30336 73712 30388
rect 73764 30376 73770 30388
rect 74350 30376 74356 30388
rect 73764 30348 74356 30376
rect 73764 30336 73770 30348
rect 74350 30336 74356 30348
rect 74408 30336 74414 30388
rect 76466 30336 76472 30388
rect 76524 30376 76530 30388
rect 77110 30376 77116 30388
rect 76524 30348 77116 30376
rect 76524 30336 76530 30348
rect 77110 30336 77116 30348
rect 77168 30336 77174 30388
rect 78122 30336 78128 30388
rect 78180 30376 78186 30388
rect 78582 30376 78588 30388
rect 78180 30348 78588 30376
rect 78180 30336 78186 30348
rect 78582 30336 78588 30348
rect 78640 30336 78646 30388
rect 79226 30336 79232 30388
rect 79284 30376 79290 30388
rect 79870 30376 79876 30388
rect 79284 30348 79876 30376
rect 79284 30336 79290 30348
rect 79870 30336 79876 30348
rect 79928 30336 79934 30388
rect 80882 30336 80888 30388
rect 80940 30376 80946 30388
rect 81342 30376 81348 30388
rect 80940 30348 81348 30376
rect 80940 30336 80946 30348
rect 81342 30336 81348 30348
rect 81400 30336 81406 30388
rect 85942 30336 85948 30388
rect 86000 30376 86006 30388
rect 86770 30376 86776 30388
rect 86000 30348 86776 30376
rect 86000 30336 86006 30348
rect 86770 30336 86776 30348
rect 86828 30336 86834 30388
rect 87598 30336 87604 30388
rect 87656 30376 87662 30388
rect 88242 30376 88248 30388
rect 87656 30348 88248 30376
rect 87656 30336 87662 30348
rect 88242 30336 88248 30348
rect 88300 30336 88306 30388
rect 91462 30336 91468 30388
rect 91520 30376 91526 30388
rect 92290 30376 92296 30388
rect 91520 30348 92296 30376
rect 91520 30336 91526 30348
rect 92290 30336 92296 30348
rect 92348 30336 92354 30388
rect 93210 30336 93216 30388
rect 93268 30376 93274 30388
rect 93762 30376 93768 30388
rect 93268 30348 93768 30376
rect 93268 30336 93274 30348
rect 93762 30336 93768 30348
rect 93820 30336 93826 30388
rect 94314 30336 94320 30388
rect 94372 30376 94378 30388
rect 94866 30376 94872 30388
rect 94372 30348 94872 30376
rect 94372 30336 94378 30348
rect 94866 30336 94872 30348
rect 94924 30336 94930 30388
rect 95970 30336 95976 30388
rect 96028 30376 96034 30388
rect 96430 30376 96436 30388
rect 96028 30348 96436 30376
rect 96028 30336 96034 30348
rect 96430 30336 96436 30348
rect 96488 30336 96494 30388
rect 97626 30336 97632 30388
rect 97684 30376 97690 30388
rect 97810 30376 97816 30388
rect 97684 30348 97816 30376
rect 97684 30336 97690 30348
rect 97810 30336 97816 30348
rect 97868 30336 97874 30388
rect 98730 30336 98736 30388
rect 98788 30376 98794 30388
rect 99282 30376 99288 30388
rect 98788 30348 99288 30376
rect 98788 30336 98794 30348
rect 99282 30336 99288 30348
rect 99340 30336 99346 30388
rect 99834 30336 99840 30388
rect 99892 30376 99898 30388
rect 100570 30376 100576 30388
rect 99892 30348 100576 30376
rect 99892 30336 99898 30348
rect 100570 30336 100576 30348
rect 100628 30336 100634 30388
rect 101490 30336 101496 30388
rect 101548 30376 101554 30388
rect 102042 30376 102048 30388
rect 101548 30348 102048 30376
rect 101548 30336 101554 30348
rect 102042 30336 102048 30348
rect 102100 30336 102106 30388
rect 102686 30336 102692 30388
rect 102744 30376 102750 30388
rect 103238 30376 103244 30388
rect 102744 30348 103244 30376
rect 102744 30336 102750 30348
rect 103238 30336 103244 30348
rect 103296 30336 103302 30388
rect 105446 30336 105452 30388
rect 105504 30376 105510 30388
rect 106182 30376 106188 30388
rect 105504 30348 106188 30376
rect 105504 30336 105510 30348
rect 106182 30336 106188 30348
rect 106240 30336 106246 30388
rect 107102 30336 107108 30388
rect 107160 30376 107166 30388
rect 107562 30376 107568 30388
rect 107160 30348 107568 30376
rect 107160 30336 107166 30348
rect 107562 30336 107568 30348
rect 107620 30336 107626 30388
rect 108206 30336 108212 30388
rect 108264 30376 108270 30388
rect 108758 30376 108764 30388
rect 108264 30348 108764 30376
rect 108264 30336 108270 30348
rect 108758 30336 108764 30348
rect 108816 30336 108822 30388
rect 113818 30336 113824 30388
rect 113876 30376 113882 30388
rect 114462 30376 114468 30388
rect 113876 30348 114468 30376
rect 113876 30336 113882 30348
rect 114462 30336 114468 30348
rect 114520 30336 114526 30388
rect 114922 30336 114928 30388
rect 114980 30376 114986 30388
rect 115750 30376 115756 30388
rect 114980 30348 115756 30376
rect 114980 30336 114986 30348
rect 115750 30336 115756 30348
rect 115808 30336 115814 30388
rect 116578 30336 116584 30388
rect 116636 30376 116642 30388
rect 117130 30376 117136 30388
rect 116636 30348 117136 30376
rect 116636 30336 116642 30348
rect 117130 30336 117136 30348
rect 117188 30336 117194 30388
rect 120442 30336 120448 30388
rect 120500 30376 120506 30388
rect 121362 30376 121368 30388
rect 120500 30348 121368 30376
rect 120500 30336 120506 30348
rect 121362 30336 121368 30348
rect 121420 30336 121426 30388
rect 122098 30336 122104 30388
rect 122156 30376 122162 30388
rect 122742 30376 122748 30388
rect 122156 30348 122748 30376
rect 122156 30336 122162 30348
rect 122742 30336 122748 30348
rect 122800 30336 122806 30388
rect 123202 30336 123208 30388
rect 123260 30376 123266 30388
rect 123938 30376 123944 30388
rect 123260 30348 123944 30376
rect 123260 30336 123266 30348
rect 123938 30336 123944 30348
rect 123996 30336 124002 30388
rect 124950 30336 124956 30388
rect 125008 30376 125014 30388
rect 125410 30376 125416 30388
rect 125008 30348 125416 30376
rect 125008 30336 125014 30348
rect 125410 30336 125416 30348
rect 125468 30336 125474 30388
rect 126054 30336 126060 30388
rect 126112 30376 126118 30388
rect 126790 30376 126796 30388
rect 126112 30348 126796 30376
rect 126112 30336 126118 30348
rect 126790 30336 126796 30348
rect 126848 30336 126854 30388
rect 127710 30336 127716 30388
rect 127768 30376 127774 30388
rect 128262 30376 128268 30388
rect 127768 30348 128268 30376
rect 127768 30336 127774 30348
rect 128262 30336 128268 30348
rect 128320 30336 128326 30388
rect 129366 30336 129372 30388
rect 129424 30376 129430 30388
rect 129550 30376 129556 30388
rect 129424 30348 129556 30376
rect 129424 30336 129430 30348
rect 129550 30336 129556 30348
rect 129608 30336 129614 30388
rect 130470 30336 130476 30388
rect 130528 30376 130534 30388
rect 131022 30376 131028 30388
rect 130528 30348 131028 30376
rect 130528 30336 130534 30348
rect 131022 30336 131028 30348
rect 131080 30336 131086 30388
rect 131574 30336 131580 30388
rect 131632 30376 131638 30388
rect 132218 30376 132224 30388
rect 131632 30348 132224 30376
rect 131632 30336 131638 30348
rect 132218 30336 132224 30348
rect 132276 30336 132282 30388
rect 133230 30336 133236 30388
rect 133288 30376 133294 30388
rect 133690 30376 133696 30388
rect 133288 30348 133696 30376
rect 133288 30336 133294 30348
rect 133690 30336 133696 30348
rect 133748 30336 133754 30388
rect 134426 30336 134432 30388
rect 134484 30376 134490 30388
rect 135070 30376 135076 30388
rect 134484 30348 135076 30376
rect 134484 30336 134490 30348
rect 135070 30336 135076 30348
rect 135128 30336 135134 30388
rect 136082 30336 136088 30388
rect 136140 30376 136146 30388
rect 136542 30376 136548 30388
rect 136140 30348 136548 30376
rect 136140 30336 136146 30348
rect 136542 30336 136548 30348
rect 136600 30336 136606 30388
rect 137186 30336 137192 30388
rect 137244 30376 137250 30388
rect 137922 30376 137928 30388
rect 137244 30348 137928 30376
rect 137244 30336 137250 30348
rect 137922 30336 137928 30348
rect 137980 30336 137986 30388
rect 140498 30336 140504 30388
rect 140556 30376 140562 30388
rect 140682 30376 140688 30388
rect 140556 30348 140688 30376
rect 140556 30336 140562 30348
rect 140682 30336 140688 30348
rect 140740 30336 140746 30388
rect 141602 30336 141608 30388
rect 141660 30376 141666 30388
rect 142062 30376 142068 30388
rect 141660 30348 142068 30376
rect 141660 30336 141666 30348
rect 142062 30336 142068 30348
rect 142120 30336 142126 30388
rect 142706 30336 142712 30388
rect 142764 30376 142770 30388
rect 142764 30348 143212 30376
rect 142764 30336 142770 30348
rect 143184 30240 143212 30348
rect 143258 30336 143264 30388
rect 143316 30376 143322 30388
rect 143442 30376 143448 30388
rect 143316 30348 143448 30376
rect 143316 30336 143322 30348
rect 143442 30336 143448 30348
rect 143500 30336 143506 30388
rect 144362 30336 144368 30388
rect 144420 30376 144426 30388
rect 144822 30376 144828 30388
rect 144420 30348 144828 30376
rect 144420 30336 144426 30348
rect 144822 30336 144828 30348
rect 144880 30336 144886 30388
rect 145558 30336 145564 30388
rect 145616 30376 145622 30388
rect 146110 30376 146116 30388
rect 145616 30348 146116 30376
rect 145616 30336 145622 30348
rect 146110 30336 146116 30348
rect 146168 30336 146174 30388
rect 146662 30336 146668 30388
rect 146720 30376 146726 30388
rect 147490 30376 147496 30388
rect 146720 30348 147496 30376
rect 146720 30336 146726 30348
rect 147490 30336 147496 30348
rect 147548 30336 147554 30388
rect 148318 30336 148324 30388
rect 148376 30376 148382 30388
rect 148962 30376 148968 30388
rect 148376 30348 148968 30376
rect 148376 30336 148382 30348
rect 148962 30336 148968 30348
rect 149020 30336 149026 30388
rect 149974 30336 149980 30388
rect 150032 30376 150038 30388
rect 150250 30376 150256 30388
rect 150032 30348 150256 30376
rect 150032 30336 150038 30348
rect 150250 30336 150256 30348
rect 150308 30336 150314 30388
rect 151078 30336 151084 30388
rect 151136 30376 151142 30388
rect 151722 30376 151728 30388
rect 151136 30348 151728 30376
rect 151136 30336 151142 30348
rect 151722 30336 151728 30348
rect 151780 30336 151786 30388
rect 152182 30336 152188 30388
rect 152240 30376 152246 30388
rect 152918 30376 152924 30388
rect 152240 30348 152924 30376
rect 152240 30336 152246 30348
rect 152918 30336 152924 30348
rect 152976 30336 152982 30388
rect 153838 30336 153844 30388
rect 153896 30376 153902 30388
rect 154390 30376 154396 30388
rect 153896 30348 154396 30376
rect 153896 30336 153902 30348
rect 154390 30336 154396 30348
rect 154448 30336 154454 30388
rect 154942 30336 154948 30388
rect 155000 30376 155006 30388
rect 155770 30376 155776 30388
rect 155000 30348 155776 30376
rect 155000 30336 155006 30348
rect 155770 30336 155776 30348
rect 155828 30336 155834 30388
rect 156690 30336 156696 30388
rect 156748 30376 156754 30388
rect 157242 30376 157248 30388
rect 156748 30348 157248 30376
rect 156748 30336 156754 30348
rect 157242 30336 157248 30348
rect 157300 30336 157306 30388
rect 157794 30336 157800 30388
rect 157852 30376 157858 30388
rect 158438 30376 158444 30388
rect 157852 30348 158444 30376
rect 157852 30336 157858 30348
rect 158438 30336 158444 30348
rect 158496 30336 158502 30388
rect 159450 30336 159456 30388
rect 159508 30376 159514 30388
rect 159910 30376 159916 30388
rect 159508 30348 159916 30376
rect 159508 30336 159514 30348
rect 159910 30336 159916 30348
rect 159968 30336 159974 30388
rect 160554 30336 160560 30388
rect 160612 30376 160618 30388
rect 161198 30376 161204 30388
rect 160612 30348 161204 30376
rect 160612 30336 160618 30348
rect 161198 30336 161204 30348
rect 161256 30336 161262 30388
rect 163866 30336 163872 30388
rect 163924 30376 163930 30388
rect 164050 30376 164056 30388
rect 163924 30348 164056 30376
rect 163924 30336 163930 30348
rect 164050 30336 164056 30348
rect 164108 30336 164114 30388
rect 164970 30336 164976 30388
rect 165028 30376 165034 30388
rect 165522 30376 165528 30388
rect 165028 30348 165528 30376
rect 165028 30336 165034 30348
rect 165522 30336 165528 30348
rect 165580 30336 165586 30388
rect 166166 30336 166172 30388
rect 166224 30376 166230 30388
rect 166902 30376 166908 30388
rect 166224 30348 166908 30376
rect 166224 30336 166230 30348
rect 166902 30336 166908 30348
rect 166960 30336 166966 30388
rect 171686 30336 171692 30388
rect 171744 30376 171750 30388
rect 172422 30376 172428 30388
rect 171744 30348 172428 30376
rect 171744 30336 171750 30348
rect 172422 30336 172428 30348
rect 172480 30336 172486 30388
rect 173342 30336 173348 30388
rect 173400 30376 173406 30388
rect 173802 30376 173808 30388
rect 173400 30348 173808 30376
rect 173400 30336 173406 30348
rect 173802 30336 173808 30348
rect 173860 30336 173866 30388
rect 174446 30336 174452 30388
rect 174504 30376 174510 30388
rect 174998 30376 175004 30388
rect 174504 30348 175004 30376
rect 174504 30336 174510 30348
rect 174998 30336 175004 30348
rect 175056 30336 175062 30388
rect 177298 30336 177304 30388
rect 177356 30376 177362 30388
rect 177850 30376 177856 30388
rect 177356 30348 177856 30376
rect 177356 30336 177362 30348
rect 177850 30336 177856 30348
rect 177908 30336 177914 30388
rect 178402 30336 178408 30388
rect 178460 30376 178466 30388
rect 179230 30376 179236 30388
rect 178460 30348 179236 30376
rect 178460 30336 178466 30348
rect 179230 30336 179236 30348
rect 179288 30336 179294 30388
rect 180058 30336 180064 30388
rect 180116 30376 180122 30388
rect 180702 30376 180708 30388
rect 180116 30348 180708 30376
rect 180116 30336 180122 30348
rect 180702 30336 180708 30348
rect 180760 30336 180766 30388
rect 181714 30336 181720 30388
rect 181772 30376 181778 30388
rect 181990 30376 181996 30388
rect 181772 30348 181996 30376
rect 181772 30336 181778 30348
rect 181990 30336 181996 30348
rect 182048 30336 182054 30388
rect 182818 30336 182824 30388
rect 182876 30376 182882 30388
rect 183462 30376 183468 30388
rect 182876 30348 183468 30376
rect 182876 30336 182882 30348
rect 183462 30336 183468 30348
rect 183520 30336 183526 30388
rect 184474 30336 184480 30388
rect 184532 30376 184538 30388
rect 184750 30376 184756 30388
rect 184532 30348 184756 30376
rect 184532 30336 184538 30348
rect 184750 30336 184756 30348
rect 184808 30336 184814 30388
rect 186682 30336 186688 30388
rect 186740 30376 186746 30388
rect 187418 30376 187424 30388
rect 186740 30348 187424 30376
rect 186740 30336 186746 30348
rect 187418 30336 187424 30348
rect 187476 30336 187482 30388
rect 189534 30336 189540 30388
rect 189592 30376 189598 30388
rect 190270 30376 190276 30388
rect 189592 30348 190276 30376
rect 189592 30336 189598 30348
rect 190270 30336 190276 30348
rect 190328 30336 190334 30388
rect 191190 30336 191196 30388
rect 191248 30376 191254 30388
rect 191742 30376 191748 30388
rect 191248 30348 191748 30376
rect 191248 30336 191254 30348
rect 191742 30336 191748 30348
rect 191800 30336 191806 30388
rect 192846 30336 192852 30388
rect 192904 30376 192910 30388
rect 193122 30376 193128 30388
rect 192904 30348 193128 30376
rect 192904 30336 192910 30348
rect 193122 30336 193128 30348
rect 193180 30336 193186 30388
rect 193950 30336 193956 30388
rect 194008 30376 194014 30388
rect 194502 30376 194508 30388
rect 194008 30348 194508 30376
rect 194008 30336 194014 30348
rect 194502 30336 194508 30348
rect 194560 30336 194566 30388
rect 196710 30336 196716 30388
rect 196768 30376 196774 30388
rect 197170 30376 197176 30388
rect 196768 30348 197176 30376
rect 196768 30336 196774 30348
rect 197170 30336 197176 30348
rect 197228 30336 197234 30388
rect 197906 30336 197912 30388
rect 197964 30376 197970 30388
rect 198642 30376 198648 30388
rect 197964 30348 198648 30376
rect 197964 30336 197970 30348
rect 198642 30336 198648 30348
rect 198700 30336 198706 30388
rect 199562 30336 199568 30388
rect 199620 30376 199626 30388
rect 200022 30376 200028 30388
rect 199620 30348 200028 30376
rect 199620 30336 199626 30348
rect 200022 30336 200028 30348
rect 200080 30336 200086 30388
rect 200666 30336 200672 30388
rect 200724 30376 200730 30388
rect 200724 30348 201172 30376
rect 200724 30336 200730 30348
rect 143442 30240 143448 30252
rect 143184 30212 143448 30240
rect 143442 30200 143448 30212
rect 143500 30200 143506 30252
rect 201144 30240 201172 30348
rect 201218 30336 201224 30388
rect 201276 30376 201282 30388
rect 201402 30376 201408 30388
rect 201276 30348 201408 30376
rect 201276 30336 201282 30348
rect 201402 30336 201408 30348
rect 201460 30336 201466 30388
rect 203886 30336 203892 30388
rect 203944 30376 203950 30388
rect 204162 30376 204168 30388
rect 203944 30348 204168 30376
rect 203944 30336 203950 30348
rect 204162 30336 204168 30348
rect 204220 30336 204226 30388
rect 205082 30336 205088 30388
rect 205140 30376 205146 30388
rect 205542 30376 205548 30388
rect 205140 30348 205548 30376
rect 205140 30336 205146 30348
rect 205542 30336 205548 30348
rect 205600 30336 205606 30388
rect 206186 30336 206192 30388
rect 206244 30376 206250 30388
rect 206738 30376 206744 30388
rect 206244 30348 206744 30376
rect 206244 30336 206250 30348
rect 206738 30336 206744 30348
rect 206796 30336 206802 30388
rect 210142 30336 210148 30388
rect 210200 30376 210206 30388
rect 210878 30376 210884 30388
rect 210200 30348 210884 30376
rect 210200 30336 210206 30348
rect 210878 30336 210884 30348
rect 210936 30336 210942 30388
rect 211798 30336 211804 30388
rect 211856 30376 211862 30388
rect 212442 30376 212448 30388
rect 211856 30348 212448 30376
rect 211856 30336 211862 30348
rect 212442 30336 212448 30348
rect 212500 30336 212506 30388
rect 212902 30336 212908 30388
rect 212960 30376 212966 30388
rect 213730 30376 213736 30388
rect 212960 30348 213736 30376
rect 212960 30336 212966 30348
rect 213730 30336 213736 30348
rect 213788 30336 213794 30388
rect 214558 30336 214564 30388
rect 214616 30376 214622 30388
rect 215202 30376 215208 30388
rect 214616 30348 215208 30376
rect 214616 30336 214622 30348
rect 215202 30336 215208 30348
rect 215260 30336 215266 30388
rect 216214 30336 216220 30388
rect 216272 30376 216278 30388
rect 216582 30376 216588 30388
rect 216272 30348 216588 30376
rect 216272 30336 216278 30348
rect 216582 30336 216588 30348
rect 216640 30336 216646 30388
rect 217318 30336 217324 30388
rect 217376 30376 217382 30388
rect 217962 30376 217968 30388
rect 217376 30348 217968 30376
rect 217376 30336 217382 30348
rect 217962 30336 217968 30348
rect 218020 30336 218026 30388
rect 218422 30336 218428 30388
rect 218480 30376 218486 30388
rect 219250 30376 219256 30388
rect 218480 30348 219256 30376
rect 218480 30336 218486 30348
rect 219250 30336 219256 30348
rect 219308 30336 219314 30388
rect 220170 30336 220176 30388
rect 220228 30376 220234 30388
rect 220630 30376 220636 30388
rect 220228 30348 220636 30376
rect 220228 30336 220234 30348
rect 220630 30336 220636 30348
rect 220688 30336 220694 30388
rect 221274 30336 221280 30388
rect 221332 30376 221338 30388
rect 222102 30376 222108 30388
rect 221332 30348 222108 30376
rect 221332 30336 221338 30348
rect 222102 30336 222108 30348
rect 222160 30336 222166 30388
rect 222930 30336 222936 30388
rect 222988 30376 222994 30388
rect 223482 30376 223488 30388
rect 222988 30348 223488 30376
rect 222988 30336 222994 30348
rect 223482 30336 223488 30348
rect 223540 30336 223546 30388
rect 224586 30336 224592 30388
rect 224644 30376 224650 30388
rect 224770 30376 224776 30388
rect 224644 30348 224776 30376
rect 224644 30336 224650 30348
rect 224770 30336 224776 30348
rect 224828 30336 224834 30388
rect 226794 30336 226800 30388
rect 226852 30376 226858 30388
rect 227438 30376 227444 30388
rect 226852 30348 227444 30376
rect 226852 30336 226858 30348
rect 227438 30336 227444 30348
rect 227496 30336 227502 30388
rect 228450 30336 228456 30388
rect 228508 30376 228514 30388
rect 229002 30376 229008 30388
rect 228508 30348 229008 30376
rect 228508 30336 228514 30348
rect 229002 30336 229008 30348
rect 229060 30336 229066 30388
rect 229646 30336 229652 30388
rect 229704 30376 229710 30388
rect 230290 30376 230296 30388
rect 229704 30348 230296 30376
rect 229704 30336 229710 30348
rect 230290 30336 230296 30348
rect 230348 30336 230354 30388
rect 231302 30336 231308 30388
rect 231360 30376 231366 30388
rect 231762 30376 231768 30388
rect 231360 30348 231768 30376
rect 231360 30336 231366 30348
rect 231762 30336 231768 30348
rect 231820 30336 231826 30388
rect 232958 30336 232964 30388
rect 233016 30376 233022 30388
rect 233142 30376 233148 30388
rect 233016 30348 233148 30376
rect 233016 30336 233022 30348
rect 233142 30336 233148 30348
rect 233200 30336 233206 30388
rect 235166 30336 235172 30388
rect 235224 30376 235230 30388
rect 235810 30376 235816 30388
rect 235224 30348 235816 30376
rect 235224 30336 235230 30348
rect 235810 30336 235816 30348
rect 235868 30336 235874 30388
rect 239493 30379 239551 30385
rect 239493 30376 239505 30379
rect 235920 30348 239505 30376
rect 235718 30268 235724 30320
rect 235776 30308 235782 30320
rect 235920 30308 235948 30348
rect 239493 30345 239505 30348
rect 239539 30345 239551 30379
rect 239493 30339 239551 30345
rect 239582 30336 239588 30388
rect 239640 30376 239646 30388
rect 240042 30376 240048 30388
rect 239640 30348 240048 30376
rect 239640 30336 239646 30348
rect 240042 30336 240048 30348
rect 240100 30336 240106 30388
rect 240778 30336 240784 30388
rect 240836 30376 240842 30388
rect 241330 30376 241336 30388
rect 240836 30348 241336 30376
rect 240836 30336 240842 30348
rect 241330 30336 241336 30348
rect 241388 30336 241394 30388
rect 241882 30336 241888 30388
rect 241940 30376 241946 30388
rect 242710 30376 242716 30388
rect 241940 30348 242716 30376
rect 241940 30336 241946 30348
rect 242710 30336 242716 30348
rect 242768 30336 242774 30388
rect 243538 30336 243544 30388
rect 243596 30376 243602 30388
rect 244182 30376 244188 30388
rect 243596 30348 244188 30376
rect 243596 30336 243602 30348
rect 244182 30336 244188 30348
rect 244240 30336 244246 30388
rect 244642 30336 244648 30388
rect 244700 30376 244706 30388
rect 245562 30376 245568 30388
rect 244700 30348 245568 30376
rect 244700 30336 244706 30348
rect 245562 30336 245568 30348
rect 245620 30336 245626 30388
rect 246298 30336 246304 30388
rect 246356 30376 246362 30388
rect 246942 30376 246948 30388
rect 246356 30348 246948 30376
rect 246356 30336 246362 30348
rect 246942 30336 246948 30348
rect 247000 30336 247006 30388
rect 247402 30336 247408 30388
rect 247460 30376 247466 30388
rect 248138 30376 248144 30388
rect 247460 30348 248144 30376
rect 247460 30336 247466 30348
rect 248138 30336 248144 30348
rect 248196 30336 248202 30388
rect 248233 30379 248291 30385
rect 248233 30345 248245 30379
rect 248279 30376 248291 30379
rect 312538 30376 312544 30388
rect 248279 30348 312544 30376
rect 248279 30345 248291 30348
rect 248233 30339 248291 30345
rect 312538 30336 312544 30348
rect 312596 30336 312602 30388
rect 235776 30280 235948 30308
rect 235776 30268 235782 30280
rect 201402 30240 201408 30252
rect 201144 30212 201408 30240
rect 201402 30200 201408 30212
rect 201460 30200 201466 30252
rect 296622 30200 296628 30252
rect 296680 30200 296686 30252
rect 296530 29996 296536 30048
rect 296588 30036 296594 30048
rect 296640 30036 296668 30200
rect 296588 30008 296668 30036
rect 296588 29996 296594 30008
rect 258534 27276 258540 27328
rect 258592 27316 258598 27328
rect 259362 27316 259368 27328
rect 258592 27288 259368 27316
rect 258592 27276 258598 27288
rect 259362 27276 259368 27288
rect 259420 27276 259426 27328
rect 302878 20612 302884 20664
rect 302936 20652 302942 20664
rect 579982 20652 579988 20664
rect 302936 20624 579988 20652
rect 302936 20612 302942 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 234430 16056 234436 16108
rect 234488 16096 234494 16108
rect 436738 16096 436744 16108
rect 234488 16068 436744 16096
rect 234488 16056 234494 16068
rect 436738 16056 436744 16068
rect 436796 16056 436802 16108
rect 241330 15988 241336 16040
rect 241388 16028 241394 16040
rect 450906 16028 450912 16040
rect 241388 16000 450912 16028
rect 241388 15988 241394 16000
rect 450906 15988 450912 16000
rect 450964 15988 450970 16040
rect 244090 15920 244096 15972
rect 244148 15960 244154 15972
rect 456794 15960 456800 15972
rect 244148 15932 456800 15960
rect 244148 15920 244154 15932
rect 456794 15920 456800 15932
rect 456852 15920 456858 15972
rect 248138 15852 248144 15904
rect 248196 15892 248202 15904
rect 465166 15892 465172 15904
rect 248196 15864 465172 15892
rect 248196 15852 248202 15864
rect 465166 15852 465172 15864
rect 465224 15852 465230 15904
rect 227438 15104 227444 15156
rect 227496 15144 227502 15156
rect 420914 15144 420920 15156
rect 227496 15116 420920 15144
rect 227496 15104 227502 15116
rect 420914 15104 420920 15116
rect 420972 15104 420978 15156
rect 229002 15036 229008 15088
rect 229060 15076 229066 15088
rect 423674 15076 423680 15088
rect 229060 15048 423680 15076
rect 229060 15036 229066 15048
rect 423674 15036 423680 15048
rect 423732 15036 423738 15088
rect 230198 14968 230204 15020
rect 230256 15008 230262 15020
rect 428458 15008 428464 15020
rect 230256 14980 428464 15008
rect 230256 14968 230262 14980
rect 428458 14968 428464 14980
rect 428516 14968 428522 15020
rect 231670 14900 231676 14952
rect 231728 14940 231734 14952
rect 432046 14940 432052 14952
rect 231728 14912 432052 14940
rect 231728 14900 231734 14912
rect 432046 14900 432052 14912
rect 432104 14900 432110 14952
rect 233050 14832 233056 14884
rect 233108 14872 233114 14884
rect 435082 14872 435088 14884
rect 233108 14844 435088 14872
rect 233108 14832 233114 14844
rect 435082 14832 435088 14844
rect 435140 14832 435146 14884
rect 248230 14764 248236 14816
rect 248288 14804 248294 14816
rect 465810 14804 465816 14816
rect 248288 14776 465816 14804
rect 248288 14764 248294 14776
rect 465810 14764 465816 14776
rect 465868 14764 465874 14816
rect 249702 14696 249708 14748
rect 249760 14736 249766 14748
rect 469858 14736 469864 14748
rect 249760 14708 469864 14736
rect 249760 14696 249766 14708
rect 469858 14696 469864 14708
rect 469916 14696 469922 14748
rect 253658 14628 253664 14680
rect 253716 14668 253722 14680
rect 476482 14668 476488 14680
rect 253716 14640 476488 14668
rect 253716 14628 253722 14640
rect 476482 14628 476488 14640
rect 476540 14628 476546 14680
rect 250898 14560 250904 14612
rect 250956 14600 250962 14612
rect 473446 14600 473452 14612
rect 250956 14572 473452 14600
rect 250956 14560 250962 14572
rect 473446 14560 473452 14572
rect 473504 14560 473510 14612
rect 290918 14492 290924 14544
rect 290976 14532 290982 14544
rect 556890 14532 556896 14544
rect 290976 14504 556896 14532
rect 290976 14492 290982 14504
rect 556890 14492 556896 14504
rect 556948 14492 556954 14544
rect 292390 14424 292396 14476
rect 292448 14464 292454 14476
rect 559282 14464 559288 14476
rect 292448 14436 559288 14464
rect 292448 14424 292454 14436
rect 559282 14424 559288 14436
rect 559340 14424 559346 14476
rect 208210 14356 208216 14408
rect 208268 14396 208274 14408
rect 381170 14396 381176 14408
rect 208268 14368 381176 14396
rect 208268 14356 208274 14368
rect 381170 14356 381176 14368
rect 381228 14356 381234 14408
rect 206738 14288 206744 14340
rect 206796 14328 206802 14340
rect 377674 14328 377680 14340
rect 206796 14300 377680 14328
rect 206796 14288 206802 14300
rect 377674 14288 377680 14300
rect 377732 14288 377738 14340
rect 184658 14220 184664 14272
rect 184716 14260 184722 14272
rect 332686 14260 332692 14272
rect 184716 14232 332692 14260
rect 184716 14220 184722 14232
rect 332686 14220 332692 14232
rect 332744 14220 332750 14272
rect 187418 14152 187424 14204
rect 187476 14192 187482 14204
rect 336274 14192 336280 14204
rect 187476 14164 336280 14192
rect 187476 14152 187482 14164
rect 336274 14152 336280 14164
rect 336332 14152 336338 14204
rect 183370 14084 183376 14136
rect 183428 14124 183434 14136
rect 328730 14124 328736 14136
rect 183428 14096 328736 14124
rect 183428 14084 183434 14096
rect 328730 14084 328736 14096
rect 328788 14084 328794 14136
rect 181898 14016 181904 14068
rect 181956 14056 181962 14068
rect 326338 14056 326344 14068
rect 181956 14028 326344 14056
rect 181956 14016 181962 14028
rect 326338 14016 326344 14028
rect 326396 14016 326402 14068
rect 181990 13948 181996 14000
rect 182048 13988 182054 14000
rect 324314 13988 324320 14000
rect 182048 13960 324320 13988
rect 182048 13948 182054 13960
rect 324314 13948 324320 13960
rect 324372 13948 324378 14000
rect 177850 13880 177856 13932
rect 177908 13920 177914 13932
rect 316034 13920 316040 13932
rect 177908 13892 316040 13920
rect 177908 13880 177914 13892
rect 316034 13880 316040 13892
rect 316092 13880 316098 13932
rect 173710 13812 173716 13864
rect 173768 13852 173774 13864
rect 307754 13852 307760 13864
rect 173768 13824 307760 13852
rect 173768 13812 173774 13824
rect 307754 13812 307760 13824
rect 307812 13812 307818 13864
rect 257890 13744 257896 13796
rect 257948 13784 257954 13796
rect 487154 13784 487160 13796
rect 257948 13756 487160 13784
rect 257948 13744 257954 13756
rect 487154 13744 487160 13756
rect 487212 13744 487218 13796
rect 259178 13676 259184 13728
rect 259236 13716 259242 13728
rect 489914 13716 489920 13728
rect 259236 13688 489920 13716
rect 259236 13676 259242 13688
rect 489914 13676 489920 13688
rect 489972 13676 489978 13728
rect 261938 13608 261944 13660
rect 261996 13648 262002 13660
rect 494698 13648 494704 13660
rect 261996 13620 494704 13648
rect 261996 13608 262002 13620
rect 494698 13608 494704 13620
rect 494756 13608 494762 13660
rect 275830 13540 275836 13592
rect 275888 13580 275894 13592
rect 525426 13580 525432 13592
rect 275888 13552 525432 13580
rect 275888 13540 275894 13552
rect 525426 13540 525432 13552
rect 525484 13540 525490 13592
rect 277118 13472 277124 13524
rect 277176 13512 277182 13524
rect 528554 13512 528560 13524
rect 277176 13484 528560 13512
rect 277176 13472 277182 13484
rect 528554 13472 528560 13484
rect 528612 13472 528618 13524
rect 158438 13404 158444 13456
rect 158496 13444 158502 13456
rect 274818 13444 274824 13456
rect 158496 13416 274824 13444
rect 158496 13404 158502 13416
rect 274818 13404 274824 13416
rect 274876 13404 274882 13456
rect 279878 13404 279884 13456
rect 279936 13444 279942 13456
rect 532050 13444 532056 13456
rect 279936 13416 532056 13444
rect 279936 13404 279942 13416
rect 532050 13404 532056 13416
rect 532108 13404 532114 13456
rect 159910 13336 159916 13388
rect 159968 13376 159974 13388
rect 278314 13376 278320 13388
rect 159968 13348 278320 13376
rect 159968 13336 159974 13348
rect 278314 13336 278320 13348
rect 278372 13336 278378 13388
rect 281350 13336 281356 13388
rect 281408 13376 281414 13388
rect 536098 13376 536104 13388
rect 281408 13348 536104 13376
rect 281408 13336 281414 13348
rect 536098 13336 536104 13348
rect 536156 13336 536162 13388
rect 162762 13268 162768 13320
rect 162820 13308 162826 13320
rect 284938 13308 284944 13320
rect 162820 13280 284944 13308
rect 162820 13268 162826 13280
rect 284938 13268 284944 13280
rect 284996 13268 285002 13320
rect 285398 13268 285404 13320
rect 285456 13308 285462 13320
rect 546678 13308 546684 13320
rect 285456 13280 546684 13308
rect 285456 13268 285462 13280
rect 546678 13268 546684 13280
rect 546736 13268 546742 13320
rect 163958 13200 163964 13252
rect 164016 13240 164022 13252
rect 288986 13240 288992 13252
rect 164016 13212 288992 13240
rect 164016 13200 164022 13212
rect 288986 13200 288992 13212
rect 289044 13200 289050 13252
rect 289630 13200 289636 13252
rect 289688 13240 289694 13252
rect 553762 13240 553768 13252
rect 289688 13212 553768 13240
rect 289688 13200 289694 13212
rect 553762 13200 553768 13212
rect 553820 13200 553826 13252
rect 169570 13132 169576 13184
rect 169628 13172 169634 13184
rect 299658 13172 299664 13184
rect 169628 13144 299664 13172
rect 169628 13132 169634 13144
rect 299658 13132 299664 13144
rect 299716 13132 299722 13184
rect 300670 13132 300676 13184
rect 300728 13172 300734 13184
rect 576946 13172 576952 13184
rect 300728 13144 576952 13172
rect 300728 13132 300734 13144
rect 576946 13132 576952 13144
rect 577004 13132 577010 13184
rect 171042 13064 171048 13116
rect 171100 13104 171106 13116
rect 303154 13104 303160 13116
rect 171100 13076 303160 13104
rect 171100 13064 171106 13076
rect 303154 13064 303160 13076
rect 303212 13064 303218 13116
rect 304258 13064 304264 13116
rect 304316 13104 304322 13116
rect 581730 13104 581736 13116
rect 304316 13076 581736 13104
rect 304316 13064 304322 13076
rect 581730 13064 581736 13076
rect 581788 13064 581794 13116
rect 256418 12996 256424 13048
rect 256476 13036 256482 13048
rect 484026 13036 484032 13048
rect 256476 13008 484032 13036
rect 256476 12996 256482 13008
rect 484026 12996 484032 13008
rect 484084 12996 484090 13048
rect 255130 12928 255136 12980
rect 255188 12968 255194 12980
rect 480530 12968 480536 12980
rect 255188 12940 480536 12968
rect 255188 12928 255194 12940
rect 480530 12928 480536 12940
rect 480588 12928 480594 12980
rect 203978 12860 203984 12912
rect 204036 12900 204042 12912
rect 374086 12900 374092 12912
rect 204036 12872 374092 12900
rect 204036 12860 204042 12872
rect 374086 12860 374092 12872
rect 374144 12860 374150 12912
rect 202782 12792 202788 12844
rect 202840 12832 202846 12844
rect 370130 12832 370136 12844
rect 202840 12804 370136 12832
rect 202840 12792 202846 12804
rect 370130 12792 370136 12804
rect 370188 12792 370194 12844
rect 177942 12724 177948 12776
rect 178000 12764 178006 12776
rect 317322 12764 317328 12776
rect 178000 12736 317328 12764
rect 178000 12724 178006 12736
rect 317322 12724 317328 12736
rect 317380 12724 317386 12776
rect 176470 12656 176476 12708
rect 176528 12696 176534 12708
rect 313826 12696 313832 12708
rect 176528 12668 313832 12696
rect 176528 12656 176534 12668
rect 313826 12656 313832 12668
rect 313884 12656 313890 12708
rect 172330 12588 172336 12640
rect 172388 12628 172394 12640
rect 306374 12628 306380 12640
rect 172388 12600 306380 12628
rect 172388 12588 172394 12600
rect 306374 12588 306380 12600
rect 306432 12588 306438 12640
rect 175090 12520 175096 12572
rect 175148 12560 175154 12572
rect 309686 12560 309692 12572
rect 175148 12532 309692 12560
rect 175148 12520 175154 12532
rect 309686 12520 309692 12532
rect 309744 12520 309750 12572
rect 168190 12452 168196 12504
rect 168248 12492 168254 12504
rect 295610 12492 295616 12504
rect 168248 12464 295616 12492
rect 168248 12452 168254 12464
rect 295610 12452 295616 12464
rect 295668 12452 295674 12504
rect 296438 12452 296444 12504
rect 296496 12492 296502 12504
rect 418798 12492 418804 12504
rect 296496 12464 418804 12492
rect 296496 12452 296502 12464
rect 418798 12452 418804 12464
rect 418856 12452 418862 12504
rect 250990 12384 250996 12436
rect 251048 12424 251054 12436
rect 470594 12424 470600 12436
rect 251048 12396 470600 12424
rect 251048 12384 251054 12396
rect 470594 12384 470600 12396
rect 470652 12384 470658 12436
rect 252462 12316 252468 12368
rect 252520 12356 252526 12368
rect 474090 12356 474096 12368
rect 252520 12328 474096 12356
rect 252520 12316 252526 12328
rect 474090 12316 474096 12328
rect 474148 12316 474154 12368
rect 253750 12248 253756 12300
rect 253808 12288 253814 12300
rect 478138 12288 478144 12300
rect 253808 12260 478144 12288
rect 253808 12248 253814 12260
rect 478138 12248 478144 12260
rect 478196 12248 478202 12300
rect 256510 12180 256516 12232
rect 256568 12220 256574 12232
rect 482370 12220 482376 12232
rect 256568 12192 482376 12220
rect 256568 12180 256574 12192
rect 482370 12180 482376 12192
rect 482428 12180 482434 12232
rect 257982 12112 257988 12164
rect 258040 12152 258046 12164
rect 486418 12152 486424 12164
rect 258040 12124 486424 12152
rect 258040 12112 258046 12124
rect 486418 12112 486424 12124
rect 486476 12112 486482 12164
rect 259270 12044 259276 12096
rect 259328 12084 259334 12096
rect 490006 12084 490012 12096
rect 259328 12056 490012 12084
rect 259328 12044 259334 12056
rect 490006 12044 490012 12056
rect 490064 12044 490070 12096
rect 260650 11976 260656 12028
rect 260708 12016 260714 12028
rect 493042 12016 493048 12028
rect 260708 11988 493048 12016
rect 260708 11976 260714 11988
rect 493042 11976 493048 11988
rect 493100 11976 493106 12028
rect 262030 11908 262036 11960
rect 262088 11948 262094 11960
rect 497090 11948 497096 11960
rect 262088 11920 497096 11948
rect 262088 11908 262094 11920
rect 497090 11908 497096 11920
rect 497148 11908 497154 11960
rect 264698 11840 264704 11892
rect 264756 11880 264762 11892
rect 500586 11880 500592 11892
rect 264756 11852 500592 11880
rect 264756 11840 264762 11852
rect 500586 11840 500592 11852
rect 500644 11840 500650 11892
rect 266170 11772 266176 11824
rect 266228 11812 266234 11824
rect 503714 11812 503720 11824
rect 266228 11784 503720 11812
rect 266228 11772 266234 11784
rect 503714 11772 503720 11784
rect 503772 11772 503778 11824
rect 267458 11704 267464 11756
rect 267516 11744 267522 11756
rect 507210 11744 507216 11756
rect 267516 11716 507216 11744
rect 267516 11704 267522 11716
rect 507210 11704 507216 11716
rect 507268 11704 507274 11756
rect 248322 11636 248328 11688
rect 248380 11676 248386 11688
rect 467466 11676 467472 11688
rect 248380 11648 467472 11676
rect 248380 11636 248386 11648
rect 467466 11636 467472 11648
rect 467524 11636 467530 11688
rect 246850 11568 246856 11620
rect 246908 11608 246914 11620
rect 463970 11608 463976 11620
rect 246908 11580 463976 11608
rect 246908 11568 246914 11580
rect 463970 11568 463976 11580
rect 464028 11568 464034 11620
rect 245470 11500 245476 11552
rect 245528 11540 245534 11552
rect 459922 11540 459928 11552
rect 245528 11512 459928 11540
rect 245528 11500 245534 11512
rect 459922 11500 459928 11512
rect 459980 11500 459986 11552
rect 244182 11432 244188 11484
rect 244240 11472 244246 11484
rect 456886 11472 456892 11484
rect 244240 11444 456892 11472
rect 244240 11432 244246 11444
rect 456886 11432 456892 11444
rect 456944 11432 456950 11484
rect 242710 11364 242716 11416
rect 242768 11404 242774 11416
rect 453298 11404 453304 11416
rect 242768 11376 453304 11404
rect 242768 11364 242774 11376
rect 453298 11364 453304 11376
rect 453356 11364 453362 11416
rect 239950 11296 239956 11348
rect 240008 11336 240014 11348
rect 448514 11336 448520 11348
rect 240008 11308 448520 11336
rect 240008 11296 240014 11308
rect 448514 11296 448520 11308
rect 448572 11296 448578 11348
rect 238570 11228 238576 11280
rect 238628 11268 238634 11280
rect 445754 11268 445760 11280
rect 238628 11240 445760 11268
rect 238628 11228 238634 11240
rect 445754 11228 445760 11240
rect 445812 11228 445818 11280
rect 235810 11160 235816 11212
rect 235868 11200 235874 11212
rect 439130 11200 439136 11212
rect 235868 11172 439136 11200
rect 235868 11160 235874 11172
rect 439130 11160 439136 11172
rect 439188 11160 439194 11212
rect 164050 11092 164056 11144
rect 164108 11132 164114 11144
rect 287330 11132 287336 11144
rect 164108 11104 287336 11132
rect 164108 11092 164114 11104
rect 287330 11092 287336 11104
rect 287388 11092 287394 11144
rect 201218 10956 201224 11008
rect 201276 10996 201282 11008
rect 367738 10996 367744 11008
rect 201276 10968 367744 10996
rect 201276 10956 201282 10968
rect 367738 10956 367744 10968
rect 367796 10956 367802 11008
rect 204070 10888 204076 10940
rect 204128 10928 204134 10940
rect 371234 10928 371240 10940
rect 204128 10900 371240 10928
rect 204128 10888 204134 10900
rect 371234 10888 371240 10900
rect 371292 10888 371298 10940
rect 205542 10820 205548 10872
rect 205600 10860 205606 10872
rect 375282 10860 375288 10872
rect 205600 10832 375288 10860
rect 205600 10820 205606 10832
rect 375282 10820 375288 10832
rect 375340 10820 375346 10872
rect 206830 10752 206836 10804
rect 206888 10792 206894 10804
rect 378410 10792 378416 10804
rect 206888 10764 378416 10792
rect 206888 10752 206894 10764
rect 378410 10752 378416 10764
rect 378468 10752 378474 10804
rect 208302 10684 208308 10736
rect 208360 10724 208366 10736
rect 382366 10724 382372 10736
rect 208360 10696 382372 10724
rect 208360 10684 208366 10696
rect 382366 10684 382372 10696
rect 382424 10684 382430 10736
rect 210878 10616 210884 10668
rect 210936 10656 210942 10668
rect 385954 10656 385960 10668
rect 210936 10628 385960 10656
rect 210936 10616 210942 10628
rect 385954 10616 385960 10628
rect 386012 10616 386018 10668
rect 212442 10548 212448 10600
rect 212500 10588 212506 10600
rect 389450 10588 389456 10600
rect 212500 10560 389456 10588
rect 212500 10548 212506 10560
rect 389450 10548 389456 10560
rect 389508 10548 389514 10600
rect 213638 10480 213644 10532
rect 213696 10520 213702 10532
rect 392578 10520 392584 10532
rect 213696 10492 392584 10520
rect 213696 10480 213702 10492
rect 392578 10480 392584 10492
rect 392636 10480 392642 10532
rect 215110 10412 215116 10464
rect 215168 10452 215174 10464
rect 396074 10452 396080 10464
rect 215168 10424 396080 10452
rect 215168 10412 215174 10424
rect 396074 10412 396080 10424
rect 396132 10412 396138 10464
rect 216490 10344 216496 10396
rect 216548 10384 216554 10396
rect 398834 10384 398840 10396
rect 216548 10356 398840 10384
rect 216548 10344 216554 10356
rect 398834 10344 398840 10356
rect 398892 10344 398898 10396
rect 219250 10276 219256 10328
rect 219308 10316 219314 10328
rect 403618 10316 403624 10328
rect 219308 10288 403624 10316
rect 219308 10276 219314 10288
rect 403618 10276 403624 10288
rect 403676 10276 403682 10328
rect 199930 10208 199936 10260
rect 199988 10248 199994 10260
rect 364610 10248 364616 10260
rect 199988 10220 364616 10248
rect 199988 10208 199994 10220
rect 364610 10208 364616 10220
rect 364668 10208 364674 10260
rect 198550 10140 198556 10192
rect 198608 10180 198614 10192
rect 361114 10180 361120 10192
rect 198608 10152 361120 10180
rect 198608 10140 198614 10152
rect 361114 10140 361120 10152
rect 361172 10140 361178 10192
rect 197170 10072 197176 10124
rect 197228 10112 197234 10124
rect 357526 10112 357532 10124
rect 197228 10084 357532 10112
rect 197228 10072 197234 10084
rect 357526 10072 357532 10084
rect 357584 10072 357590 10124
rect 195790 10004 195796 10056
rect 195848 10044 195854 10056
rect 353570 10044 353576 10056
rect 195848 10016 353576 10044
rect 195848 10004 195854 10016
rect 353570 10004 353576 10016
rect 353628 10004 353634 10056
rect 193030 9936 193036 9988
rect 193088 9976 193094 9988
rect 349154 9976 349160 9988
rect 193088 9948 349160 9976
rect 193088 9936 193094 9948
rect 349154 9936 349160 9948
rect 349212 9936 349218 9988
rect 191650 9868 191656 9920
rect 191708 9908 191714 9920
rect 346946 9908 346952 9920
rect 191708 9880 346952 9908
rect 191708 9868 191714 9880
rect 346946 9868 346952 9880
rect 347004 9868 347010 9920
rect 190178 9800 190184 9852
rect 190236 9840 190242 9852
rect 342898 9840 342904 9852
rect 190236 9812 342904 9840
rect 190236 9800 190242 9812
rect 342898 9800 342904 9812
rect 342956 9800 342962 9852
rect 188982 9732 188988 9784
rect 189040 9772 189046 9784
rect 339494 9772 339500 9784
rect 189040 9744 339500 9772
rect 189040 9732 189046 9744
rect 339494 9732 339500 9744
rect 339552 9732 339558 9784
rect 244918 9664 244924 9716
rect 244976 9704 244982 9716
rect 305546 9704 305552 9716
rect 244976 9676 305552 9704
rect 244976 9664 244982 9676
rect 305546 9664 305552 9676
rect 305604 9664 305610 9716
rect 157150 9596 157156 9648
rect 157208 9636 157214 9648
rect 273622 9636 273628 9648
rect 157208 9608 273628 9636
rect 157208 9596 157214 9608
rect 273622 9596 273628 9608
rect 273680 9596 273686 9648
rect 274450 9596 274456 9648
rect 274508 9636 274514 9648
rect 520734 9636 520740 9648
rect 274508 9608 520740 9636
rect 274508 9596 274514 9608
rect 520734 9596 520740 9608
rect 520792 9596 520798 9648
rect 158530 9528 158536 9580
rect 158588 9568 158594 9580
rect 277118 9568 277124 9580
rect 158588 9540 277124 9568
rect 158588 9528 158594 9540
rect 277118 9528 277124 9540
rect 277176 9528 277182 9580
rect 277210 9528 277216 9580
rect 277268 9568 277274 9580
rect 527818 9568 527824 9580
rect 277268 9540 527824 9568
rect 277268 9528 277274 9540
rect 527818 9528 527824 9540
rect 527876 9528 527882 9580
rect 160002 9460 160008 9512
rect 160060 9500 160066 9512
rect 279510 9500 279516 9512
rect 160060 9472 279516 9500
rect 160060 9460 160066 9472
rect 279510 9460 279516 9472
rect 279568 9460 279574 9512
rect 280706 9500 280712 9512
rect 279620 9472 280712 9500
rect 161198 9392 161204 9444
rect 161256 9432 161262 9444
rect 279620 9432 279648 9472
rect 280706 9460 280712 9472
rect 280764 9460 280770 9512
rect 282730 9460 282736 9512
rect 282788 9500 282794 9512
rect 286873 9503 286931 9509
rect 282788 9472 286824 9500
rect 282788 9460 282794 9472
rect 161256 9404 279648 9432
rect 161256 9392 161262 9404
rect 279970 9392 279976 9444
rect 280028 9432 280034 9444
rect 280028 9404 283328 9432
rect 280028 9392 280034 9404
rect 164142 9324 164148 9376
rect 164200 9364 164206 9376
rect 283193 9367 283251 9373
rect 283193 9364 283205 9367
rect 164200 9336 283205 9364
rect 164200 9324 164206 9336
rect 283193 9333 283205 9336
rect 283239 9333 283251 9367
rect 283193 9327 283251 9333
rect 161290 9256 161296 9308
rect 161348 9296 161354 9308
rect 283098 9296 283104 9308
rect 161348 9268 283104 9296
rect 161348 9256 161354 9268
rect 283098 9256 283104 9268
rect 283156 9256 283162 9308
rect 283300 9296 283328 9404
rect 284202 9392 284208 9444
rect 284260 9432 284266 9444
rect 286796 9432 286824 9472
rect 286873 9469 286885 9503
rect 286919 9500 286931 9503
rect 534902 9500 534908 9512
rect 286919 9472 534908 9500
rect 286919 9469 286931 9472
rect 286873 9463 286931 9469
rect 534902 9460 534908 9472
rect 534960 9460 534966 9512
rect 538398 9432 538404 9444
rect 284260 9404 286732 9432
rect 286796 9404 538404 9432
rect 284260 9392 284266 9404
rect 283377 9367 283435 9373
rect 283377 9333 283389 9367
rect 283423 9364 283435 9367
rect 286594 9364 286600 9376
rect 283423 9336 286600 9364
rect 283423 9333 283435 9336
rect 283377 9327 283435 9333
rect 286594 9324 286600 9336
rect 286652 9324 286658 9376
rect 286704 9364 286732 9404
rect 538398 9392 538404 9404
rect 538456 9392 538462 9444
rect 541986 9364 541992 9376
rect 286704 9336 541992 9364
rect 541986 9324 541992 9336
rect 542044 9324 542050 9376
rect 286781 9299 286839 9305
rect 286781 9296 286793 9299
rect 283300 9268 286793 9296
rect 286781 9265 286793 9268
rect 286827 9265 286839 9299
rect 286781 9259 286839 9265
rect 286870 9256 286876 9308
rect 286928 9296 286934 9308
rect 549070 9296 549076 9308
rect 286928 9268 549076 9296
rect 286928 9256 286934 9268
rect 549070 9256 549076 9268
rect 549128 9256 549134 9308
rect 165522 9188 165528 9240
rect 165580 9228 165586 9240
rect 290182 9228 290188 9240
rect 165580 9200 290188 9228
rect 165580 9188 165586 9200
rect 290182 9188 290188 9200
rect 290240 9188 290246 9240
rect 293770 9188 293776 9240
rect 293828 9228 293834 9240
rect 563238 9228 563244 9240
rect 293828 9200 563244 9228
rect 293828 9188 293834 9200
rect 563238 9188 563244 9200
rect 563296 9188 563302 9240
rect 166810 9120 166816 9172
rect 166868 9160 166874 9172
rect 293678 9160 293684 9172
rect 166868 9132 293684 9160
rect 166868 9120 166874 9132
rect 293678 9120 293684 9132
rect 293736 9120 293742 9172
rect 295150 9120 295156 9172
rect 295208 9160 295214 9172
rect 566826 9160 566832 9172
rect 295208 9132 566832 9160
rect 295208 9120 295214 9132
rect 566826 9120 566832 9132
rect 566884 9120 566890 9172
rect 173802 9052 173808 9104
rect 173860 9092 173866 9104
rect 307938 9092 307944 9104
rect 173860 9064 307944 9092
rect 173860 9052 173866 9064
rect 307938 9052 307944 9064
rect 307996 9052 308002 9104
rect 308398 9052 308404 9104
rect 308456 9092 308462 9104
rect 580994 9092 581000 9104
rect 308456 9064 581000 9092
rect 308456 9052 308462 9064
rect 580994 9052 581000 9064
rect 581052 9052 581058 9104
rect 168282 8984 168288 9036
rect 168340 9024 168346 9036
rect 297266 9024 297272 9036
rect 168340 8996 297272 9024
rect 168340 8984 168346 8996
rect 297266 8984 297272 8996
rect 297324 8984 297330 9036
rect 299290 8984 299296 9036
rect 299348 9024 299354 9036
rect 300581 9027 300639 9033
rect 300581 9024 300593 9027
rect 299348 8996 300593 9024
rect 299348 8984 299354 8996
rect 300581 8993 300593 8996
rect 300627 8993 300639 9027
rect 300581 8987 300639 8993
rect 300670 8984 300676 9036
rect 300728 9024 300734 9036
rect 300949 9027 301007 9033
rect 300728 8996 300900 9024
rect 300728 8984 300734 8996
rect 169662 8916 169668 8968
rect 169720 8956 169726 8968
rect 300762 8956 300768 8968
rect 169720 8928 300768 8956
rect 169720 8916 169726 8928
rect 300762 8916 300768 8928
rect 300820 8916 300826 8968
rect 300872 8956 300900 8996
rect 300949 8993 300961 9027
rect 300995 9024 301007 9027
rect 573910 9024 573916 9036
rect 300995 8996 573916 9024
rect 300995 8993 301007 8996
rect 300949 8987 301007 8993
rect 573910 8984 573916 8996
rect 573968 8984 573974 9036
rect 578602 8956 578608 8968
rect 300872 8928 578608 8956
rect 578602 8916 578608 8928
rect 578660 8916 578666 8968
rect 155678 8848 155684 8900
rect 155736 8888 155742 8900
rect 270034 8888 270040 8900
rect 155736 8860 270040 8888
rect 155736 8848 155742 8860
rect 270034 8848 270040 8860
rect 270092 8848 270098 8900
rect 270310 8848 270316 8900
rect 270368 8888 270374 8900
rect 513558 8888 513564 8900
rect 270368 8860 513564 8888
rect 270368 8848 270374 8860
rect 513558 8848 513564 8860
rect 513616 8848 513622 8900
rect 154390 8780 154396 8832
rect 154448 8820 154454 8832
rect 266538 8820 266544 8832
rect 154448 8792 266544 8820
rect 154448 8780 154454 8792
rect 266538 8780 266544 8792
rect 266596 8780 266602 8832
rect 267550 8780 267556 8832
rect 267608 8820 267614 8832
rect 506474 8820 506480 8832
rect 267608 8792 506480 8820
rect 267608 8780 267614 8792
rect 506474 8780 506480 8792
rect 506532 8780 506538 8832
rect 150158 8712 150164 8764
rect 150216 8752 150222 8764
rect 259454 8752 259460 8764
rect 150216 8724 259460 8752
rect 150216 8712 150222 8724
rect 259454 8712 259460 8724
rect 259512 8712 259518 8764
rect 262122 8712 262128 8764
rect 262180 8752 262186 8764
rect 262180 8724 263088 8752
rect 262180 8712 262186 8724
rect 152918 8644 152924 8696
rect 152976 8684 152982 8696
rect 262950 8684 262956 8696
rect 152976 8656 262956 8684
rect 152976 8644 152982 8656
rect 262950 8644 262956 8656
rect 263008 8644 263014 8696
rect 263060 8684 263088 8724
rect 263410 8712 263416 8764
rect 263468 8752 263474 8764
rect 499390 8752 499396 8764
rect 263468 8724 499396 8752
rect 263468 8712 263474 8724
rect 499390 8712 499396 8724
rect 499448 8712 499454 8764
rect 495894 8684 495900 8696
rect 263060 8656 495900 8684
rect 495894 8644 495900 8656
rect 495952 8644 495958 8696
rect 148870 8576 148876 8628
rect 148928 8616 148934 8628
rect 255866 8616 255872 8628
rect 148928 8588 255872 8616
rect 148928 8576 148934 8588
rect 255866 8576 255872 8588
rect 255924 8576 255930 8628
rect 259362 8576 259368 8628
rect 259420 8616 259426 8628
rect 488810 8616 488816 8628
rect 259420 8588 488816 8616
rect 259420 8576 259426 8588
rect 488810 8576 488816 8588
rect 488868 8576 488874 8628
rect 147398 8508 147404 8560
rect 147456 8548 147462 8560
rect 252370 8548 252376 8560
rect 147456 8520 252376 8548
rect 147456 8508 147462 8520
rect 252370 8508 252376 8520
rect 252428 8508 252434 8560
rect 256602 8508 256608 8560
rect 256660 8548 256666 8560
rect 485222 8548 485228 8560
rect 256660 8520 485228 8548
rect 256660 8508 256666 8520
rect 485222 8508 485228 8520
rect 485280 8508 485286 8560
rect 146110 8440 146116 8492
rect 146168 8480 146174 8492
rect 248782 8480 248788 8492
rect 146168 8452 248788 8480
rect 146168 8440 146174 8452
rect 248782 8440 248788 8452
rect 248840 8440 248846 8492
rect 255222 8440 255228 8492
rect 255280 8480 255286 8492
rect 481726 8480 481732 8492
rect 255280 8452 481732 8480
rect 255280 8440 255286 8452
rect 481726 8440 481732 8452
rect 481784 8440 481790 8492
rect 175182 8372 175188 8424
rect 175240 8412 175246 8424
rect 311434 8412 311440 8424
rect 175240 8384 311440 8412
rect 175240 8372 175246 8384
rect 311434 8372 311440 8384
rect 311492 8372 311498 8424
rect 172422 8304 172428 8356
rect 172480 8344 172486 8356
rect 304350 8344 304356 8356
rect 172480 8316 304356 8344
rect 172480 8304 172486 8316
rect 304350 8304 304356 8316
rect 304408 8304 304414 8356
rect 223482 8236 223488 8288
rect 223540 8276 223546 8288
rect 413094 8276 413100 8288
rect 223540 8248 413100 8276
rect 223540 8236 223546 8248
rect 413094 8236 413100 8248
rect 413152 8236 413158 8288
rect 123938 8168 123944 8220
rect 123996 8208 124002 8220
rect 201494 8208 201500 8220
rect 123996 8180 201500 8208
rect 123996 8168 124002 8180
rect 201494 8168 201500 8180
rect 201552 8168 201558 8220
rect 224770 8168 224776 8220
rect 224828 8208 224834 8220
rect 416682 8208 416688 8220
rect 224828 8180 416688 8208
rect 224828 8168 224834 8180
rect 416682 8168 416688 8180
rect 416740 8168 416746 8220
rect 125410 8100 125416 8152
rect 125468 8140 125474 8152
rect 205082 8140 205088 8152
rect 125468 8112 205088 8140
rect 125468 8100 125474 8112
rect 205082 8100 205088 8112
rect 205140 8100 205146 8152
rect 226242 8100 226248 8152
rect 226300 8140 226306 8152
rect 420178 8140 420184 8152
rect 226300 8112 420184 8140
rect 226300 8100 226306 8112
rect 420178 8100 420184 8112
rect 420236 8100 420242 8152
rect 126698 8032 126704 8084
rect 126756 8072 126762 8084
rect 208578 8072 208584 8084
rect 126756 8044 208584 8072
rect 126756 8032 126762 8044
rect 208578 8032 208584 8044
rect 208636 8032 208642 8084
rect 230290 8032 230296 8084
rect 230348 8072 230354 8084
rect 427262 8072 427268 8084
rect 230348 8044 427268 8072
rect 230348 8032 230354 8044
rect 427262 8032 427268 8044
rect 427320 8032 427326 8084
rect 132218 7964 132224 8016
rect 132276 8004 132282 8016
rect 219250 8004 219256 8016
rect 132276 7976 219256 8004
rect 132276 7964 132282 7976
rect 219250 7964 219256 7976
rect 219308 7964 219314 8016
rect 227530 7964 227536 8016
rect 227588 8004 227594 8016
rect 423766 8004 423772 8016
rect 227588 7976 423772 8004
rect 227588 7964 227594 7976
rect 423766 7964 423772 7976
rect 423824 7964 423830 8016
rect 129458 7896 129464 7948
rect 129516 7936 129522 7948
rect 215662 7936 215668 7948
rect 129516 7908 215668 7936
rect 129516 7896 129522 7908
rect 215662 7896 215668 7908
rect 215720 7896 215726 7948
rect 231762 7896 231768 7948
rect 231820 7936 231826 7948
rect 430850 7936 430856 7948
rect 231820 7908 430856 7936
rect 231820 7896 231826 7908
rect 430850 7896 430856 7908
rect 430908 7896 430914 7948
rect 133690 7828 133696 7880
rect 133748 7868 133754 7880
rect 222746 7868 222752 7880
rect 133748 7840 222752 7868
rect 133748 7828 133754 7840
rect 222746 7828 222752 7840
rect 222804 7828 222810 7880
rect 233142 7828 233148 7880
rect 233200 7868 233206 7880
rect 434438 7868 434444 7880
rect 233200 7840 434444 7868
rect 233200 7828 233206 7840
rect 434438 7828 434444 7840
rect 434496 7828 434502 7880
rect 134978 7760 134984 7812
rect 135036 7800 135042 7812
rect 226334 7800 226340 7812
rect 135036 7772 226340 7800
rect 135036 7760 135042 7772
rect 226334 7760 226340 7772
rect 226392 7760 226398 7812
rect 234522 7760 234528 7812
rect 234580 7800 234586 7812
rect 437934 7800 437940 7812
rect 234580 7772 437940 7800
rect 234580 7760 234586 7772
rect 437934 7760 437940 7772
rect 437992 7760 437998 7812
rect 139210 7692 139216 7744
rect 139268 7732 139274 7744
rect 234614 7732 234620 7744
rect 139268 7704 234620 7732
rect 139268 7692 139274 7704
rect 234614 7692 234620 7704
rect 234672 7692 234678 7744
rect 235902 7692 235908 7744
rect 235960 7732 235966 7744
rect 441522 7732 441528 7744
rect 235960 7704 441528 7732
rect 235960 7692 235966 7704
rect 441522 7692 441528 7704
rect 441580 7692 441586 7744
rect 141970 7624 141976 7676
rect 142028 7664 142034 7676
rect 241698 7664 241704 7676
rect 142028 7636 241704 7664
rect 142028 7624 142034 7636
rect 241698 7624 241704 7636
rect 241756 7624 241762 7676
rect 242802 7624 242808 7676
rect 242860 7664 242866 7676
rect 455690 7664 455696 7676
rect 242860 7636 455696 7664
rect 242860 7624 242866 7636
rect 455690 7624 455696 7636
rect 455748 7624 455754 7676
rect 143258 7556 143264 7608
rect 143316 7596 143322 7608
rect 245194 7596 245200 7608
rect 143316 7568 245200 7596
rect 143316 7556 143322 7568
rect 245194 7556 245200 7568
rect 245252 7556 245258 7608
rect 245562 7556 245568 7608
rect 245620 7596 245626 7608
rect 459186 7596 459192 7608
rect 245620 7568 459192 7596
rect 245620 7556 245626 7568
rect 459186 7556 459192 7568
rect 459244 7556 459250 7608
rect 222102 7488 222108 7540
rect 222160 7528 222166 7540
rect 409598 7528 409604 7540
rect 222160 7500 409604 7528
rect 222160 7488 222166 7500
rect 409598 7488 409604 7500
rect 409656 7488 409662 7540
rect 219342 7420 219348 7472
rect 219400 7460 219406 7472
rect 406010 7460 406016 7472
rect 219400 7432 406016 7460
rect 219400 7420 219406 7432
rect 406010 7420 406016 7432
rect 406068 7420 406074 7472
rect 217870 7352 217876 7404
rect 217928 7392 217934 7404
rect 402514 7392 402520 7404
rect 217928 7364 402520 7392
rect 217928 7352 217934 7364
rect 402514 7352 402520 7364
rect 402572 7352 402578 7404
rect 216582 7284 216588 7336
rect 216640 7324 216646 7336
rect 398926 7324 398932 7336
rect 216640 7296 398932 7324
rect 216640 7284 216646 7296
rect 398926 7284 398932 7296
rect 398984 7284 398990 7336
rect 215202 7216 215208 7268
rect 215260 7256 215266 7268
rect 395338 7256 395344 7268
rect 215260 7228 395344 7256
rect 215260 7216 215266 7228
rect 395338 7216 395344 7228
rect 395396 7216 395402 7268
rect 213730 7148 213736 7200
rect 213788 7188 213794 7200
rect 391842 7188 391848 7200
rect 213788 7160 391848 7188
rect 213788 7148 213794 7160
rect 391842 7148 391848 7160
rect 391900 7148 391906 7200
rect 210970 7080 210976 7132
rect 211028 7120 211034 7132
rect 388254 7120 388260 7132
rect 211028 7092 388260 7120
rect 211028 7080 211034 7092
rect 388254 7080 388260 7092
rect 388312 7080 388318 7132
rect 209682 7012 209688 7064
rect 209740 7052 209746 7064
rect 384758 7052 384764 7064
rect 209740 7024 384764 7052
rect 209740 7012 209746 7024
rect 384758 7012 384764 7024
rect 384816 7012 384822 7064
rect 158622 6944 158628 6996
rect 158680 6984 158686 6996
rect 276014 6984 276020 6996
rect 158680 6956 276020 6984
rect 158680 6944 158686 6956
rect 276014 6944 276020 6956
rect 276072 6944 276078 6996
rect 276658 6944 276664 6996
rect 276716 6984 276722 6996
rect 319714 6984 319720 6996
rect 276716 6956 319720 6984
rect 276716 6944 276722 6956
rect 319714 6944 319720 6956
rect 319772 6944 319778 6996
rect 142062 6808 142068 6860
rect 142120 6848 142126 6860
rect 240502 6848 240508 6860
rect 142120 6820 240508 6848
rect 142120 6808 142126 6820
rect 240502 6808 240508 6820
rect 240560 6808 240566 6860
rect 242158 6808 242164 6860
rect 242216 6848 242222 6860
rect 301406 6848 301412 6860
rect 242216 6820 301412 6848
rect 242216 6808 242222 6820
rect 301406 6808 301412 6820
rect 301464 6808 301470 6860
rect 301498 6808 301504 6860
rect 301556 6848 301562 6860
rect 312630 6848 312636 6860
rect 301556 6820 312636 6848
rect 301556 6808 301562 6820
rect 312630 6808 312636 6820
rect 312688 6808 312694 6860
rect 315298 6808 315304 6860
rect 315356 6848 315362 6860
rect 580166 6848 580172 6860
rect 315356 6820 580172 6848
rect 315356 6808 315362 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 117130 6740 117136 6792
rect 117188 6780 117194 6792
rect 187326 6780 187332 6792
rect 117188 6752 187332 6780
rect 117188 6740 117194 6752
rect 187326 6740 187332 6752
rect 187384 6740 187390 6792
rect 198642 6740 198648 6792
rect 198700 6780 198706 6792
rect 359918 6780 359924 6792
rect 198700 6752 359924 6780
rect 198700 6740 198706 6752
rect 359918 6740 359924 6752
rect 359976 6740 359982 6792
rect 118510 6672 118516 6724
rect 118568 6712 118574 6724
rect 190822 6712 190828 6724
rect 118568 6684 190828 6712
rect 118568 6672 118574 6684
rect 190822 6672 190828 6684
rect 190880 6672 190886 6724
rect 200022 6672 200028 6724
rect 200080 6712 200086 6724
rect 363506 6712 363512 6724
rect 200080 6684 363512 6712
rect 200080 6672 200086 6684
rect 363506 6672 363512 6684
rect 363564 6672 363570 6724
rect 119982 6604 119988 6656
rect 120040 6644 120046 6656
rect 194318 6644 194324 6656
rect 120040 6616 194324 6644
rect 120040 6604 120046 6616
rect 194318 6604 194324 6616
rect 194376 6604 194382 6656
rect 201310 6604 201316 6656
rect 201368 6644 201374 6656
rect 367002 6644 367008 6656
rect 201368 6616 367008 6644
rect 201368 6604 201374 6616
rect 367002 6604 367008 6616
rect 367060 6604 367066 6656
rect 121270 6536 121276 6588
rect 121328 6576 121334 6588
rect 197906 6576 197912 6588
rect 121328 6548 197912 6576
rect 121328 6536 121334 6548
rect 197906 6536 197912 6548
rect 197964 6536 197970 6588
rect 237190 6536 237196 6588
rect 237248 6576 237254 6588
rect 442626 6576 442632 6588
rect 237248 6548 442632 6576
rect 237248 6536 237254 6548
rect 442626 6536 442632 6548
rect 442684 6536 442690 6588
rect 143350 6468 143356 6520
rect 143408 6508 143414 6520
rect 244090 6508 244096 6520
rect 143408 6480 244096 6508
rect 143408 6468 143414 6480
rect 244090 6468 244096 6480
rect 244148 6468 244154 6520
rect 260742 6468 260748 6520
rect 260800 6508 260806 6520
rect 492306 6508 492312 6520
rect 260800 6480 492312 6508
rect 260800 6468 260806 6480
rect 492306 6468 492312 6480
rect 492364 6468 492370 6520
rect 144730 6400 144736 6452
rect 144788 6440 144794 6452
rect 247586 6440 247592 6452
rect 144788 6412 247592 6440
rect 144788 6400 144794 6412
rect 247586 6400 247592 6412
rect 247644 6400 247650 6452
rect 264790 6400 264796 6452
rect 264848 6440 264854 6452
rect 502978 6440 502984 6452
rect 264848 6412 502984 6440
rect 264848 6400 264854 6412
rect 502978 6400 502984 6412
rect 503036 6400 503042 6452
rect 147490 6332 147496 6384
rect 147548 6372 147554 6384
rect 251174 6372 251180 6384
rect 147548 6344 251180 6372
rect 147548 6332 147554 6344
rect 251174 6332 251180 6344
rect 251232 6332 251238 6384
rect 269022 6332 269028 6384
rect 269080 6372 269086 6384
rect 510062 6372 510068 6384
rect 269080 6344 510068 6372
rect 269080 6332 269086 6344
rect 510062 6332 510068 6344
rect 510120 6332 510126 6384
rect 99190 6264 99196 6316
rect 99248 6304 99254 6316
rect 150618 6304 150624 6316
rect 99248 6276 150624 6304
rect 99248 6264 99254 6276
rect 150618 6264 150624 6276
rect 150676 6264 150682 6316
rect 151630 6264 151636 6316
rect 151688 6304 151694 6316
rect 261754 6304 261760 6316
rect 151688 6276 261760 6304
rect 151688 6264 151694 6276
rect 261754 6264 261760 6276
rect 261812 6264 261818 6316
rect 271690 6264 271696 6316
rect 271748 6304 271754 6316
rect 517146 6304 517152 6316
rect 271748 6276 517152 6304
rect 271748 6264 271754 6276
rect 517146 6264 517152 6276
rect 517204 6264 517210 6316
rect 100478 6196 100484 6248
rect 100536 6236 100542 6248
rect 154206 6236 154212 6248
rect 100536 6208 154212 6236
rect 100536 6196 100542 6208
rect 154206 6196 154212 6208
rect 154264 6196 154270 6248
rect 155770 6196 155776 6248
rect 155828 6236 155834 6248
rect 268838 6236 268844 6248
rect 155828 6208 268844 6236
rect 155828 6196 155834 6208
rect 268838 6196 268844 6208
rect 268896 6196 268902 6248
rect 275922 6196 275928 6248
rect 275980 6236 275986 6248
rect 524230 6236 524236 6248
rect 275980 6208 524236 6236
rect 275980 6196 275986 6208
rect 524230 6196 524236 6208
rect 524288 6196 524294 6248
rect 111610 6128 111616 6180
rect 111668 6168 111674 6180
rect 176654 6168 176660 6180
rect 111668 6140 176660 6168
rect 111668 6128 111674 6140
rect 176654 6128 176660 6140
rect 176712 6128 176718 6180
rect 179322 6128 179328 6180
rect 179380 6168 179386 6180
rect 320910 6168 320916 6180
rect 179380 6140 320916 6168
rect 179380 6128 179386 6140
rect 320910 6128 320916 6140
rect 320968 6128 320974 6180
rect 322198 6128 322204 6180
rect 322256 6168 322262 6180
rect 583389 6171 583447 6177
rect 583389 6168 583401 6171
rect 322256 6140 583401 6168
rect 322256 6128 322262 6140
rect 583389 6137 583401 6140
rect 583435 6137 583447 6171
rect 583389 6131 583447 6137
rect 115750 6060 115756 6112
rect 115808 6100 115814 6112
rect 183738 6100 183744 6112
rect 115808 6072 183744 6100
rect 115808 6060 115814 6072
rect 183738 6060 183744 6072
rect 183796 6060 183802 6112
rect 194410 6060 194416 6112
rect 194468 6100 194474 6112
rect 352834 6100 352840 6112
rect 194468 6072 352840 6100
rect 194468 6060 194474 6072
rect 352834 6060 352840 6072
rect 352892 6060 352898 6112
rect 113082 5992 113088 6044
rect 113140 6032 113146 6044
rect 180242 6032 180248 6044
rect 113140 6004 180248 6032
rect 113140 5992 113146 6004
rect 180242 5992 180248 6004
rect 180300 5992 180306 6044
rect 193122 5992 193128 6044
rect 193180 6032 193186 6044
rect 349246 6032 349252 6044
rect 193180 6004 349252 6032
rect 193180 5992 193186 6004
rect 349246 5992 349252 6004
rect 349304 5992 349310 6044
rect 114462 5924 114468 5976
rect 114520 5964 114526 5976
rect 181438 5964 181444 5976
rect 114520 5936 181444 5964
rect 114520 5924 114526 5936
rect 181438 5924 181444 5936
rect 181496 5924 181502 5976
rect 191742 5924 191748 5976
rect 191800 5964 191806 5976
rect 345750 5964 345756 5976
rect 191800 5936 345756 5964
rect 191800 5924 191806 5936
rect 345750 5924 345756 5936
rect 345808 5924 345814 5976
rect 110230 5856 110236 5908
rect 110288 5896 110294 5908
rect 173158 5896 173164 5908
rect 110288 5868 173164 5896
rect 110288 5856 110294 5868
rect 173158 5856 173164 5868
rect 173216 5856 173222 5908
rect 190270 5856 190276 5908
rect 190328 5896 190334 5908
rect 342162 5896 342168 5908
rect 190328 5868 342168 5896
rect 190328 5856 190334 5868
rect 342162 5856 342168 5868
rect 342220 5856 342226 5908
rect 108942 5788 108948 5840
rect 109000 5828 109006 5840
rect 170766 5828 170772 5840
rect 109000 5800 170772 5828
rect 109000 5788 109006 5800
rect 170766 5788 170772 5800
rect 170824 5788 170830 5840
rect 187510 5788 187516 5840
rect 187568 5828 187574 5840
rect 338666 5828 338672 5840
rect 187568 5800 338672 5828
rect 187568 5788 187574 5800
rect 338666 5788 338672 5800
rect 338724 5788 338730 5840
rect 108850 5720 108856 5772
rect 108908 5760 108914 5772
rect 169570 5760 169576 5772
rect 108908 5732 169576 5760
rect 108908 5720 108914 5732
rect 169570 5720 169576 5732
rect 169628 5720 169634 5772
rect 186222 5720 186228 5772
rect 186280 5760 186286 5772
rect 335078 5760 335084 5772
rect 186280 5732 335084 5760
rect 186280 5720 186286 5732
rect 335078 5720 335084 5732
rect 335136 5720 335142 5772
rect 106090 5652 106096 5704
rect 106148 5692 106154 5704
rect 166074 5692 166080 5704
rect 106148 5664 166080 5692
rect 106148 5652 106154 5664
rect 166074 5652 166080 5664
rect 166132 5652 166138 5704
rect 184750 5652 184756 5704
rect 184808 5692 184814 5704
rect 331582 5692 331588 5704
rect 184808 5664 331588 5692
rect 184808 5652 184814 5664
rect 331582 5652 331588 5664
rect 331640 5652 331646 5704
rect 104802 5584 104808 5636
rect 104860 5624 104866 5636
rect 162486 5624 162492 5636
rect 104860 5596 162492 5624
rect 104860 5584 104866 5596
rect 162486 5584 162492 5596
rect 162544 5584 162550 5636
rect 183462 5584 183468 5636
rect 183520 5624 183526 5636
rect 327994 5624 328000 5636
rect 183520 5596 328000 5624
rect 183520 5584 183526 5596
rect 327994 5584 328000 5596
rect 328052 5584 328058 5636
rect 103238 5516 103244 5568
rect 103296 5556 103302 5568
rect 157794 5556 157800 5568
rect 103296 5528 157800 5556
rect 103296 5516 103302 5528
rect 157794 5516 157800 5528
rect 157852 5516 157858 5568
rect 182082 5516 182088 5568
rect 182140 5556 182146 5568
rect 324406 5556 324412 5568
rect 182140 5528 324412 5556
rect 182140 5516 182146 5528
rect 324406 5516 324412 5528
rect 324464 5516 324470 5568
rect 93762 5448 93768 5500
rect 93820 5488 93826 5500
rect 137646 5488 137652 5500
rect 93820 5460 137652 5488
rect 93820 5448 93826 5460
rect 137646 5448 137652 5460
rect 137704 5448 137710 5500
rect 137830 5448 137836 5500
rect 137888 5488 137894 5500
rect 232222 5488 232228 5500
rect 137888 5460 232228 5488
rect 137888 5448 137894 5460
rect 232222 5448 232228 5460
rect 232280 5448 232286 5500
rect 278682 5448 278688 5500
rect 278740 5488 278746 5500
rect 530118 5488 530124 5500
rect 278740 5460 530124 5488
rect 278740 5448 278746 5460
rect 530118 5448 530124 5460
rect 530176 5448 530182 5500
rect 94958 5380 94964 5432
rect 95016 5420 95022 5432
rect 140038 5420 140044 5432
rect 95016 5392 140044 5420
rect 95016 5380 95022 5392
rect 140038 5380 140044 5392
rect 140096 5380 140102 5432
rect 140590 5380 140596 5432
rect 140648 5420 140654 5432
rect 239306 5420 239312 5432
rect 140648 5392 239312 5420
rect 140648 5380 140654 5392
rect 239306 5380 239312 5392
rect 239364 5380 239370 5432
rect 274542 5380 274548 5432
rect 274600 5420 274606 5432
rect 278501 5423 278559 5429
rect 278501 5420 278513 5423
rect 274600 5392 278513 5420
rect 274600 5380 274606 5392
rect 278501 5389 278513 5392
rect 278547 5389 278559 5423
rect 278501 5383 278559 5389
rect 280062 5380 280068 5432
rect 280120 5420 280126 5432
rect 533706 5420 533712 5432
rect 280120 5392 533712 5420
rect 280120 5380 280126 5392
rect 533706 5380 533712 5392
rect 533764 5380 533770 5432
rect 95050 5312 95056 5364
rect 95108 5352 95114 5364
rect 141234 5352 141240 5364
rect 95108 5324 141240 5352
rect 95108 5312 95114 5324
rect 141234 5312 141240 5324
rect 141292 5312 141298 5364
rect 143442 5312 143448 5364
rect 143500 5352 143506 5364
rect 242894 5352 242900 5364
rect 143500 5324 242900 5352
rect 143500 5312 143506 5324
rect 242894 5312 242900 5324
rect 242952 5312 242958 5364
rect 277302 5312 277308 5364
rect 277360 5352 277366 5364
rect 278317 5355 278375 5361
rect 278317 5352 278329 5355
rect 277360 5324 278329 5352
rect 277360 5312 277366 5324
rect 278317 5321 278329 5324
rect 278363 5321 278375 5355
rect 278317 5315 278375 5321
rect 282822 5312 282828 5364
rect 282880 5352 282886 5364
rect 291933 5355 291991 5361
rect 282880 5324 291884 5352
rect 282880 5312 282886 5324
rect 96522 5244 96528 5296
rect 96580 5284 96586 5296
rect 144730 5284 144736 5296
rect 96580 5256 144736 5284
rect 96580 5244 96586 5256
rect 144730 5244 144736 5256
rect 144788 5244 144794 5296
rect 144822 5244 144828 5296
rect 144880 5284 144886 5296
rect 246390 5284 246396 5296
rect 144880 5256 246396 5284
rect 144880 5244 144886 5256
rect 246390 5244 246396 5256
rect 246448 5244 246454 5296
rect 277857 5287 277915 5293
rect 277857 5253 277869 5287
rect 277903 5284 277915 5287
rect 284294 5284 284300 5296
rect 277903 5256 284300 5284
rect 277903 5253 277915 5256
rect 277857 5247 277915 5253
rect 284294 5244 284300 5256
rect 284352 5244 284358 5296
rect 285582 5244 285588 5296
rect 285640 5284 285646 5296
rect 291856 5284 291884 5324
rect 291933 5321 291945 5355
rect 291979 5352 291991 5355
rect 537202 5352 537208 5364
rect 291979 5324 537208 5352
rect 291979 5321 291991 5324
rect 291933 5315 291991 5321
rect 537202 5312 537208 5324
rect 537260 5312 537266 5364
rect 540790 5284 540796 5296
rect 285640 5256 291792 5284
rect 291856 5256 540796 5284
rect 285640 5244 285646 5256
rect 96430 5176 96436 5228
rect 96488 5216 96494 5228
rect 143534 5216 143540 5228
rect 96488 5188 143540 5216
rect 96488 5176 96494 5188
rect 143534 5176 143540 5188
rect 143592 5176 143598 5228
rect 146202 5176 146208 5228
rect 146260 5216 146266 5228
rect 249978 5216 249984 5228
rect 146260 5188 249984 5216
rect 146260 5176 146266 5188
rect 249978 5176 249984 5188
rect 250036 5176 250042 5228
rect 277581 5219 277639 5225
rect 277581 5185 277593 5219
rect 277627 5216 277639 5219
rect 281902 5216 281908 5228
rect 277627 5188 281908 5216
rect 277627 5185 277639 5188
rect 277581 5179 277639 5185
rect 281902 5176 281908 5188
rect 281960 5176 281966 5228
rect 288342 5176 288348 5228
rect 288400 5216 288406 5228
rect 291654 5216 291660 5228
rect 288400 5188 291660 5216
rect 288400 5176 288406 5188
rect 291654 5176 291660 5188
rect 291712 5176 291718 5228
rect 291764 5216 291792 5256
rect 540790 5244 540796 5256
rect 540848 5244 540854 5296
rect 544378 5216 544384 5228
rect 291764 5188 544384 5216
rect 544378 5176 544384 5188
rect 544436 5176 544442 5228
rect 97810 5108 97816 5160
rect 97868 5148 97874 5160
rect 147122 5148 147128 5160
rect 97868 5120 147128 5148
rect 97868 5108 97874 5120
rect 147122 5108 147128 5120
rect 147180 5108 147186 5160
rect 147582 5108 147588 5160
rect 147640 5148 147646 5160
rect 253474 5148 253480 5160
rect 147640 5120 253480 5148
rect 147640 5108 147646 5120
rect 253474 5108 253480 5120
rect 253532 5108 253538 5160
rect 271782 5108 271788 5160
rect 271840 5148 271846 5160
rect 278041 5151 278099 5157
rect 278041 5148 278053 5151
rect 271840 5120 278053 5148
rect 271840 5108 271846 5120
rect 278041 5117 278053 5120
rect 278087 5117 278099 5151
rect 278041 5111 278099 5117
rect 286962 5108 286968 5160
rect 287020 5148 287026 5160
rect 547874 5148 547880 5160
rect 287020 5120 547880 5148
rect 287020 5108 287026 5120
rect 547874 5108 547880 5120
rect 547932 5108 547938 5160
rect 97718 5040 97724 5092
rect 97776 5080 97782 5092
rect 148318 5080 148324 5092
rect 97776 5052 148324 5080
rect 97776 5040 97782 5052
rect 148318 5040 148324 5052
rect 148376 5040 148382 5092
rect 150342 5040 150348 5092
rect 150400 5080 150406 5092
rect 257062 5080 257068 5092
rect 150400 5052 257068 5080
rect 150400 5040 150406 5052
rect 257062 5040 257068 5052
rect 257120 5040 257126 5092
rect 264882 5040 264888 5092
rect 264940 5080 264946 5092
rect 268657 5083 268715 5089
rect 268657 5080 268669 5083
rect 264940 5052 268669 5080
rect 264940 5040 264946 5052
rect 268657 5049 268669 5052
rect 268703 5049 268715 5083
rect 268657 5043 268715 5049
rect 273162 5040 273168 5092
rect 273220 5080 273226 5092
rect 277949 5083 278007 5089
rect 273220 5040 273254 5080
rect 277949 5049 277961 5083
rect 277995 5080 278007 5083
rect 277995 5052 291884 5080
rect 277995 5049 278007 5052
rect 277949 5043 278007 5049
rect 100570 4972 100576 5024
rect 100628 5012 100634 5024
rect 151814 5012 151820 5024
rect 100628 4984 151820 5012
rect 100628 4972 100634 4984
rect 151814 4972 151820 4984
rect 151872 4972 151878 5024
rect 153102 4972 153108 5024
rect 153160 5012 153166 5024
rect 264146 5012 264152 5024
rect 153160 4984 264152 5012
rect 153160 4972 153166 4984
rect 264146 4972 264152 4984
rect 264204 4972 264210 5024
rect 266262 4972 266268 5024
rect 266320 5012 266326 5024
rect 268565 5015 268623 5021
rect 268565 5012 268577 5015
rect 266320 4984 268577 5012
rect 266320 4972 266326 4984
rect 268565 4981 268577 4984
rect 268611 4981 268623 5015
rect 273226 5012 273254 5040
rect 278225 5015 278283 5021
rect 278225 5012 278237 5015
rect 273226 4984 278237 5012
rect 268565 4975 268623 4981
rect 278225 4981 278237 4984
rect 278271 4981 278283 5015
rect 278225 4975 278283 4981
rect 281442 4972 281448 5024
rect 281500 5012 281506 5024
rect 291749 5015 291807 5021
rect 291749 5012 291761 5015
rect 281500 4984 291761 5012
rect 281500 4972 281506 4984
rect 291749 4981 291761 4984
rect 291795 4981 291807 5015
rect 291749 4975 291807 4981
rect 102042 4904 102048 4956
rect 102100 4944 102106 4956
rect 155402 4944 155408 4956
rect 102100 4916 155408 4944
rect 102100 4904 102106 4916
rect 155402 4904 155408 4916
rect 155460 4904 155466 4956
rect 155862 4904 155868 4956
rect 155920 4944 155926 4956
rect 271230 4944 271236 4956
rect 155920 4916 271236 4944
rect 155920 4904 155926 4916
rect 271230 4904 271236 4916
rect 271288 4904 271294 4956
rect 277305 4947 277363 4953
rect 277305 4913 277317 4947
rect 277351 4944 277363 4947
rect 291856 4944 291884 5052
rect 291930 5040 291936 5092
rect 291988 5080 291994 5092
rect 551462 5080 551468 5092
rect 291988 5052 551468 5080
rect 291988 5040 291994 5052
rect 551462 5040 551468 5052
rect 551520 5040 551526 5092
rect 295242 4972 295248 5024
rect 295300 5012 295306 5024
rect 301593 5015 301651 5021
rect 295300 4984 301544 5012
rect 295300 4972 295306 4984
rect 298462 4944 298468 4956
rect 277351 4916 291792 4944
rect 291856 4916 298468 4944
rect 277351 4913 277363 4916
rect 277305 4907 277363 4913
rect 103330 4836 103336 4888
rect 103388 4876 103394 4888
rect 158898 4876 158904 4888
rect 103388 4848 158904 4876
rect 103388 4836 103394 4848
rect 158898 4836 158904 4848
rect 158956 4836 158962 4888
rect 161382 4836 161388 4888
rect 161440 4876 161446 4888
rect 277581 4879 277639 4885
rect 277581 4876 277593 4879
rect 161440 4848 277593 4876
rect 161440 4836 161446 4848
rect 277581 4845 277593 4848
rect 277627 4845 277639 4879
rect 277581 4839 277639 4845
rect 278133 4879 278191 4885
rect 278133 4845 278145 4879
rect 278179 4876 278191 4879
rect 291378 4876 291384 4888
rect 278179 4848 291384 4876
rect 278179 4845 278191 4848
rect 278133 4839 278191 4845
rect 291378 4836 291384 4848
rect 291436 4836 291442 4888
rect 291764 4876 291792 4916
rect 298462 4904 298468 4916
rect 298520 4904 298526 4956
rect 299382 4904 299388 4956
rect 299440 4944 299446 4956
rect 301409 4947 301467 4953
rect 301409 4944 301421 4947
rect 299440 4916 301421 4944
rect 299440 4904 299446 4916
rect 301409 4913 301421 4916
rect 301455 4913 301467 4947
rect 301516 4944 301544 4984
rect 301593 4981 301605 5015
rect 301639 5012 301651 5015
rect 562042 5012 562048 5024
rect 301639 4984 562048 5012
rect 301639 4981 301651 4984
rect 301593 4975 301651 4981
rect 562042 4972 562048 4984
rect 562100 4972 562106 5024
rect 565630 4944 565636 4956
rect 301516 4916 565636 4944
rect 301409 4907 301467 4913
rect 565630 4904 565636 4916
rect 565688 4904 565694 4956
rect 294874 4876 294880 4888
rect 291764 4848 294880 4876
rect 294874 4836 294880 4848
rect 294932 4836 294938 4888
rect 296622 4836 296628 4888
rect 296680 4876 296686 4888
rect 569126 4876 569132 4888
rect 296680 4848 569132 4876
rect 296680 4836 296686 4848
rect 569126 4836 569132 4848
rect 569184 4836 569190 4888
rect 106182 4768 106188 4820
rect 106240 4808 106246 4820
rect 163682 4808 163688 4820
rect 106240 4780 163688 4808
rect 106240 4768 106246 4780
rect 163682 4768 163688 4780
rect 163740 4768 163746 4820
rect 166902 4768 166908 4820
rect 166960 4808 166966 4820
rect 292574 4808 292580 4820
rect 166960 4780 278084 4808
rect 166960 4768 166966 4780
rect 92290 4700 92296 4752
rect 92348 4740 92354 4752
rect 134150 4740 134156 4752
rect 92348 4712 134156 4740
rect 92348 4700 92354 4712
rect 134150 4700 134156 4712
rect 134208 4700 134214 4752
rect 136542 4700 136548 4752
rect 136600 4740 136606 4752
rect 228726 4740 228732 4752
rect 136600 4712 228732 4740
rect 136600 4700 136606 4712
rect 228726 4700 228732 4712
rect 228784 4700 228790 4752
rect 268381 4743 268439 4749
rect 268381 4709 268393 4743
rect 268427 4740 268439 4743
rect 277949 4743 278007 4749
rect 277949 4740 277961 4743
rect 268427 4712 277961 4740
rect 268427 4709 268439 4712
rect 268381 4703 268439 4709
rect 277949 4709 277961 4712
rect 277995 4709 278007 4743
rect 278056 4740 278084 4780
rect 278424 4780 292580 4808
rect 278424 4740 278452 4780
rect 292574 4768 292580 4780
rect 292632 4768 292638 4820
rect 293862 4768 293868 4820
rect 293920 4808 293926 4820
rect 301593 4811 301651 4817
rect 301593 4808 301605 4811
rect 293920 4780 301605 4808
rect 293920 4768 293926 4780
rect 301593 4777 301605 4780
rect 301639 4777 301651 4811
rect 301593 4771 301651 4777
rect 301685 4811 301743 4817
rect 301685 4777 301697 4811
rect 301731 4808 301743 4811
rect 576302 4808 576308 4820
rect 301731 4780 576308 4808
rect 301731 4777 301743 4780
rect 301685 4771 301743 4777
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 278056 4712 278452 4740
rect 278501 4743 278559 4749
rect 277949 4703 278007 4709
rect 278501 4709 278513 4743
rect 278547 4740 278559 4743
rect 523034 4740 523040 4752
rect 278547 4712 523040 4740
rect 278547 4709 278559 4712
rect 278501 4703 278559 4709
rect 523034 4700 523040 4712
rect 523092 4700 523098 4752
rect 89622 4632 89628 4684
rect 89680 4672 89686 4684
rect 129366 4672 129372 4684
rect 89680 4644 129372 4672
rect 89680 4632 89686 4644
rect 129366 4632 129372 4644
rect 129424 4632 129430 4684
rect 135070 4632 135076 4684
rect 135128 4672 135134 4684
rect 225138 4672 225144 4684
rect 135128 4644 225144 4672
rect 135128 4632 135134 4644
rect 225138 4632 225144 4644
rect 225196 4632 225202 4684
rect 263502 4632 263508 4684
rect 263560 4672 263566 4684
rect 268197 4675 268255 4681
rect 268197 4672 268209 4675
rect 263560 4644 268209 4672
rect 263560 4632 263566 4644
rect 268197 4641 268209 4644
rect 268243 4641 268255 4675
rect 268197 4635 268255 4641
rect 268289 4675 268347 4681
rect 268289 4641 268301 4675
rect 268335 4672 268347 4675
rect 277305 4675 277363 4681
rect 277305 4672 277317 4675
rect 268335 4644 277317 4672
rect 268335 4641 268347 4644
rect 268289 4635 268347 4641
rect 277305 4641 277317 4644
rect 277351 4641 277363 4675
rect 277305 4635 277363 4641
rect 278317 4675 278375 4681
rect 278317 4641 278329 4675
rect 278363 4672 278375 4675
rect 526622 4672 526628 4684
rect 278363 4644 526628 4672
rect 278363 4641 278375 4644
rect 278317 4635 278375 4641
rect 526622 4632 526628 4644
rect 526680 4632 526686 4684
rect 88242 4564 88248 4616
rect 88300 4604 88306 4616
rect 125870 4604 125876 4616
rect 88300 4576 125876 4604
rect 88300 4564 88306 4576
rect 125870 4564 125876 4576
rect 125928 4564 125934 4616
rect 132310 4564 132316 4616
rect 132368 4604 132374 4616
rect 221550 4604 221556 4616
rect 132368 4576 221556 4604
rect 132368 4564 132374 4576
rect 221550 4564 221556 4576
rect 221608 4564 221614 4616
rect 278133 4607 278191 4613
rect 278133 4604 278145 4607
rect 263566 4576 278145 4604
rect 130930 4496 130936 4548
rect 130988 4536 130994 4548
rect 218054 4536 218060 4548
rect 130988 4508 218060 4536
rect 130988 4496 130994 4508
rect 218054 4496 218060 4508
rect 218112 4496 218118 4548
rect 124030 4428 124036 4480
rect 124088 4468 124094 4480
rect 203886 4468 203892 4480
rect 124088 4440 203892 4468
rect 124088 4428 124094 4440
rect 203886 4428 203892 4440
rect 203944 4428 203950 4480
rect 204898 4428 204904 4480
rect 204956 4468 204962 4480
rect 263566 4468 263594 4576
rect 278133 4573 278145 4576
rect 278179 4573 278191 4607
rect 278133 4567 278191 4573
rect 278225 4607 278283 4613
rect 278225 4573 278237 4607
rect 278271 4604 278283 4607
rect 519538 4604 519544 4616
rect 278271 4576 519544 4604
rect 278271 4573 278283 4576
rect 278225 4567 278283 4573
rect 519538 4564 519544 4576
rect 519596 4564 519602 4616
rect 268473 4539 268531 4545
rect 268473 4505 268485 4539
rect 268519 4536 268531 4539
rect 277857 4539 277915 4545
rect 277857 4536 277869 4539
rect 268519 4508 277869 4536
rect 268519 4505 268531 4508
rect 268473 4499 268531 4505
rect 277857 4505 277869 4508
rect 277903 4505 277915 4539
rect 277857 4499 277915 4505
rect 278041 4539 278099 4545
rect 278041 4505 278053 4539
rect 278087 4536 278099 4539
rect 515950 4536 515956 4548
rect 278087 4508 515956 4536
rect 278087 4505 278099 4508
rect 278041 4499 278099 4505
rect 515950 4496 515956 4508
rect 516008 4496 516014 4548
rect 204956 4440 263594 4468
rect 204956 4428 204962 4440
rect 267642 4428 267648 4480
rect 267700 4468 267706 4480
rect 267700 4440 268608 4468
rect 267700 4428 267706 4440
rect 128262 4360 128268 4412
rect 128320 4400 128326 4412
rect 210970 4400 210976 4412
rect 128320 4372 210976 4400
rect 128320 4360 128326 4372
rect 210970 4360 210976 4372
rect 211028 4360 211034 4412
rect 213178 4360 213184 4412
rect 213236 4400 213242 4412
rect 268381 4403 268439 4409
rect 268381 4400 268393 4403
rect 213236 4372 268393 4400
rect 213236 4360 213242 4372
rect 268381 4369 268393 4372
rect 268427 4369 268439 4403
rect 268580 4400 268608 4440
rect 270402 4428 270408 4480
rect 270460 4468 270466 4480
rect 512454 4468 512460 4480
rect 270460 4440 512460 4468
rect 270460 4428 270466 4440
rect 512454 4428 512460 4440
rect 512512 4428 512518 4480
rect 508866 4400 508872 4412
rect 268580 4372 508872 4400
rect 268381 4363 268439 4369
rect 508866 4360 508872 4372
rect 508924 4360 508930 4412
rect 126790 4292 126796 4344
rect 126848 4332 126854 4344
rect 207382 4332 207388 4344
rect 126848 4304 207388 4332
rect 126848 4292 126854 4304
rect 207382 4292 207388 4304
rect 207440 4292 207446 4344
rect 209038 4292 209044 4344
rect 209096 4332 209102 4344
rect 268289 4335 268347 4341
rect 268289 4332 268301 4335
rect 209096 4304 268301 4332
rect 209096 4292 209102 4304
rect 268289 4301 268301 4304
rect 268335 4301 268347 4335
rect 268289 4295 268347 4301
rect 268565 4335 268623 4341
rect 268565 4301 268577 4335
rect 268611 4332 268623 4335
rect 505370 4332 505376 4344
rect 268611 4304 505376 4332
rect 268611 4301 268623 4304
rect 268565 4295 268623 4301
rect 505370 4292 505376 4304
rect 505428 4292 505434 4344
rect 129550 4224 129556 4276
rect 129608 4264 129614 4276
rect 214466 4264 214472 4276
rect 129608 4236 214472 4264
rect 129608 4224 129614 4236
rect 214466 4224 214472 4236
rect 214524 4224 214530 4276
rect 268197 4267 268255 4273
rect 268197 4233 268209 4267
rect 268243 4264 268255 4267
rect 268657 4267 268715 4273
rect 268243 4236 268608 4264
rect 268243 4233 268255 4236
rect 268197 4227 268255 4233
rect 103517 4199 103575 4205
rect 103517 4165 103529 4199
rect 103563 4196 103575 4199
rect 108393 4199 108451 4205
rect 108393 4196 108405 4199
rect 103563 4168 104664 4196
rect 103563 4165 103575 4168
rect 103517 4159 103575 4165
rect 63310 4088 63316 4140
rect 63368 4128 63374 4140
rect 74994 4128 75000 4140
rect 63368 4100 75000 4128
rect 63368 4088 63374 4100
rect 74994 4088 75000 4100
rect 75052 4088 75058 4140
rect 77202 4088 77208 4140
rect 77260 4128 77266 4140
rect 104526 4128 104532 4140
rect 77260 4100 104532 4128
rect 77260 4088 77266 4100
rect 104526 4088 104532 4100
rect 104584 4088 104590 4140
rect 104636 4128 104664 4168
rect 108132 4168 108405 4196
rect 108132 4128 108160 4168
rect 108393 4165 108405 4168
rect 108439 4165 108451 4199
rect 108393 4159 108451 4165
rect 110322 4156 110328 4208
rect 110380 4196 110386 4208
rect 113085 4199 113143 4205
rect 113085 4196 113097 4199
rect 110380 4168 113097 4196
rect 110380 4156 110386 4168
rect 113085 4165 113097 4168
rect 113131 4165 113143 4199
rect 113085 4159 113143 4165
rect 122650 4156 122656 4208
rect 122708 4196 122714 4208
rect 200298 4196 200304 4208
rect 122708 4168 200304 4196
rect 122708 4156 122714 4168
rect 200298 4156 200304 4168
rect 200356 4156 200362 4208
rect 200758 4156 200764 4208
rect 200816 4196 200822 4208
rect 268473 4199 268531 4205
rect 268473 4196 268485 4199
rect 200816 4168 268485 4196
rect 200816 4156 200822 4168
rect 268473 4165 268485 4168
rect 268519 4165 268531 4199
rect 268580 4196 268608 4236
rect 268657 4233 268669 4267
rect 268703 4264 268715 4267
rect 501782 4264 501788 4276
rect 268703 4236 501788 4264
rect 268703 4233 268715 4236
rect 268657 4227 268715 4233
rect 501782 4224 501788 4236
rect 501840 4224 501846 4276
rect 498194 4196 498200 4208
rect 268580 4168 498200 4196
rect 268473 4159 268531 4165
rect 498194 4156 498200 4168
rect 498252 4156 498258 4208
rect 111610 4128 111616 4140
rect 104636 4100 108160 4128
rect 108224 4100 111616 4128
rect 65978 4020 65984 4072
rect 66036 4060 66042 4072
rect 78582 4060 78588 4072
rect 66036 4032 78588 4060
rect 66036 4020 66042 4032
rect 78582 4020 78588 4032
rect 78640 4020 78646 4072
rect 79870 4020 79876 4072
rect 79928 4060 79934 4072
rect 108114 4060 108120 4072
rect 79928 4032 108120 4060
rect 79928 4020 79934 4032
rect 108114 4020 108120 4032
rect 108172 4020 108178 4072
rect 26329 3995 26387 4001
rect 26329 3961 26341 3995
rect 26375 3992 26387 3995
rect 29086 3992 29092 4004
rect 26375 3964 29092 3992
rect 26375 3961 26387 3964
rect 26329 3955 26387 3961
rect 29086 3952 29092 3964
rect 29144 3952 29150 4004
rect 60642 3952 60648 4004
rect 60700 3992 60706 4004
rect 66714 3992 66720 4004
rect 60700 3964 66720 3992
rect 60700 3952 60706 3964
rect 66714 3952 66720 3964
rect 66772 3952 66778 4004
rect 67542 3952 67548 4004
rect 67600 3992 67606 4004
rect 81161 3995 81219 4001
rect 81161 3992 81173 3995
rect 67600 3964 81173 3992
rect 67600 3952 67606 3964
rect 81161 3961 81173 3964
rect 81207 3961 81219 3995
rect 81161 3955 81219 3961
rect 81342 3952 81348 4004
rect 81400 3992 81406 4004
rect 108224 3992 108252 4100
rect 111610 4088 111616 4100
rect 111668 4088 111674 4140
rect 111705 4131 111763 4137
rect 111705 4097 111717 4131
rect 111751 4128 111763 4131
rect 117958 4128 117964 4140
rect 111751 4100 117964 4128
rect 111751 4097 111763 4100
rect 111705 4091 111763 4097
rect 117958 4088 117964 4100
rect 118016 4088 118022 4140
rect 184934 4128 184940 4140
rect 118068 4100 184940 4128
rect 108301 4063 108359 4069
rect 108301 4029 108313 4063
rect 108347 4060 108359 4063
rect 115198 4060 115204 4072
rect 108347 4032 115204 4060
rect 108347 4029 108359 4032
rect 108301 4023 108359 4029
rect 115198 4020 115204 4032
rect 115256 4020 115262 4072
rect 115842 4020 115848 4072
rect 115900 4060 115906 4072
rect 118068 4060 118096 4100
rect 184934 4088 184940 4100
rect 184992 4088 184998 4140
rect 185578 4088 185584 4140
rect 185636 4128 185642 4140
rect 196897 4131 196955 4137
rect 196897 4128 196909 4131
rect 185636 4100 196909 4128
rect 185636 4088 185642 4100
rect 196897 4097 196909 4100
rect 196943 4097 196955 4131
rect 196897 4091 196955 4097
rect 201402 4088 201408 4140
rect 201460 4128 201466 4140
rect 365806 4128 365812 4140
rect 201460 4100 365812 4128
rect 201460 4088 201466 4100
rect 365806 4088 365812 4100
rect 365864 4088 365870 4140
rect 366358 4088 366364 4140
rect 366416 4128 366422 4140
rect 368845 4131 368903 4137
rect 368845 4128 368857 4131
rect 366416 4100 368857 4128
rect 366416 4088 366422 4100
rect 368845 4097 368857 4100
rect 368891 4097 368903 4131
rect 368845 4091 368903 4097
rect 368937 4131 368995 4137
rect 368937 4097 368949 4131
rect 368983 4128 368995 4131
rect 373077 4131 373135 4137
rect 368983 4100 373028 4128
rect 368983 4097 368995 4100
rect 368937 4091 368995 4097
rect 115900 4032 118096 4060
rect 118145 4063 118203 4069
rect 115900 4020 115906 4032
rect 118145 4029 118157 4063
rect 118191 4060 118203 4063
rect 121181 4063 121239 4069
rect 121181 4060 121193 4063
rect 118191 4032 121193 4060
rect 118191 4029 118203 4032
rect 118145 4023 118203 4029
rect 121181 4029 121193 4032
rect 121227 4029 121239 4063
rect 121181 4023 121239 4029
rect 121362 4020 121368 4072
rect 121420 4060 121426 4072
rect 127713 4063 127771 4069
rect 121420 4032 127664 4060
rect 121420 4020 121426 4032
rect 81400 3964 108252 3992
rect 108393 3995 108451 4001
rect 81400 3952 81406 3964
rect 108393 3961 108405 3995
rect 108439 3992 108451 3995
rect 111705 3995 111763 4001
rect 111705 3992 111717 3995
rect 108439 3964 111717 3992
rect 108439 3961 108451 3964
rect 108393 3955 108451 3961
rect 111705 3961 111717 3964
rect 111751 3961 111763 3995
rect 111705 3955 111763 3961
rect 111797 3995 111855 4001
rect 111797 3961 111809 3995
rect 111843 3992 111855 3995
rect 114002 3992 114008 4004
rect 111843 3964 114008 3992
rect 111843 3961 111855 3964
rect 111797 3955 111855 3961
rect 114002 3952 114008 3964
rect 114060 3952 114066 4004
rect 117222 3952 117228 4004
rect 117280 3992 117286 4004
rect 117869 3995 117927 4001
rect 117869 3992 117881 3995
rect 117280 3964 117881 3992
rect 117280 3952 117286 3964
rect 117869 3961 117881 3964
rect 117915 3961 117927 3995
rect 117869 3955 117927 3961
rect 117958 3952 117964 4004
rect 118016 3992 118022 4004
rect 123478 3992 123484 4004
rect 118016 3964 123484 3992
rect 118016 3952 118022 3964
rect 123478 3952 123484 3964
rect 123536 3952 123542 4004
rect 124122 3952 124128 4004
rect 124180 3992 124186 4004
rect 127434 3992 127440 4004
rect 124180 3964 127440 3992
rect 124180 3952 124186 3964
rect 127434 3952 127440 3964
rect 127492 3952 127498 4004
rect 127636 3992 127664 4032
rect 127713 4029 127725 4063
rect 127759 4060 127771 4063
rect 188522 4060 188528 4072
rect 127759 4032 188528 4060
rect 127759 4029 127771 4032
rect 127713 4023 127771 4029
rect 188522 4020 188528 4032
rect 188580 4020 188586 4072
rect 204162 4020 204168 4072
rect 204220 4060 204226 4072
rect 372890 4060 372896 4072
rect 204220 4032 372896 4060
rect 204220 4020 204226 4032
rect 372890 4020 372896 4032
rect 372948 4020 372954 4072
rect 373000 4060 373028 4100
rect 373077 4097 373089 4131
rect 373123 4128 373135 4131
rect 383470 4128 383476 4140
rect 373123 4100 383476 4128
rect 373123 4097 373135 4100
rect 373077 4091 373135 4097
rect 383470 4088 383476 4100
rect 383528 4088 383534 4140
rect 383565 4131 383623 4137
rect 383565 4097 383577 4131
rect 383611 4128 383623 4131
rect 433242 4128 433248 4140
rect 383611 4100 433248 4128
rect 383611 4097 383623 4100
rect 383565 4091 383623 4097
rect 433242 4088 433248 4100
rect 433300 4088 433306 4140
rect 376478 4060 376484 4072
rect 373000 4032 376484 4060
rect 376478 4020 376484 4032
rect 376536 4020 376542 4072
rect 376570 4020 376576 4072
rect 376628 4060 376634 4072
rect 376628 4032 380112 4060
rect 376628 4020 376634 4032
rect 195606 3992 195612 4004
rect 127636 3964 195612 3992
rect 195606 3952 195612 3964
rect 195664 3952 195670 4004
rect 200117 3995 200175 4001
rect 200117 3961 200129 3995
rect 200163 3992 200175 3995
rect 206186 3992 206192 4004
rect 200163 3964 206192 3992
rect 200163 3961 200175 3964
rect 200117 3955 200175 3961
rect 206186 3952 206192 3964
rect 206244 3952 206250 4004
rect 206922 3952 206928 4004
rect 206980 3992 206986 4004
rect 379974 3992 379980 4004
rect 206980 3964 379980 3992
rect 206980 3952 206986 3964
rect 379974 3952 379980 3964
rect 380032 3952 380038 4004
rect 380084 3992 380112 4032
rect 380158 4020 380164 4072
rect 380216 4060 380222 4072
rect 383381 4063 383439 4069
rect 383381 4060 383393 4063
rect 380216 4032 383393 4060
rect 380216 4020 380222 4032
rect 383381 4029 383393 4032
rect 383427 4029 383439 4063
rect 383381 4023 383439 4029
rect 383657 4063 383715 4069
rect 383657 4029 383669 4063
rect 383703 4060 383715 4063
rect 447410 4060 447416 4072
rect 383703 4032 447416 4060
rect 383703 4029 383715 4032
rect 383657 4023 383715 4029
rect 447410 4020 447416 4032
rect 447468 4020 447474 4072
rect 382829 3995 382887 4001
rect 382829 3992 382841 3995
rect 380084 3964 382841 3992
rect 382829 3961 382841 3964
rect 382875 3961 382887 3995
rect 382829 3955 382887 3961
rect 382918 3952 382924 4004
rect 382976 3992 382982 4004
rect 475746 3992 475752 4004
rect 382976 3964 475752 3992
rect 382976 3952 382982 3964
rect 475746 3952 475752 3964
rect 475804 3952 475810 4004
rect 26237 3927 26295 3933
rect 26237 3893 26249 3927
rect 26283 3924 26295 3927
rect 30558 3924 30564 3936
rect 26283 3896 30564 3924
rect 26283 3893 26295 3896
rect 26237 3887 26295 3893
rect 30558 3884 30564 3896
rect 30616 3884 30622 3936
rect 64782 3884 64788 3936
rect 64840 3924 64846 3936
rect 77386 3924 77392 3936
rect 64840 3896 77392 3924
rect 64840 3884 64846 3896
rect 77386 3884 77392 3896
rect 77444 3884 77450 3936
rect 79778 3884 79784 3936
rect 79836 3924 79842 3936
rect 109310 3924 109316 3936
rect 79836 3896 109316 3924
rect 79836 3884 79842 3896
rect 109310 3884 109316 3896
rect 109368 3884 109374 3936
rect 109405 3927 109463 3933
rect 109405 3893 109417 3927
rect 109451 3924 109463 3927
rect 119890 3924 119896 3936
rect 109451 3896 119896 3924
rect 109451 3893 109463 3896
rect 109405 3887 109463 3893
rect 119890 3884 119896 3896
rect 119948 3884 119954 3936
rect 122742 3884 122748 3936
rect 122800 3924 122806 3936
rect 127529 3927 127587 3933
rect 127529 3924 127541 3927
rect 122800 3896 127541 3924
rect 122800 3884 122806 3896
rect 127529 3893 127541 3896
rect 127575 3893 127587 3927
rect 192018 3924 192024 3936
rect 127529 3887 127587 3893
rect 127636 3896 192024 3924
rect 17034 3816 17040 3868
rect 17092 3856 17098 3868
rect 17092 3828 26234 3856
rect 17092 3816 17098 3828
rect 19426 3748 19432 3800
rect 19484 3788 19490 3800
rect 20530 3788 20536 3800
rect 19484 3760 20536 3788
rect 19484 3748 19490 3760
rect 20530 3748 20536 3760
rect 20588 3748 20594 3800
rect 26206 3788 26234 3828
rect 66162 3816 66168 3868
rect 66220 3856 66226 3868
rect 79686 3856 79692 3868
rect 66220 3828 79692 3856
rect 66220 3816 66226 3828
rect 79686 3816 79692 3828
rect 79744 3816 79750 3868
rect 81250 3816 81256 3868
rect 81308 3856 81314 3868
rect 112806 3856 112812 3868
rect 81308 3828 112812 3856
rect 81308 3816 81314 3828
rect 112806 3816 112812 3828
rect 112864 3816 112870 3868
rect 112993 3859 113051 3865
rect 112993 3825 113005 3859
rect 113039 3856 113051 3859
rect 118053 3859 118111 3865
rect 118053 3856 118065 3859
rect 113039 3828 118065 3856
rect 113039 3825 113051 3828
rect 112993 3819 113051 3825
rect 118053 3825 118065 3828
rect 118099 3825 118111 3859
rect 118053 3819 118111 3825
rect 118602 3816 118608 3868
rect 118660 3856 118666 3868
rect 127636 3856 127664 3896
rect 192018 3884 192024 3896
rect 192076 3884 192082 3936
rect 194502 3884 194508 3936
rect 194560 3924 194566 3936
rect 204993 3927 205051 3933
rect 204993 3924 205005 3927
rect 194560 3896 205005 3924
rect 194560 3884 194566 3896
rect 204993 3893 205005 3896
rect 205039 3893 205051 3927
rect 204993 3887 205051 3893
rect 211062 3884 211068 3936
rect 211120 3924 211126 3936
rect 387150 3924 387156 3936
rect 211120 3896 387156 3924
rect 211120 3884 211126 3896
rect 387150 3884 387156 3896
rect 387208 3884 387214 3936
rect 199102 3856 199108 3868
rect 118660 3828 127664 3856
rect 127728 3828 199108 3856
rect 118660 3816 118666 3828
rect 36078 3788 36084 3800
rect 26206 3760 36084 3788
rect 36078 3748 36084 3760
rect 36136 3748 36142 3800
rect 70210 3748 70216 3800
rect 70268 3788 70274 3800
rect 71593 3791 71651 3797
rect 70268 3760 71544 3788
rect 70268 3748 70274 3760
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 33318 3720 33324 3732
rect 12308 3692 33324 3720
rect 12308 3680 12314 3692
rect 33318 3680 33324 3692
rect 33376 3680 33382 3732
rect 62022 3680 62028 3732
rect 62080 3720 62086 3732
rect 70302 3720 70308 3732
rect 62080 3692 70308 3720
rect 62080 3680 62086 3692
rect 70302 3680 70308 3692
rect 70360 3680 70366 3732
rect 71516 3720 71544 3760
rect 71593 3757 71605 3791
rect 71639 3788 71651 3791
rect 80882 3788 80888 3800
rect 71639 3760 80888 3788
rect 71639 3757 71651 3760
rect 71593 3751 71651 3757
rect 80882 3748 80888 3760
rect 80940 3748 80946 3800
rect 81161 3791 81219 3797
rect 81161 3757 81173 3791
rect 81207 3788 81219 3791
rect 82078 3788 82084 3800
rect 81207 3760 82084 3788
rect 81207 3757 81219 3760
rect 81161 3751 81219 3757
rect 82078 3748 82084 3760
rect 82136 3748 82142 3800
rect 82722 3748 82728 3800
rect 82780 3788 82786 3800
rect 108301 3791 108359 3797
rect 108301 3788 108313 3791
rect 82780 3760 108313 3788
rect 82780 3748 82786 3760
rect 108301 3757 108313 3760
rect 108347 3757 108359 3791
rect 108301 3751 108359 3757
rect 108390 3748 108396 3800
rect 108448 3788 108454 3800
rect 111797 3791 111855 3797
rect 111797 3788 111809 3791
rect 108448 3760 111809 3788
rect 108448 3748 108454 3760
rect 111797 3757 111809 3760
rect 111843 3757 111855 3791
rect 111797 3751 111855 3757
rect 114557 3791 114615 3797
rect 114557 3757 114569 3791
rect 114603 3788 114615 3791
rect 124674 3788 124680 3800
rect 114603 3760 124680 3788
rect 114603 3757 114615 3760
rect 114557 3751 114615 3757
rect 124674 3748 124680 3760
rect 124732 3748 124738 3800
rect 125502 3748 125508 3800
rect 125560 3788 125566 3800
rect 127437 3791 127495 3797
rect 127437 3788 127449 3791
rect 125560 3760 127449 3788
rect 125560 3748 125566 3760
rect 127437 3757 127449 3760
rect 127483 3757 127495 3791
rect 127437 3751 127495 3757
rect 127529 3791 127587 3797
rect 127529 3757 127541 3791
rect 127575 3788 127587 3791
rect 127728 3788 127756 3828
rect 199102 3816 199108 3828
rect 199160 3816 199166 3868
rect 202690 3856 202696 3868
rect 200086 3828 202696 3856
rect 127575 3760 127756 3788
rect 127575 3757 127587 3760
rect 127529 3751 127587 3757
rect 127802 3748 127808 3800
rect 127860 3788 127866 3800
rect 200086 3788 200114 3828
rect 202690 3816 202696 3828
rect 202748 3816 202754 3868
rect 213822 3816 213828 3868
rect 213880 3856 213886 3868
rect 394234 3856 394240 3868
rect 213880 3828 394240 3856
rect 213880 3816 213886 3828
rect 394234 3816 394240 3828
rect 394292 3816 394298 3868
rect 401318 3856 401324 3868
rect 398668 3828 401324 3856
rect 209774 3788 209780 3800
rect 127860 3760 200114 3788
rect 200408 3760 209780 3788
rect 127860 3748 127866 3760
rect 89162 3720 89168 3732
rect 71516 3692 89168 3720
rect 89162 3680 89168 3692
rect 89220 3680 89226 3732
rect 89257 3723 89315 3729
rect 89257 3689 89269 3723
rect 89303 3720 89315 3723
rect 89303 3692 92980 3720
rect 89303 3689 89315 3692
rect 89257 3683 89315 3689
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 26237 3655 26295 3661
rect 26237 3652 26249 3655
rect 7708 3624 26249 3652
rect 7708 3612 7714 3624
rect 26237 3621 26249 3624
rect 26283 3621 26295 3655
rect 27798 3652 27804 3664
rect 26237 3615 26295 3621
rect 26436 3624 27804 3652
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 26329 3587 26387 3593
rect 26329 3584 26341 3587
rect 2924 3556 26341 3584
rect 2924 3544 2930 3556
rect 26329 3553 26341 3556
rect 26375 3553 26387 3587
rect 26329 3547 26387 3553
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 26436 3516 26464 3624
rect 27798 3612 27804 3624
rect 27856 3612 27862 3664
rect 60458 3612 60464 3664
rect 60516 3652 60522 3664
rect 64417 3655 64475 3661
rect 64417 3652 64429 3655
rect 60516 3624 64429 3652
rect 60516 3612 60522 3624
rect 64417 3621 64429 3624
rect 64463 3621 64475 3655
rect 64417 3615 64475 3621
rect 68922 3612 68928 3664
rect 68980 3652 68986 3664
rect 84470 3652 84476 3664
rect 68980 3624 84476 3652
rect 68980 3612 68986 3624
rect 84470 3612 84476 3624
rect 84528 3612 84534 3664
rect 86862 3612 86868 3664
rect 86920 3652 86926 3664
rect 87509 3655 87567 3661
rect 87509 3652 87521 3655
rect 86920 3624 87521 3652
rect 86920 3612 86926 3624
rect 87509 3621 87521 3624
rect 87555 3621 87567 3655
rect 87509 3615 87567 3621
rect 87598 3612 87604 3664
rect 87656 3652 87662 3664
rect 92952 3652 92980 3692
rect 93118 3680 93124 3732
rect 93176 3720 93182 3732
rect 128170 3720 128176 3732
rect 93176 3692 128176 3720
rect 93176 3680 93182 3692
rect 128170 3680 128176 3692
rect 128228 3680 128234 3732
rect 132037 3723 132095 3729
rect 128280 3692 131988 3720
rect 122282 3652 122288 3664
rect 87656 3624 92888 3652
rect 92952 3624 122288 3652
rect 87656 3612 87662 3624
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28810 3584 28816 3596
rect 27764 3556 28816 3584
rect 27764 3544 27770 3556
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 37090 3584 37096 3596
rect 36044 3556 37096 3584
rect 36044 3544 36050 3556
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45370 3584 45376 3596
rect 44324 3556 45376 3584
rect 44324 3544 44330 3556
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 60550 3544 60556 3596
rect 60608 3584 60614 3596
rect 69106 3584 69112 3596
rect 60608 3556 69112 3584
rect 60608 3544 60614 3556
rect 69106 3544 69112 3556
rect 69164 3544 69170 3596
rect 71590 3544 71596 3596
rect 71648 3584 71654 3596
rect 92750 3584 92756 3596
rect 71648 3556 92756 3584
rect 71648 3544 71654 3556
rect 92750 3544 92756 3556
rect 92808 3544 92814 3596
rect 92860 3584 92888 3624
rect 122282 3612 122288 3624
rect 122340 3612 122346 3664
rect 126882 3612 126888 3664
rect 126940 3652 126946 3664
rect 128280 3652 128308 3692
rect 126940 3624 128308 3652
rect 126940 3612 126946 3624
rect 129642 3612 129648 3664
rect 129700 3652 129706 3664
rect 131960 3652 131988 3692
rect 132037 3689 132049 3723
rect 132083 3720 132095 3723
rect 200117 3723 200175 3729
rect 200117 3720 200129 3723
rect 132083 3692 200129 3720
rect 132083 3689 132095 3692
rect 132037 3683 132095 3689
rect 200117 3689 200129 3692
rect 200163 3689 200175 3723
rect 200117 3683 200175 3689
rect 200408 3652 200436 3760
rect 209774 3748 209780 3760
rect 209832 3748 209838 3800
rect 217962 3748 217968 3800
rect 218020 3788 218026 3800
rect 398668 3788 398696 3828
rect 401318 3816 401324 3828
rect 401376 3816 401382 3868
rect 218020 3760 398696 3788
rect 218020 3748 218026 3760
rect 398834 3748 398840 3800
rect 398892 3788 398898 3800
rect 400122 3788 400128 3800
rect 398892 3760 400128 3788
rect 398892 3748 398898 3760
rect 400122 3748 400128 3760
rect 400180 3748 400186 3800
rect 220722 3680 220728 3732
rect 220780 3720 220786 3732
rect 408402 3720 408408 3732
rect 220780 3692 408408 3720
rect 220780 3680 220786 3692
rect 408402 3680 408408 3692
rect 408460 3680 408466 3732
rect 129700 3624 131896 3652
rect 131960 3624 200436 3652
rect 200577 3655 200635 3661
rect 129700 3612 129706 3624
rect 93946 3584 93952 3596
rect 92860 3556 93952 3584
rect 93946 3544 93952 3556
rect 94004 3544 94010 3596
rect 94498 3544 94504 3596
rect 94556 3584 94562 3596
rect 131758 3584 131764 3596
rect 94556 3556 131764 3584
rect 94556 3544 94562 3556
rect 131758 3544 131764 3556
rect 131816 3544 131822 3596
rect 131868 3584 131896 3624
rect 200577 3621 200589 3655
rect 200623 3652 200635 3655
rect 212166 3652 212172 3664
rect 200623 3624 212172 3652
rect 200623 3621 200635 3624
rect 200577 3615 200635 3621
rect 212166 3612 212172 3624
rect 212224 3612 212230 3664
rect 224862 3612 224868 3664
rect 224920 3652 224926 3664
rect 415486 3652 415492 3664
rect 224920 3624 415492 3652
rect 224920 3612 224926 3624
rect 415486 3612 415492 3624
rect 415544 3612 415550 3664
rect 418798 3612 418804 3664
rect 418856 3652 418862 3664
rect 568022 3652 568028 3664
rect 418856 3624 568028 3652
rect 418856 3612 418862 3624
rect 568022 3612 568028 3624
rect 568080 3612 568086 3664
rect 213362 3584 213368 3596
rect 131868 3556 213368 3584
rect 213362 3544 213368 3556
rect 213420 3544 213426 3596
rect 227622 3544 227628 3596
rect 227680 3584 227686 3596
rect 422570 3584 422576 3596
rect 227680 3556 422576 3584
rect 227680 3544 227686 3556
rect 422570 3544 422576 3556
rect 422628 3544 422634 3596
rect 429654 3584 429660 3596
rect 423600 3556 429660 3584
rect 1728 3488 26464 3516
rect 1728 3476 1734 3488
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53742 3516 53748 3528
rect 52512 3488 53748 3516
rect 52512 3476 52518 3488
rect 53742 3476 53748 3488
rect 53800 3476 53806 3528
rect 54018 3476 54024 3528
rect 54076 3516 54082 3528
rect 54938 3516 54944 3528
rect 54076 3488 54944 3516
rect 54076 3476 54082 3488
rect 54938 3476 54944 3488
rect 54996 3476 55002 3528
rect 56410 3476 56416 3528
rect 56468 3516 56474 3528
rect 58434 3516 58440 3528
rect 56468 3488 58440 3516
rect 56468 3476 56474 3488
rect 58434 3476 58440 3488
rect 58492 3476 58498 3528
rect 59170 3476 59176 3528
rect 59228 3516 59234 3528
rect 64322 3516 64328 3528
rect 59228 3488 64328 3516
rect 59228 3476 59234 3488
rect 64322 3476 64328 3488
rect 64380 3476 64386 3528
rect 64417 3519 64475 3525
rect 64417 3485 64429 3519
rect 64463 3516 64475 3519
rect 67910 3516 67916 3528
rect 64463 3488 67916 3516
rect 64463 3485 64475 3488
rect 64417 3479 64475 3485
rect 67910 3476 67916 3488
rect 67968 3476 67974 3528
rect 70394 3476 70400 3528
rect 70452 3516 70458 3528
rect 71777 3519 71835 3525
rect 71777 3516 71789 3519
rect 70452 3488 71789 3516
rect 70452 3476 70458 3488
rect 71777 3485 71789 3488
rect 71823 3485 71835 3519
rect 71777 3479 71835 3485
rect 71869 3519 71927 3525
rect 71869 3485 71881 3519
rect 71915 3516 71927 3519
rect 85666 3516 85672 3528
rect 71915 3488 85672 3516
rect 71915 3485 71927 3488
rect 71869 3479 71927 3485
rect 85666 3476 85672 3488
rect 85724 3476 85730 3528
rect 86770 3476 86776 3528
rect 86828 3516 86834 3528
rect 88889 3519 88947 3525
rect 88889 3516 88901 3519
rect 86828 3488 88901 3516
rect 86828 3476 86834 3488
rect 88889 3485 88901 3488
rect 88935 3485 88947 3519
rect 88889 3479 88947 3485
rect 88978 3476 88984 3528
rect 89036 3516 89042 3528
rect 90358 3516 90364 3528
rect 89036 3488 90364 3516
rect 89036 3476 89042 3488
rect 90358 3476 90364 3488
rect 90416 3476 90422 3528
rect 90453 3519 90511 3525
rect 90453 3485 90465 3519
rect 90499 3516 90511 3519
rect 114557 3519 114615 3525
rect 114557 3516 114569 3519
rect 90499 3488 114569 3516
rect 90499 3485 90511 3488
rect 90453 3479 90511 3485
rect 114557 3485 114569 3488
rect 114603 3485 114615 3519
rect 114557 3479 114615 3485
rect 119338 3476 119344 3528
rect 119396 3516 119402 3528
rect 121086 3516 121092 3528
rect 119396 3488 121092 3516
rect 119396 3476 119402 3488
rect 121086 3476 121092 3488
rect 121144 3476 121150 3528
rect 121181 3519 121239 3525
rect 121181 3485 121193 3519
rect 121227 3516 121239 3519
rect 127713 3519 127771 3525
rect 127713 3516 127725 3519
rect 121227 3488 127725 3516
rect 121227 3485 121239 3488
rect 121181 3479 121239 3485
rect 127713 3485 127725 3488
rect 127759 3485 127771 3519
rect 127713 3479 127771 3485
rect 127805 3519 127863 3525
rect 127805 3485 127817 3519
rect 127851 3516 127863 3519
rect 132037 3519 132095 3525
rect 132037 3516 132049 3519
rect 127851 3488 132049 3516
rect 127851 3485 127863 3488
rect 127805 3479 127863 3485
rect 132037 3485 132049 3488
rect 132083 3485 132095 3519
rect 132037 3479 132095 3485
rect 132402 3476 132408 3528
rect 132460 3516 132466 3528
rect 220446 3516 220452 3528
rect 132460 3488 220452 3516
rect 132460 3476 132466 3488
rect 220446 3476 220452 3488
rect 220504 3476 220510 3528
rect 230382 3476 230388 3528
rect 230440 3516 230446 3528
rect 423600 3516 423628 3556
rect 429654 3544 429660 3556
rect 429712 3544 429718 3596
rect 489914 3544 489920 3596
rect 489972 3584 489978 3596
rect 491110 3584 491116 3596
rect 489972 3556 491116 3584
rect 489972 3544 489978 3556
rect 491110 3544 491116 3556
rect 491168 3544 491174 3596
rect 230440 3488 423628 3516
rect 230440 3476 230446 3488
rect 423674 3476 423680 3528
rect 423732 3516 423738 3528
rect 424962 3516 424968 3528
rect 423732 3488 424968 3516
rect 423732 3476 423738 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 448514 3476 448520 3528
rect 448572 3516 448578 3528
rect 449802 3516 449808 3528
rect 448572 3488 449808 3516
rect 448572 3476 448578 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 456794 3476 456800 3528
rect 456852 3516 456858 3528
rect 458082 3516 458088 3528
rect 456852 3488 458088 3516
rect 456852 3476 456858 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 27614 3448 27620 3460
rect 624 3420 27620 3448
rect 624 3408 630 3420
rect 27614 3408 27620 3420
rect 27672 3408 27678 3460
rect 57790 3408 57796 3460
rect 57848 3448 57854 3460
rect 60826 3448 60832 3460
rect 57848 3420 60832 3448
rect 57848 3408 57854 3420
rect 60826 3408 60832 3420
rect 60884 3408 60890 3460
rect 61930 3408 61936 3460
rect 61988 3448 61994 3460
rect 71498 3448 71504 3460
rect 61988 3420 71504 3448
rect 61988 3408 61994 3420
rect 71498 3408 71504 3420
rect 71556 3408 71562 3460
rect 71682 3408 71688 3460
rect 71740 3448 71746 3460
rect 91554 3448 91560 3460
rect 71740 3420 91560 3448
rect 71740 3408 71746 3420
rect 91554 3408 91560 3420
rect 91612 3408 91618 3460
rect 92382 3408 92388 3460
rect 92440 3448 92446 3460
rect 135254 3448 135260 3460
rect 92440 3420 135260 3448
rect 92440 3408 92446 3420
rect 135254 3408 135260 3420
rect 135312 3408 135318 3460
rect 137922 3408 137928 3460
rect 137980 3448 137986 3460
rect 231026 3448 231032 3460
rect 137980 3420 231032 3448
rect 137980 3408 137986 3420
rect 231026 3408 231032 3420
rect 231084 3408 231090 3460
rect 237282 3408 237288 3460
rect 237340 3448 237346 3460
rect 443822 3448 443828 3460
rect 237340 3420 443828 3448
rect 237340 3408 237346 3420
rect 443822 3408 443828 3420
rect 443880 3408 443886 3460
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 9582 3380 9588 3392
rect 8812 3352 9588 3380
rect 8812 3340 8818 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 10962 3380 10968 3392
rect 10008 3352 10968 3380
rect 10008 3340 10014 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 12342 3380 12348 3392
rect 11204 3352 12348 3380
rect 11204 3340 11210 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 16482 3380 16488 3392
rect 15988 3352 16488 3380
rect 15988 3340 15994 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 19242 3380 19248 3392
rect 18288 3352 19248 3380
rect 18288 3340 18294 3352
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 24762 3380 24768 3392
rect 24268 3352 24768 3380
rect 24268 3340 24274 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25314 3340 25320 3392
rect 25372 3380 25378 3392
rect 26142 3380 26148 3392
rect 25372 3352 26148 3380
rect 25372 3340 25378 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 57882 3340 57888 3392
rect 57940 3380 57946 3392
rect 63218 3380 63224 3392
rect 57940 3352 63224 3380
rect 57940 3340 57946 3352
rect 63218 3340 63224 3352
rect 63276 3340 63282 3392
rect 64690 3340 64696 3392
rect 64748 3380 64754 3392
rect 76190 3380 76196 3392
rect 64748 3352 76196 3380
rect 64748 3340 64754 3352
rect 76190 3340 76196 3352
rect 76248 3340 76254 3392
rect 78490 3340 78496 3392
rect 78548 3380 78554 3392
rect 78548 3352 104112 3380
rect 78548 3340 78554 3352
rect 55122 3272 55128 3324
rect 55180 3312 55186 3324
rect 56042 3312 56048 3324
rect 55180 3284 56048 3312
rect 55180 3272 55186 3284
rect 56042 3272 56048 3284
rect 56100 3272 56106 3324
rect 66070 3272 66076 3324
rect 66128 3312 66134 3324
rect 71593 3315 71651 3321
rect 71593 3312 71605 3315
rect 66128 3284 71605 3312
rect 66128 3272 66134 3284
rect 71593 3281 71605 3284
rect 71639 3281 71651 3315
rect 71593 3275 71651 3281
rect 71777 3315 71835 3321
rect 71777 3281 71789 3315
rect 71823 3312 71835 3315
rect 87966 3312 87972 3324
rect 71823 3284 87972 3312
rect 71823 3281 71835 3284
rect 71777 3275 71835 3281
rect 87966 3272 87972 3284
rect 88024 3272 88030 3324
rect 88061 3315 88119 3321
rect 88061 3281 88073 3315
rect 88107 3312 88119 3315
rect 90361 3315 90419 3321
rect 90361 3312 90373 3315
rect 88107 3284 90373 3312
rect 88107 3281 88119 3284
rect 88061 3275 88119 3281
rect 90361 3281 90373 3284
rect 90407 3281 90419 3315
rect 90361 3275 90419 3281
rect 90450 3272 90456 3324
rect 90508 3312 90514 3324
rect 90508 3284 103514 3312
rect 90508 3272 90514 3284
rect 57698 3204 57704 3256
rect 57756 3244 57762 3256
rect 62022 3244 62028 3256
rect 57756 3216 62028 3244
rect 57756 3204 57762 3216
rect 62022 3204 62028 3216
rect 62080 3204 62086 3256
rect 63402 3204 63408 3256
rect 63460 3244 63466 3256
rect 73798 3244 73804 3256
rect 63460 3216 73804 3244
rect 63460 3204 63466 3216
rect 73798 3204 73804 3216
rect 73856 3204 73862 3256
rect 77110 3204 77116 3256
rect 77168 3244 77174 3256
rect 102226 3244 102232 3256
rect 77168 3216 102232 3244
rect 77168 3204 77174 3216
rect 102226 3204 102232 3216
rect 102284 3204 102290 3256
rect 103486 3244 103514 3284
rect 103977 3247 104035 3253
rect 103977 3244 103989 3247
rect 103486 3216 103989 3244
rect 103977 3213 103989 3216
rect 104023 3213 104035 3247
rect 104084 3244 104112 3352
rect 104158 3340 104164 3392
rect 104216 3380 104222 3392
rect 106918 3380 106924 3392
rect 104216 3352 106924 3380
rect 104216 3340 104222 3352
rect 106918 3340 106924 3352
rect 106976 3340 106982 3392
rect 109405 3383 109463 3389
rect 109405 3380 109417 3383
rect 107028 3352 109417 3380
rect 104253 3315 104311 3321
rect 104253 3281 104265 3315
rect 104299 3312 104311 3315
rect 106829 3315 106887 3321
rect 106829 3312 106841 3315
rect 104299 3284 106841 3312
rect 104299 3281 104311 3284
rect 104253 3275 104311 3281
rect 106829 3281 106841 3284
rect 106875 3281 106887 3315
rect 106829 3275 106887 3281
rect 105722 3244 105728 3256
rect 104084 3216 105728 3244
rect 103977 3207 104035 3213
rect 105722 3204 105728 3216
rect 105780 3204 105786 3256
rect 105814 3204 105820 3256
rect 105872 3244 105878 3256
rect 107028 3244 107056 3352
rect 109405 3349 109417 3352
rect 109451 3349 109463 3383
rect 109405 3343 109463 3349
rect 111702 3340 111708 3392
rect 111760 3380 111766 3392
rect 177850 3380 177856 3392
rect 111760 3352 177856 3380
rect 111760 3340 111766 3352
rect 177850 3340 177856 3352
rect 177908 3340 177914 3392
rect 200577 3383 200635 3389
rect 200577 3380 200589 3383
rect 177960 3352 200589 3380
rect 107105 3315 107163 3321
rect 107105 3281 107117 3315
rect 107151 3312 107163 3315
rect 116394 3312 116400 3324
rect 107151 3284 116400 3312
rect 107151 3281 107163 3284
rect 107105 3275 107163 3281
rect 116394 3272 116400 3284
rect 116452 3272 116458 3324
rect 174262 3312 174268 3324
rect 117976 3284 174268 3312
rect 105872 3216 107056 3244
rect 105872 3204 105878 3216
rect 107562 3204 107568 3256
rect 107620 3244 107626 3256
rect 112993 3247 113051 3253
rect 112993 3244 113005 3247
rect 107620 3216 113005 3244
rect 107620 3204 107626 3216
rect 112993 3213 113005 3216
rect 113039 3213 113051 3247
rect 112993 3207 113051 3213
rect 113085 3247 113143 3253
rect 113085 3213 113097 3247
rect 113131 3244 113143 3247
rect 117976 3244 118004 3284
rect 174262 3272 174268 3284
rect 174320 3272 174326 3324
rect 177390 3272 177396 3324
rect 177448 3312 177454 3324
rect 177960 3312 177988 3352
rect 200577 3349 200589 3352
rect 200623 3349 200635 3383
rect 355873 3383 355931 3389
rect 355873 3380 355885 3383
rect 200577 3343 200635 3349
rect 204916 3352 355885 3380
rect 177448 3284 177988 3312
rect 178037 3315 178095 3321
rect 177448 3272 177454 3284
rect 178037 3281 178049 3315
rect 178083 3312 178095 3315
rect 193214 3312 193220 3324
rect 178083 3284 193220 3312
rect 178083 3281 178095 3284
rect 178037 3275 178095 3281
rect 193214 3272 193220 3284
rect 193272 3272 193278 3324
rect 194229 3315 194287 3321
rect 194229 3281 194241 3315
rect 194275 3312 194287 3315
rect 194275 3284 195376 3312
rect 194275 3281 194287 3284
rect 194229 3275 194287 3281
rect 113131 3216 118004 3244
rect 118053 3247 118111 3253
rect 113131 3213 113143 3216
rect 113085 3207 113143 3213
rect 118053 3213 118065 3247
rect 118099 3244 118111 3247
rect 167178 3244 167184 3256
rect 118099 3216 167184 3244
rect 118099 3213 118111 3216
rect 118053 3207 118111 3213
rect 167178 3204 167184 3216
rect 167236 3204 167242 3256
rect 175918 3204 175924 3256
rect 175976 3244 175982 3256
rect 195149 3247 195207 3253
rect 195149 3244 195161 3247
rect 175976 3216 195161 3244
rect 175976 3204 175982 3216
rect 195149 3213 195161 3216
rect 195195 3213 195207 3247
rect 195149 3207 195207 3213
rect 55030 3136 55036 3188
rect 55088 3176 55094 3188
rect 57238 3176 57244 3188
rect 55088 3148 57244 3176
rect 55088 3136 55094 3148
rect 57238 3136 57244 3148
rect 57296 3136 57302 3188
rect 63310 3136 63316 3188
rect 63368 3176 63374 3188
rect 72602 3176 72608 3188
rect 63368 3148 72608 3176
rect 63368 3136 63374 3148
rect 72602 3136 72608 3148
rect 72660 3136 72666 3188
rect 75822 3136 75828 3188
rect 75880 3176 75886 3188
rect 101030 3176 101036 3188
rect 75880 3148 101036 3176
rect 75880 3136 75886 3148
rect 101030 3136 101036 3148
rect 101088 3136 101094 3188
rect 101398 3136 101404 3188
rect 101456 3176 101462 3188
rect 103517 3179 103575 3185
rect 103517 3176 103529 3179
rect 101456 3148 103529 3176
rect 101456 3136 101462 3148
rect 103517 3145 103529 3148
rect 103563 3145 103575 3179
rect 103517 3139 103575 3145
rect 103606 3136 103612 3188
rect 103664 3176 103670 3188
rect 160094 3176 160100 3188
rect 103664 3148 160100 3176
rect 103664 3136 103670 3148
rect 160094 3136 160100 3148
rect 160152 3136 160158 3188
rect 160738 3136 160744 3188
rect 160796 3176 160802 3188
rect 160796 3148 161474 3176
rect 160796 3136 160802 3148
rect 56502 3068 56508 3120
rect 56560 3108 56566 3120
rect 59630 3108 59636 3120
rect 56560 3080 59636 3108
rect 56560 3068 56566 3080
rect 59630 3068 59636 3080
rect 59688 3068 59694 3120
rect 68830 3068 68836 3120
rect 68888 3108 68894 3120
rect 71869 3111 71927 3117
rect 71869 3108 71881 3111
rect 68888 3080 71881 3108
rect 68888 3068 68894 3080
rect 71869 3077 71881 3080
rect 71915 3077 71927 3111
rect 71869 3071 71927 3077
rect 75730 3068 75736 3120
rect 75788 3108 75794 3120
rect 99834 3108 99840 3120
rect 75788 3080 99840 3108
rect 75788 3068 75794 3080
rect 99834 3068 99840 3080
rect 99892 3068 99898 3120
rect 103241 3111 103299 3117
rect 103241 3108 103253 3111
rect 99944 3080 103253 3108
rect 74442 3000 74448 3052
rect 74500 3040 74506 3052
rect 98638 3040 98644 3052
rect 74500 3012 98644 3040
rect 74500 3000 74506 3012
rect 98638 3000 98644 3012
rect 98696 3000 98702 3052
rect 99944 3040 99972 3080
rect 103241 3077 103253 3080
rect 103287 3077 103299 3111
rect 153010 3108 153016 3120
rect 103241 3071 103299 3077
rect 103486 3080 153016 3108
rect 98748 3012 99972 3040
rect 74258 2932 74264 2984
rect 74316 2972 74322 2984
rect 97442 2972 97448 2984
rect 74316 2944 97448 2972
rect 74316 2932 74322 2944
rect 97442 2932 97448 2944
rect 97500 2932 97506 2984
rect 98748 2972 98776 3012
rect 100662 3000 100668 3052
rect 100720 3040 100726 3052
rect 103486 3040 103514 3080
rect 153010 3068 153016 3080
rect 153068 3068 153074 3120
rect 155218 3068 155224 3120
rect 155276 3108 155282 3120
rect 161290 3108 161296 3120
rect 155276 3080 161296 3108
rect 155276 3068 155282 3080
rect 161290 3068 161296 3080
rect 161348 3068 161354 3120
rect 161446 3108 161474 3148
rect 170398 3136 170404 3188
rect 170456 3176 170462 3188
rect 189718 3176 189724 3188
rect 170456 3148 189724 3176
rect 170456 3136 170462 3148
rect 189718 3136 189724 3148
rect 189776 3136 189782 3188
rect 190362 3136 190368 3188
rect 190420 3176 190426 3188
rect 195241 3179 195299 3185
rect 195241 3176 195253 3179
rect 190420 3148 195253 3176
rect 190420 3136 190426 3148
rect 195241 3145 195253 3148
rect 195287 3145 195299 3179
rect 195348 3176 195376 3284
rect 197262 3272 197268 3324
rect 197320 3312 197326 3324
rect 204916 3312 204944 3352
rect 355873 3349 355885 3352
rect 355919 3349 355931 3383
rect 355873 3343 355931 3349
rect 355962 3340 355968 3392
rect 356020 3380 356026 3392
rect 356020 3352 356192 3380
rect 356020 3340 356026 3352
rect 197320 3284 204944 3312
rect 204993 3315 205051 3321
rect 197320 3272 197326 3284
rect 204993 3281 205005 3315
rect 205039 3312 205051 3315
rect 349065 3315 349123 3321
rect 349065 3312 349077 3315
rect 205039 3284 349077 3312
rect 205039 3281 205051 3284
rect 204993 3275 205051 3281
rect 349065 3281 349077 3284
rect 349111 3281 349123 3315
rect 349065 3275 349123 3281
rect 349154 3272 349160 3324
rect 349212 3312 349218 3324
rect 350442 3312 350448 3324
rect 349212 3284 350448 3312
rect 349212 3272 349218 3284
rect 350442 3272 350448 3284
rect 350500 3272 350506 3324
rect 351178 3272 351184 3324
rect 351236 3312 351242 3324
rect 351236 3284 351776 3312
rect 351236 3272 351242 3284
rect 195425 3247 195483 3253
rect 195425 3213 195437 3247
rect 195471 3244 195483 3247
rect 344554 3244 344560 3256
rect 195471 3216 344560 3244
rect 195471 3213 195483 3216
rect 195425 3207 195483 3213
rect 344554 3204 344560 3216
rect 344612 3204 344618 3256
rect 344649 3247 344707 3253
rect 344649 3213 344661 3247
rect 344695 3244 344707 3247
rect 349801 3247 349859 3253
rect 349801 3244 349813 3247
rect 344695 3216 349813 3244
rect 344695 3213 344707 3216
rect 344649 3207 344707 3213
rect 349801 3213 349813 3216
rect 349847 3213 349859 3247
rect 349801 3207 349859 3213
rect 349893 3247 349951 3253
rect 349893 3213 349905 3247
rect 349939 3244 349951 3247
rect 351638 3244 351644 3256
rect 349939 3216 351644 3244
rect 349939 3213 349951 3216
rect 349893 3207 349951 3213
rect 351638 3204 351644 3216
rect 351696 3204 351702 3256
rect 351748 3244 351776 3284
rect 351822 3272 351828 3324
rect 351880 3312 351886 3324
rect 356164 3312 356192 3352
rect 358078 3340 358084 3392
rect 358136 3380 358142 3392
rect 369213 3383 369271 3389
rect 369213 3380 369225 3383
rect 358136 3352 369225 3380
rect 358136 3340 358142 3352
rect 369213 3349 369225 3352
rect 369259 3349 369271 3383
rect 369213 3343 369271 3349
rect 369486 3340 369492 3392
rect 369544 3380 369550 3392
rect 373077 3383 373135 3389
rect 373077 3380 373089 3383
rect 369544 3352 373089 3380
rect 369544 3340 369550 3352
rect 373077 3349 373089 3352
rect 373123 3349 373135 3383
rect 373077 3343 373135 3349
rect 373258 3340 373264 3392
rect 373316 3380 373322 3392
rect 426158 3380 426164 3392
rect 373316 3352 426164 3380
rect 373316 3340 373322 3352
rect 426158 3340 426164 3352
rect 426216 3340 426222 3392
rect 383470 3312 383476 3324
rect 351880 3284 356100 3312
rect 356164 3284 383476 3312
rect 351880 3272 351886 3284
rect 355870 3244 355876 3256
rect 351748 3216 355876 3244
rect 355870 3204 355876 3216
rect 355928 3204 355934 3256
rect 356072 3244 356100 3284
rect 383470 3272 383476 3284
rect 383528 3272 383534 3324
rect 383562 3272 383568 3324
rect 383620 3312 383626 3324
rect 418982 3312 418988 3324
rect 383620 3284 418988 3312
rect 383620 3272 383626 3284
rect 418982 3272 418988 3284
rect 419040 3272 419046 3324
rect 368937 3247 368995 3253
rect 368937 3244 368949 3247
rect 356072 3216 368949 3244
rect 368937 3213 368949 3216
rect 368983 3213 368995 3247
rect 369394 3244 369400 3256
rect 368937 3207 368995 3213
rect 369044 3216 369400 3244
rect 337470 3176 337476 3188
rect 195348 3148 337476 3176
rect 195241 3139 195299 3145
rect 337470 3136 337476 3148
rect 337528 3136 337534 3188
rect 337562 3136 337568 3188
rect 337620 3176 337626 3188
rect 344189 3179 344247 3185
rect 344189 3176 344201 3179
rect 337620 3148 344201 3176
rect 337620 3136 337626 3148
rect 344189 3145 344201 3148
rect 344235 3145 344247 3179
rect 344189 3139 344247 3145
rect 344278 3136 344284 3188
rect 344336 3176 344342 3188
rect 369044 3176 369072 3216
rect 369394 3204 369400 3216
rect 369452 3204 369458 3256
rect 369489 3247 369547 3253
rect 369489 3213 369501 3247
rect 369535 3244 369547 3247
rect 411898 3244 411904 3256
rect 369535 3216 411904 3244
rect 369535 3213 369547 3216
rect 369489 3207 369547 3213
rect 411898 3204 411904 3216
rect 411956 3204 411962 3256
rect 344336 3148 369072 3176
rect 369121 3179 369179 3185
rect 344336 3136 344342 3148
rect 369121 3145 369133 3179
rect 369167 3176 369179 3179
rect 404814 3176 404820 3188
rect 369167 3148 404820 3176
rect 369167 3145 369179 3148
rect 369121 3139 369179 3145
rect 404814 3136 404820 3148
rect 404872 3136 404878 3188
rect 175458 3108 175464 3120
rect 161446 3080 175464 3108
rect 175458 3068 175464 3080
rect 175516 3068 175522 3120
rect 177298 3068 177304 3120
rect 177356 3108 177362 3120
rect 178129 3111 178187 3117
rect 178129 3108 178141 3111
rect 177356 3080 178141 3108
rect 177356 3068 177362 3080
rect 178129 3077 178141 3080
rect 178175 3077 178187 3111
rect 178129 3071 178187 3077
rect 181530 3068 181536 3120
rect 181588 3108 181594 3120
rect 237006 3108 237012 3120
rect 181588 3080 237012 3108
rect 181588 3068 181594 3080
rect 237006 3068 237012 3080
rect 237064 3068 237070 3120
rect 307754 3068 307760 3120
rect 307812 3108 307818 3120
rect 309042 3108 309048 3120
rect 307812 3080 309048 3108
rect 307812 3068 307818 3080
rect 309042 3068 309048 3080
rect 309100 3068 309106 3120
rect 309778 3068 309784 3120
rect 309836 3108 309842 3120
rect 320637 3111 320695 3117
rect 320637 3108 320649 3111
rect 309836 3080 320649 3108
rect 309836 3068 309842 3080
rect 320637 3077 320649 3080
rect 320683 3077 320695 3111
rect 320637 3071 320695 3077
rect 320729 3111 320787 3117
rect 320729 3077 320741 3111
rect 320775 3108 320787 3111
rect 461578 3108 461584 3120
rect 320775 3080 461584 3108
rect 320775 3077 320787 3080
rect 320729 3071 320787 3077
rect 461578 3068 461584 3080
rect 461636 3068 461642 3120
rect 583386 3108 583392 3120
rect 583347 3080 583392 3108
rect 583386 3068 583392 3080
rect 583444 3068 583450 3120
rect 149514 3040 149520 3052
rect 100720 3012 103514 3040
rect 104912 3012 149520 3040
rect 100720 3000 100726 3012
rect 97644 2944 98776 2972
rect 59262 2864 59268 2916
rect 59320 2904 59326 2916
rect 65518 2904 65524 2916
rect 59320 2876 65524 2904
rect 59320 2864 59326 2876
rect 65518 2864 65524 2876
rect 65576 2864 65582 2916
rect 73062 2864 73068 2916
rect 73120 2904 73126 2916
rect 95142 2904 95148 2916
rect 73120 2876 95148 2904
rect 73120 2864 73126 2876
rect 95142 2864 95148 2876
rect 95200 2864 95206 2916
rect 95878 2864 95884 2916
rect 95936 2904 95942 2916
rect 97537 2907 97595 2913
rect 97537 2904 97549 2907
rect 95936 2876 97549 2904
rect 95936 2864 95942 2876
rect 97537 2873 97549 2876
rect 97583 2873 97595 2907
rect 97537 2867 97595 2873
rect 74350 2796 74356 2848
rect 74408 2836 74414 2848
rect 96246 2836 96252 2848
rect 74408 2808 96252 2836
rect 74408 2796 74414 2808
rect 96246 2796 96252 2808
rect 96304 2796 96310 2848
rect 97644 2836 97672 2944
rect 99282 2932 99288 2984
rect 99340 2972 99346 2984
rect 104912 2972 104940 3012
rect 149514 3000 149520 3012
rect 149572 3000 149578 3052
rect 156598 3000 156604 3052
rect 156656 3040 156662 3052
rect 164878 3040 164884 3052
rect 156656 3012 164884 3040
rect 156656 3000 156662 3012
rect 164878 3000 164884 3012
rect 164936 3000 164942 3052
rect 167638 3000 167644 3052
rect 167696 3040 167702 3052
rect 182542 3040 182548 3052
rect 167696 3012 182548 3040
rect 167696 3000 167702 3012
rect 182542 3000 182548 3012
rect 182600 3000 182606 3052
rect 184842 3000 184848 3052
rect 184900 3040 184906 3052
rect 184900 3012 186360 3040
rect 184900 3000 184906 3012
rect 99340 2944 104940 2972
rect 104989 2975 105047 2981
rect 99340 2932 99346 2944
rect 104989 2941 105001 2975
rect 105035 2972 105047 2975
rect 145926 2972 145932 2984
rect 105035 2944 145932 2972
rect 105035 2941 105047 2944
rect 104989 2935 105047 2941
rect 145926 2932 145932 2944
rect 145984 2932 145990 2984
rect 166258 2932 166264 2984
rect 166316 2972 166322 2984
rect 179046 2972 179052 2984
rect 166316 2944 179052 2972
rect 166316 2932 166322 2944
rect 179046 2932 179052 2944
rect 179104 2932 179110 2984
rect 180058 2932 180064 2984
rect 180116 2972 180122 2984
rect 186225 2975 186283 2981
rect 186225 2972 186237 2975
rect 180116 2944 186237 2972
rect 180116 2932 180122 2944
rect 186225 2941 186237 2944
rect 186271 2941 186283 2975
rect 186225 2935 186283 2941
rect 97721 2907 97779 2913
rect 97721 2873 97733 2907
rect 97767 2904 97779 2907
rect 103333 2907 103391 2913
rect 103333 2904 103345 2907
rect 97767 2876 103345 2904
rect 97767 2873 97779 2876
rect 97721 2867 97779 2873
rect 103333 2873 103345 2876
rect 103379 2873 103391 2907
rect 103333 2867 103391 2873
rect 103517 2907 103575 2913
rect 103517 2873 103529 2907
rect 103563 2904 103575 2907
rect 142430 2904 142436 2916
rect 103563 2876 142436 2904
rect 103563 2873 103575 2876
rect 103517 2867 103575 2873
rect 142430 2864 142436 2876
rect 142488 2864 142494 2916
rect 142798 2864 142804 2916
rect 142856 2904 142862 2916
rect 156598 2904 156604 2916
rect 142856 2876 156604 2904
rect 142856 2864 142862 2876
rect 156598 2864 156604 2876
rect 156656 2864 156662 2916
rect 157978 2864 157984 2916
rect 158036 2904 158042 2916
rect 168374 2904 168380 2916
rect 158036 2876 168380 2904
rect 158036 2864 158042 2876
rect 168374 2864 168380 2876
rect 168432 2864 168438 2916
rect 169018 2864 169024 2916
rect 169076 2904 169082 2916
rect 186130 2904 186136 2916
rect 169076 2876 186136 2904
rect 169076 2864 169082 2876
rect 186130 2864 186136 2876
rect 186188 2864 186194 2916
rect 186332 2904 186360 3012
rect 187602 3000 187608 3052
rect 187660 3040 187666 3052
rect 194229 3043 194287 3049
rect 194229 3040 194241 3043
rect 187660 3012 194241 3040
rect 187660 3000 187666 3012
rect 194229 3009 194241 3012
rect 194275 3009 194287 3043
rect 194229 3003 194287 3009
rect 194321 3043 194379 3049
rect 194321 3009 194333 3043
rect 194367 3040 194379 3043
rect 330386 3040 330392 3052
rect 194367 3012 330392 3040
rect 194367 3009 194379 3012
rect 194321 3003 194379 3009
rect 330386 3000 330392 3012
rect 330444 3000 330450 3052
rect 330478 3000 330484 3052
rect 330536 3040 330542 3052
rect 333149 3043 333207 3049
rect 333149 3040 333161 3043
rect 330536 3012 333161 3040
rect 330536 3000 330542 3012
rect 333149 3009 333161 3012
rect 333195 3009 333207 3043
rect 333149 3003 333207 3009
rect 333238 3000 333244 3052
rect 333296 3040 333302 3052
rect 348050 3040 348056 3052
rect 333296 3012 348056 3040
rect 333296 3000 333302 3012
rect 348050 3000 348056 3012
rect 348108 3000 348114 3052
rect 349065 3043 349123 3049
rect 349065 3009 349077 3043
rect 349111 3040 349123 3043
rect 349709 3043 349767 3049
rect 349709 3040 349721 3043
rect 349111 3012 349721 3040
rect 349111 3009 349123 3012
rect 349065 3003 349123 3009
rect 349709 3009 349721 3012
rect 349755 3009 349767 3043
rect 349709 3003 349767 3009
rect 349801 3043 349859 3049
rect 349801 3009 349813 3043
rect 349847 3040 349859 3043
rect 362310 3040 362316 3052
rect 349847 3012 362316 3040
rect 349847 3009 349859 3012
rect 349801 3003 349859 3009
rect 362310 3000 362316 3012
rect 362368 3000 362374 3052
rect 362402 3000 362408 3052
rect 362460 3040 362466 3052
rect 369121 3043 369179 3049
rect 369121 3040 369133 3043
rect 362460 3012 369133 3040
rect 362460 3000 362466 3012
rect 369121 3009 369133 3012
rect 369167 3009 369179 3043
rect 369121 3003 369179 3009
rect 369213 3043 369271 3049
rect 369213 3009 369225 3043
rect 369259 3040 369271 3043
rect 397730 3040 397736 3052
rect 369259 3012 397736 3040
rect 369259 3009 369271 3012
rect 369213 3003 369271 3009
rect 397730 3000 397736 3012
rect 397788 3000 397794 3052
rect 186501 2975 186559 2981
rect 186501 2941 186513 2975
rect 186547 2972 186559 2975
rect 233418 2972 233424 2984
rect 186547 2944 233424 2972
rect 186547 2941 186559 2944
rect 186501 2935 186559 2941
rect 233418 2932 233424 2944
rect 233476 2932 233482 2984
rect 315390 2932 315396 2984
rect 315448 2972 315454 2984
rect 320729 2975 320787 2981
rect 320729 2972 320741 2975
rect 315448 2944 320741 2972
rect 315448 2932 315454 2944
rect 320729 2941 320741 2944
rect 320775 2941 320787 2975
rect 320729 2935 320787 2941
rect 320821 2975 320879 2981
rect 320821 2941 320833 2975
rect 320867 2972 320879 2975
rect 454494 2972 454500 2984
rect 320867 2944 454500 2972
rect 320867 2941 320879 2944
rect 320821 2935 320879 2941
rect 454494 2932 454500 2944
rect 454552 2932 454558 2984
rect 194321 2907 194379 2913
rect 194321 2904 194333 2907
rect 186332 2876 194333 2904
rect 194321 2873 194333 2876
rect 194367 2873 194379 2907
rect 194321 2867 194379 2873
rect 195149 2907 195207 2913
rect 195149 2873 195161 2907
rect 195195 2904 195207 2907
rect 196802 2904 196808 2916
rect 195195 2876 196808 2904
rect 195195 2873 195207 2876
rect 195149 2867 195207 2873
rect 196802 2864 196808 2876
rect 196860 2864 196866 2916
rect 196897 2907 196955 2913
rect 196897 2873 196909 2907
rect 196943 2904 196955 2907
rect 323302 2904 323308 2916
rect 196943 2876 323308 2904
rect 196943 2873 196955 2876
rect 196897 2867 196955 2873
rect 323302 2864 323308 2876
rect 323360 2864 323366 2916
rect 323670 2864 323676 2916
rect 323728 2904 323734 2916
rect 333882 2904 333888 2916
rect 323728 2876 333888 2904
rect 323728 2864 323734 2876
rect 333882 2864 333888 2876
rect 333940 2864 333946 2916
rect 340966 2904 340972 2916
rect 334084 2876 340972 2904
rect 96356 2808 97672 2836
rect 95234 2728 95240 2780
rect 95292 2768 95298 2780
rect 96356 2768 96384 2808
rect 97902 2796 97908 2848
rect 97960 2836 97966 2848
rect 103425 2839 103483 2845
rect 97960 2808 103376 2836
rect 97960 2796 97966 2808
rect 95292 2740 96384 2768
rect 103348 2768 103376 2808
rect 103425 2805 103437 2839
rect 103471 2836 103483 2839
rect 138842 2836 138848 2848
rect 103471 2808 138848 2836
rect 103471 2805 103483 2808
rect 103425 2799 103483 2805
rect 138842 2796 138848 2808
rect 138900 2796 138906 2848
rect 159358 2796 159364 2848
rect 159416 2836 159422 2848
rect 171962 2836 171968 2848
rect 159416 2808 171968 2836
rect 159416 2796 159422 2808
rect 171962 2796 171968 2808
rect 172020 2796 172026 2848
rect 173250 2796 173256 2848
rect 173308 2836 173314 2848
rect 178037 2839 178095 2845
rect 178037 2836 178049 2839
rect 173308 2808 178049 2836
rect 173308 2796 173314 2808
rect 178037 2805 178049 2808
rect 178083 2805 178095 2839
rect 178037 2799 178095 2805
rect 178129 2839 178187 2845
rect 178129 2805 178141 2839
rect 178175 2836 178187 2839
rect 229830 2836 229836 2848
rect 178175 2808 229836 2836
rect 178175 2805 178187 2808
rect 178129 2799 178187 2805
rect 229830 2796 229836 2808
rect 229888 2796 229894 2848
rect 312538 2796 312544 2848
rect 312596 2836 312602 2848
rect 320821 2839 320879 2845
rect 320821 2836 320833 2839
rect 312596 2808 320833 2836
rect 312596 2796 312602 2808
rect 320821 2805 320833 2808
rect 320867 2805 320879 2839
rect 333977 2839 334035 2845
rect 333977 2836 333989 2839
rect 320821 2799 320879 2805
rect 320928 2808 333989 2836
rect 104989 2771 105047 2777
rect 104989 2768 105001 2771
rect 103348 2740 105001 2768
rect 95292 2728 95298 2740
rect 104989 2737 105001 2740
rect 105035 2737 105047 2771
rect 104989 2731 105047 2737
rect 320637 2771 320695 2777
rect 320637 2737 320649 2771
rect 320683 2768 320695 2771
rect 320928 2768 320956 2808
rect 333977 2805 333989 2808
rect 334023 2805 334035 2839
rect 333977 2799 334035 2805
rect 320683 2740 320956 2768
rect 320683 2737 320695 2740
rect 320637 2731 320695 2737
rect 324314 2728 324320 2780
rect 324372 2768 324378 2780
rect 325602 2768 325608 2780
rect 324372 2740 325608 2768
rect 324372 2728 324378 2740
rect 325602 2728 325608 2740
rect 325660 2728 325666 2780
rect 333149 2771 333207 2777
rect 333149 2737 333161 2771
rect 333195 2768 333207 2771
rect 334084 2768 334112 2876
rect 340966 2864 340972 2876
rect 341024 2864 341030 2916
rect 341518 2864 341524 2916
rect 341576 2904 341582 2916
rect 344649 2907 344707 2913
rect 344649 2904 344661 2907
rect 341576 2876 344661 2904
rect 341576 2864 341582 2876
rect 344649 2873 344661 2876
rect 344695 2873 344707 2907
rect 344649 2867 344707 2873
rect 344741 2907 344799 2913
rect 344741 2873 344753 2907
rect 344787 2904 344799 2907
rect 355226 2904 355232 2916
rect 344787 2876 355232 2904
rect 344787 2873 344799 2876
rect 344741 2867 344799 2873
rect 355226 2864 355232 2876
rect 355284 2864 355290 2916
rect 355318 2864 355324 2916
rect 355376 2904 355382 2916
rect 355873 2907 355931 2913
rect 355376 2876 355824 2904
rect 355376 2864 355382 2876
rect 334161 2839 334219 2845
rect 334161 2805 334173 2839
rect 334207 2836 334219 2839
rect 355689 2839 355747 2845
rect 355689 2836 355701 2839
rect 334207 2808 355701 2836
rect 334207 2805 334219 2808
rect 334161 2799 334219 2805
rect 355689 2805 355701 2808
rect 355735 2805 355747 2839
rect 355689 2799 355747 2805
rect 333195 2740 334112 2768
rect 355796 2768 355824 2876
rect 355873 2873 355885 2907
rect 355919 2904 355931 2907
rect 358722 2904 358728 2916
rect 355919 2876 358728 2904
rect 355919 2873 355931 2876
rect 355873 2867 355931 2873
rect 358722 2864 358728 2876
rect 358780 2864 358786 2916
rect 390646 2904 390652 2916
rect 358924 2876 390652 2904
rect 355965 2839 356023 2845
rect 355965 2805 355977 2839
rect 356011 2836 356023 2839
rect 358817 2839 358875 2845
rect 358817 2836 358829 2839
rect 356011 2808 358829 2836
rect 356011 2805 356023 2808
rect 355965 2799 356023 2805
rect 358817 2805 358829 2808
rect 358863 2805 358875 2839
rect 358817 2799 358875 2805
rect 358924 2768 358952 2876
rect 390646 2864 390652 2876
rect 390704 2864 390710 2916
rect 359001 2839 359059 2845
rect 359001 2805 359013 2839
rect 359047 2836 359059 2839
rect 440326 2836 440332 2848
rect 359047 2808 440332 2836
rect 359047 2805 359059 2808
rect 359001 2799 359059 2805
rect 440326 2796 440332 2808
rect 440384 2796 440390 2848
rect 355796 2740 358952 2768
rect 333195 2737 333207 2740
rect 333149 2731 333207 2737
rect 103241 2703 103299 2709
rect 103241 2669 103253 2703
rect 103287 2700 103299 2703
rect 103517 2703 103575 2709
rect 103517 2700 103529 2703
rect 103287 2672 103529 2700
rect 103287 2669 103299 2672
rect 103241 2663 103299 2669
rect 103517 2669 103529 2672
rect 103563 2669 103575 2703
rect 103517 2663 103575 2669
<< via1 >>
rect 166908 700952 166960 701004
rect 300124 700952 300176 701004
rect 24308 700884 24360 700936
rect 185124 700884 185176 700936
rect 162768 700816 162820 700868
rect 332508 700816 332560 700868
rect 164148 700748 164200 700800
rect 348792 700748 348844 700800
rect 40500 700680 40552 700732
rect 236000 700680 236052 700732
rect 154488 700612 154540 700664
rect 397460 700612 397512 700664
rect 157248 700544 157300 700596
rect 413652 700544 413704 700596
rect 147588 700476 147640 700528
rect 462320 700476 462372 700528
rect 105452 700408 105504 700460
rect 147312 700408 147364 700460
rect 150348 700408 150400 700460
rect 478512 700408 478564 700460
rect 72976 700340 73028 700392
rect 147128 700340 147180 700392
rect 147220 700340 147272 700392
rect 494796 700340 494848 700392
rect 89168 700272 89220 700324
rect 146944 700272 146996 700324
rect 147036 700272 147088 700324
rect 527180 700272 527232 700324
rect 172428 700204 172480 700256
rect 283840 700204 283892 700256
rect 169668 700136 169720 700188
rect 267648 700136 267700 700188
rect 173808 700068 173860 700120
rect 235172 700068 235224 700120
rect 137836 700000 137888 700052
rect 182180 700000 182232 700052
rect 179328 699932 179380 699984
rect 218980 699932 219032 699984
rect 154120 699864 154172 699916
rect 180064 699864 180116 699916
rect 176568 699796 176620 699848
rect 202788 699796 202840 699848
rect 170312 699728 170364 699780
rect 180800 699728 180852 699780
rect 251456 699660 251508 699712
rect 252468 699660 252520 699712
rect 381176 699660 381228 699712
rect 382188 699660 382240 699712
rect 443736 688644 443788 688696
rect 463332 688644 463384 688696
rect 3424 683136 3476 683188
rect 230480 683136 230532 683188
rect 3516 670692 3568 670744
rect 193128 670692 193180 670744
rect 252468 666476 252520 666528
rect 300768 666476 300820 666528
rect 542360 666408 542412 666460
rect 542360 661716 542412 661768
rect 196992 650360 197044 650412
rect 236000 650564 236052 650616
rect 4804 650020 4856 650072
rect 40132 650020 40184 650072
rect 230480 646119 230532 646128
rect 230480 646085 230489 646119
rect 230489 646085 230523 646119
rect 230523 646085 230532 646119
rect 230480 646076 230532 646085
rect 230480 645507 230532 645516
rect 230480 645473 230489 645507
rect 230489 645473 230523 645507
rect 230523 645473 230532 645507
rect 230480 645464 230532 645473
rect 202696 645396 202748 645448
rect 443828 644784 443880 644836
rect 443736 644580 443788 644632
rect 3792 644444 3844 644496
rect 104716 644444 104768 644496
rect 98644 644240 98696 644292
rect 104256 644240 104308 644292
rect 204536 644240 204588 644292
rect 236184 644240 236236 644292
rect 240692 644240 240744 644292
rect 429200 644308 429252 644360
rect 193128 643671 193180 643680
rect 193128 643637 193137 643671
rect 193137 643637 193171 643671
rect 193171 643637 193180 643671
rect 193128 643628 193180 643637
rect 199384 643628 199436 643680
rect 199568 643628 199620 643680
rect 185124 643560 185176 643612
rect 196624 643560 196676 643612
rect 198004 643560 198056 643612
rect 204536 643560 204588 643612
rect 185124 643288 185176 643340
rect 3608 643220 3660 643272
rect 133788 643220 133840 643272
rect 193128 643263 193180 643272
rect 193128 643229 193137 643263
rect 193137 643229 193171 643263
rect 193171 643229 193180 643263
rect 193128 643220 193180 643229
rect 208400 643152 208452 643204
rect 220176 643152 220228 643204
rect 192208 643084 192260 643136
rect 206560 643084 206612 643136
rect 209688 643084 209740 643136
rect 220084 643084 220136 643136
rect 160008 642880 160060 642932
rect 190920 642880 190972 642932
rect 196992 642812 197044 642864
rect 201776 642404 201828 642456
rect 201776 642200 201828 642252
rect 192208 642132 192260 642184
rect 236184 642268 236236 642320
rect 241612 642268 241664 642320
rect 364340 642268 364392 642320
rect 471796 640840 471848 640892
rect 580540 641656 580592 641708
rect 459560 640296 459612 640348
rect 196900 640203 196952 640212
rect 196900 640169 196909 640203
rect 196909 640169 196943 640203
rect 196943 640169 196952 640203
rect 196900 640160 196952 640169
rect 185124 639956 185176 640008
rect 193128 639999 193180 640008
rect 193128 639965 193137 639999
rect 193137 639965 193171 639999
rect 193171 639965 193180 639999
rect 193128 639956 193180 639965
rect 185124 639684 185176 639736
rect 443736 639616 443788 639668
rect 193128 639591 193180 639600
rect 193128 639557 193137 639591
rect 193137 639557 193171 639591
rect 193171 639557 193180 639591
rect 193128 639548 193180 639557
rect 224868 639548 224920 639600
rect 230480 639548 230532 639600
rect 202236 639208 202288 639260
rect 443644 639183 443696 639192
rect 443644 639149 443653 639183
rect 443653 639149 443687 639183
rect 443687 639149 443696 639183
rect 443644 639140 443696 639149
rect 443736 639140 443788 639192
rect 193128 636191 193180 636200
rect 193128 636157 193137 636191
rect 193137 636157 193171 636191
rect 193171 636157 193180 636191
rect 193128 636148 193180 636157
rect 185124 636080 185176 636132
rect 185124 635808 185176 635860
rect 193128 635783 193180 635792
rect 193128 635749 193137 635783
rect 193137 635749 193171 635783
rect 193171 635749 193180 635783
rect 193128 635740 193180 635749
rect 220084 634652 220136 634704
rect 220268 634695 220320 634704
rect 220268 634661 220277 634695
rect 220277 634661 220311 634695
rect 220311 634661 220320 634695
rect 220268 634652 220320 634661
rect 193128 632519 193180 632528
rect 193128 632485 193137 632519
rect 193137 632485 193171 632519
rect 193171 632485 193180 632519
rect 193128 632476 193180 632485
rect 185124 632408 185176 632460
rect 185124 632136 185176 632188
rect 193128 632111 193180 632120
rect 193128 632077 193137 632111
rect 193137 632077 193171 632111
rect 193171 632077 193180 632111
rect 193128 632068 193180 632077
rect 219900 631975 219952 631984
rect 219900 631941 219909 631975
rect 219909 631941 219943 631975
rect 219943 631941 219952 631975
rect 219900 631932 219952 631941
rect 220360 631932 220412 631984
rect 193128 628983 193180 628992
rect 193128 628949 193137 628983
rect 193137 628949 193171 628983
rect 193171 628949 193180 628983
rect 193128 628940 193180 628949
rect 185124 628872 185176 628924
rect 196900 628668 196952 628720
rect 185124 628600 185176 628652
rect 193128 628507 193180 628516
rect 193128 628473 193137 628507
rect 193137 628473 193171 628507
rect 193171 628473 193180 628507
rect 193128 628464 193180 628473
rect 196992 628328 197044 628380
rect 542360 617856 542412 617908
rect 382188 615476 382240 615528
rect 542360 613368 542412 613420
rect 114468 606364 114520 606416
rect 118976 606364 119028 606416
rect 119988 606364 120040 606416
rect 211160 606364 211212 606416
rect 3148 593308 3200 593360
rect 40040 593308 40092 593360
rect 167460 591268 167512 591320
rect 580172 591268 580224 591320
rect 167460 579640 167512 579692
rect 210424 579640 210476 579692
rect 167460 577464 167512 577516
rect 580172 577464 580224 577516
rect 424968 570596 425020 570648
rect 443736 570596 443788 570648
rect 410340 569916 410392 569968
rect 424324 569916 424376 569968
rect 424968 569916 425020 569968
rect 404268 566856 404320 566908
rect 427820 566448 427872 566500
rect 92388 558900 92440 558952
rect 391848 558900 391900 558952
rect 3332 553392 3384 553444
rect 218060 553392 218112 553444
rect 99288 542376 99340 542428
rect 391388 542376 391440 542428
rect 391756 542376 391808 542428
rect 3332 540880 3384 540932
rect 40224 540880 40276 540932
rect 111708 536800 111760 536852
rect 580172 536800 580224 536852
rect 417700 534012 417752 534064
rect 580724 534012 580776 534064
rect 401600 533944 401652 533996
rect 402060 533944 402112 533996
rect 542360 533944 542412 533996
rect 143448 533400 143500 533452
rect 401600 533400 401652 533452
rect 115848 533332 115900 533384
rect 417700 533332 417752 533384
rect 3332 527144 3384 527196
rect 223580 527144 223632 527196
rect 114468 524424 114520 524476
rect 580172 524424 580224 524476
rect 108948 510620 109000 510672
rect 580172 510620 580224 510672
rect 3332 500964 3384 501016
rect 226340 500964 226392 501016
rect 3148 489812 3200 489864
rect 40132 489812 40184 489864
rect 104808 484372 104860 484424
rect 579620 484372 579672 484424
rect 3056 474716 3108 474768
rect 230480 474716 230532 474768
rect 106188 470568 106240 470620
rect 579988 470568 580040 470620
rect 3332 462340 3384 462392
rect 200764 462340 200816 462392
rect 424324 458124 424376 458176
rect 424968 458124 425020 458176
rect 580172 458124 580224 458176
rect 100760 457444 100812 457496
rect 424968 457444 425020 457496
rect 3332 448536 3384 448588
rect 233240 448536 233292 448588
rect 3332 437384 3384 437436
rect 40040 437384 40092 437436
rect 96528 430584 96580 430636
rect 580172 430584 580224 430636
rect 3148 422288 3200 422340
rect 237380 422288 237432 422340
rect 391756 419432 391808 419484
rect 579620 419432 579672 419484
rect 3332 409844 3384 409896
rect 217324 409844 217376 409896
rect 95148 404336 95200 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 240140 397468 240192 397520
rect 89628 378156 89680 378208
rect 579620 378156 579672 378208
rect 3332 371220 3384 371272
rect 245660 371220 245712 371272
rect 391848 365644 391900 365696
rect 580172 365644 580224 365696
rect 88248 351908 88300 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 247040 345040 247092 345092
rect 82544 324300 82596 324352
rect 579988 324300 580040 324352
rect 3608 318792 3660 318844
rect 252744 318792 252796 318844
rect 147128 314576 147180 314628
rect 190460 314576 190512 314628
rect 8208 314508 8260 314560
rect 197452 314508 197504 314560
rect 3424 314440 3476 314492
rect 204628 314440 204680 314492
rect 3516 314372 3568 314424
rect 209780 314372 209832 314424
rect 135076 314304 135128 314356
rect 443644 314304 443696 314356
rect 137836 314236 137888 314288
rect 558920 314236 558972 314288
rect 133052 314168 133104 314220
rect 580264 314168 580316 314220
rect 130660 314100 130712 314152
rect 580356 314100 580408 314152
rect 128268 314032 128320 314084
rect 580540 314032 580592 314084
rect 125508 313964 125560 314016
rect 580448 313964 580500 314016
rect 123392 313896 123444 313948
rect 580632 313896 580684 313948
rect 147312 313828 147364 313880
rect 187792 313828 187844 313880
rect 220084 313352 220136 313404
rect 228732 313352 228784 313404
rect 144736 313284 144788 313336
rect 147220 313284 147272 313336
rect 195704 313284 195756 313336
rect 196992 313284 197044 313336
rect 220176 313284 220228 313336
rect 221556 313284 221608 313336
rect 185124 313216 185176 313268
rect 185676 313216 185728 313268
rect 146944 313148 146996 313200
rect 140320 313080 140372 313132
rect 147036 313080 147088 313132
rect 87328 313012 87380 313064
rect 88248 313012 88300 313064
rect 94504 313012 94556 313064
rect 95148 313012 95200 313064
rect 104164 313012 104216 313064
rect 104808 313012 104860 313064
rect 113824 313012 113876 313064
rect 114468 313012 114520 313064
rect 142712 313012 142764 313064
rect 143448 313012 143500 313064
rect 149888 313012 149940 313064
rect 150348 313012 150400 313064
rect 152280 313080 152332 313132
rect 153108 313080 153160 313132
rect 159548 313080 159600 313132
rect 160008 313080 160060 313132
rect 161940 313080 161992 313132
rect 162768 313080 162820 313132
rect 169208 313080 169260 313132
rect 169668 313080 169720 313132
rect 171600 313080 171652 313132
rect 172428 313080 172480 313132
rect 178776 313080 178828 313132
rect 179328 313080 179380 313132
rect 180064 313080 180116 313132
rect 185400 313080 185452 313132
rect 192576 313148 192628 313200
rect 193128 313148 193180 313200
rect 185676 313080 185728 313132
rect 200120 313080 200172 313132
rect 201776 313148 201828 313200
rect 214288 313148 214340 313200
rect 207020 313080 207072 313132
rect 210424 313080 210476 313132
rect 216680 313080 216732 313132
rect 217324 313080 217376 313132
rect 243176 313080 243228 313132
rect 200764 313012 200816 313064
rect 236000 313012 236052 313064
rect 77668 312944 77720 312996
rect 304632 312944 304684 312996
rect 3884 312876 3936 312928
rect 250444 312876 250496 312928
rect 6368 312808 6420 312860
rect 257620 312808 257672 312860
rect 5448 312740 5500 312792
rect 260012 312740 260064 312792
rect 5356 312672 5408 312724
rect 267280 312672 267332 312724
rect 3332 312604 3384 312656
rect 264980 312604 265032 312656
rect 3976 312536 4028 312588
rect 272064 312536 272116 312588
rect 5264 312468 5316 312520
rect 274640 312468 274692 312520
rect 3700 312400 3752 312452
rect 276940 312400 276992 312452
rect 3792 312332 3844 312384
rect 279332 312332 279384 312384
rect 5172 312264 5224 312316
rect 281724 312264 281776 312316
rect 5080 312196 5132 312248
rect 284300 312196 284352 312248
rect 6276 312128 6328 312180
rect 286508 312128 286560 312180
rect 4988 312060 5040 312112
rect 288900 312060 288952 312112
rect 6184 311992 6236 312044
rect 291384 311992 291436 312044
rect 3608 311924 3660 311976
rect 293960 311924 294012 311976
rect 84936 311856 84988 311908
rect 580172 311856 580224 311908
rect 79968 310428 80020 310480
rect 75276 310360 75328 310412
rect 70308 310335 70360 310344
rect 70308 310301 70317 310335
rect 70317 310301 70351 310335
rect 70351 310301 70360 310335
rect 70308 310292 70360 310301
rect 72884 310292 72936 310344
rect 304540 310428 304592 310480
rect 303528 310360 303580 310412
rect 304356 310292 304408 310344
rect 60648 310267 60700 310276
rect 60648 310233 60657 310267
rect 60657 310233 60691 310267
rect 60691 310233 60700 310267
rect 60648 310224 60700 310233
rect 63224 310267 63276 310276
rect 63224 310233 63233 310267
rect 63233 310233 63267 310267
rect 63267 310233 63276 310267
rect 63224 310224 63276 310233
rect 65616 310224 65668 310276
rect 303436 310224 303488 310276
rect 55956 310199 56008 310208
rect 55956 310165 55965 310199
rect 55965 310165 55999 310199
rect 55999 310165 56008 310199
rect 55956 310156 56008 310165
rect 58440 310156 58492 310208
rect 303252 310156 303304 310208
rect 36728 310131 36780 310140
rect 36728 310097 36737 310131
rect 36737 310097 36771 310131
rect 36771 310097 36780 310131
rect 36728 310088 36780 310097
rect 39120 310131 39172 310140
rect 39120 310097 39129 310131
rect 39129 310097 39163 310131
rect 39163 310097 39172 310131
rect 39120 310088 39172 310097
rect 41328 310131 41380 310140
rect 41328 310097 41337 310131
rect 41337 310097 41371 310131
rect 41371 310097 41380 310131
rect 41328 310088 41380 310097
rect 46388 310131 46440 310140
rect 46388 310097 46397 310131
rect 46397 310097 46431 310131
rect 46431 310097 46440 310131
rect 46388 310088 46440 310097
rect 48780 310131 48832 310140
rect 48780 310097 48789 310131
rect 48789 310097 48823 310131
rect 48823 310097 48832 310131
rect 48780 310088 48832 310097
rect 53564 310088 53616 310140
rect 4712 310020 4764 310072
rect 255320 310020 255372 310072
rect 4068 309952 4120 310004
rect 262496 309952 262548 310004
rect 269672 309995 269724 310004
rect 269672 309961 269681 309995
rect 269681 309961 269715 309995
rect 269715 309961 269724 309995
rect 269672 309952 269724 309961
rect 296168 309995 296220 310004
rect 296168 309961 296177 309995
rect 296177 309961 296211 309995
rect 296211 309961 296220 309995
rect 296168 309952 296220 309961
rect 304264 310088 304316 310140
rect 3884 309816 3936 309868
rect 303068 310020 303120 310072
rect 298560 309952 298612 310004
rect 304724 309952 304776 310004
rect 4896 309680 4948 309732
rect 3424 309612 3476 309664
rect 580816 309544 580868 309596
rect 580632 309476 580684 309528
rect 580724 309408 580776 309460
rect 580540 309340 580592 309392
rect 580356 309272 580408 309324
rect 580448 309204 580500 309256
rect 580264 309136 580316 309188
rect 2964 306212 3016 306264
rect 6368 306212 6420 306264
rect 304724 299412 304776 299464
rect 580172 299412 580224 299464
rect 2780 293224 2832 293276
rect 4712 293224 4764 293276
rect 303528 273164 303580 273216
rect 579988 273164 580040 273216
rect 2780 267180 2832 267232
rect 5448 267180 5500 267232
rect 304632 259360 304684 259412
rect 579804 259360 579856 259412
rect 304540 245556 304592 245608
rect 580172 245556 580224 245608
rect 304448 233180 304500 233232
rect 579988 233180 580040 233232
rect 2780 214956 2832 215008
rect 5356 214956 5408 215008
rect 303436 206932 303488 206984
rect 579620 206932 579672 206984
rect 303252 166948 303304 167000
rect 580172 166948 580224 167000
rect 2780 163344 2832 163396
rect 5264 163344 5316 163396
rect 304356 153144 304408 153196
rect 580172 153144 580224 153196
rect 303344 126896 303396 126948
rect 579620 126896 579672 126948
rect 2780 123836 2832 123888
rect 4804 123836 4856 123888
rect 2780 110712 2832 110764
rect 5172 110712 5224 110764
rect 2780 97724 2832 97776
rect 6276 97724 6328 97776
rect 303160 86912 303212 86964
rect 580172 86912 580224 86964
rect 2780 85144 2832 85196
rect 5080 85144 5132 85196
rect 304264 73108 304316 73160
rect 579988 73108 580040 73160
rect 2780 71612 2832 71664
rect 4988 71612 5040 71664
rect 303068 46860 303120 46912
rect 580172 46860 580224 46912
rect 3148 45500 3200 45552
rect 6184 45500 6236 45552
rect 107338 33804 107390 33856
rect 302976 33056 303028 33108
rect 580172 33056 580224 33108
rect 2780 32852 2832 32904
rect 4896 32852 4948 32904
rect 250812 31764 250864 31816
rect 251088 31764 251140 31816
rect 261944 31764 261996 31816
rect 262128 31764 262180 31816
rect 264704 31764 264756 31816
rect 264888 31764 264940 31816
rect 19248 31696 19300 31748
rect 36268 31696 36320 31748
rect 41328 31696 41380 31748
rect 46940 31696 46992 31748
rect 110972 31696 111024 31748
rect 160744 31696 160796 31748
rect 188988 31696 189040 31748
rect 330484 31696 330536 31748
rect 16488 31628 16540 31680
rect 35164 31628 35216 31680
rect 44088 31628 44140 31680
rect 47952 31628 48004 31680
rect 68836 31628 68888 31680
rect 20536 31560 20588 31612
rect 37372 31560 37424 31612
rect 42708 31560 42760 31612
rect 47400 31560 47452 31612
rect 83188 31628 83240 31680
rect 90272 31628 90324 31680
rect 90364 31628 90416 31680
rect 94504 31628 94556 31680
rect 106004 31628 106056 31680
rect 156604 31628 156656 31680
rect 200764 31628 200816 31680
rect 215668 31628 215720 31680
rect 358084 31628 358136 31680
rect 85764 31560 85816 31612
rect 93676 31560 93728 31612
rect 95884 31560 95936 31612
rect 104348 31560 104400 31612
rect 155224 31560 155276 31612
rect 165528 31560 165580 31612
rect 15108 31492 15160 31544
rect 34612 31492 34664 31544
rect 38568 31492 38620 31544
rect 45744 31492 45796 31544
rect 72608 31492 72660 31544
rect 87512 31492 87564 31544
rect 157984 31492 158036 31544
rect 162216 31492 162268 31544
rect 204904 31560 204956 31612
rect 209044 31560 209096 31612
rect 351184 31560 351236 31612
rect 205548 31492 205600 31544
rect 348424 31492 348476 31544
rect 13728 31424 13780 31476
rect 34060 31424 34112 31476
rect 86500 31424 86552 31476
rect 101404 31424 101456 31476
rect 10968 31356 11020 31408
rect 32404 31356 32456 31408
rect 70952 31356 71004 31408
rect 88984 31356 89036 31408
rect 12348 31288 12400 31340
rect 33140 31288 33192 31340
rect 34428 31288 34480 31340
rect 43536 31288 43588 31340
rect 45468 31288 45520 31340
rect 48504 31288 48556 31340
rect 84844 31288 84896 31340
rect 105544 31356 105596 31408
rect 109316 31356 109368 31408
rect 159364 31424 159416 31476
rect 166908 31424 166960 31476
rect 209044 31424 209096 31476
rect 237932 31424 237984 31476
rect 238668 31424 238720 31476
rect 376024 31424 376076 31476
rect 170404 31356 170456 31408
rect 219072 31356 219124 31408
rect 362224 31356 362276 31408
rect 115848 31288 115900 31340
rect 169024 31288 169076 31340
rect 198648 31288 198700 31340
rect 341524 31288 341576 31340
rect 9588 31220 9640 31272
rect 31852 31220 31904 31272
rect 35808 31220 35860 31272
rect 44180 31220 44232 31272
rect 77024 31220 77076 31272
rect 102324 31220 102376 31272
rect 225696 31220 225748 31272
rect 369124 31220 369176 31272
rect 6828 31152 6880 31204
rect 30748 31152 30800 31204
rect 33048 31152 33100 31204
rect 42984 31152 43036 31204
rect 45376 31152 45428 31204
rect 49148 31152 49200 31204
rect 78588 31152 78640 31204
rect 104164 31152 104216 31204
rect 114376 31152 114428 31204
rect 167644 31152 167696 31204
rect 212356 31152 212408 31204
rect 355324 31152 355376 31204
rect 5448 31084 5500 31136
rect 30380 31084 30432 31136
rect 31668 31084 31720 31136
rect 42432 31084 42484 31136
rect 82084 31084 82136 31136
rect 108304 31084 108356 31136
rect 112628 31084 112680 31136
rect 166264 31084 166316 31136
rect 168932 31084 168984 31136
rect 213184 31084 213236 31136
rect 222016 31084 222068 31136
rect 366364 31084 366416 31136
rect 4068 31016 4120 31068
rect 29644 31016 29696 31068
rect 30288 31016 30340 31068
rect 41880 31016 41932 31068
rect 67548 31016 67600 31068
rect 83004 31016 83056 31068
rect 85396 31016 85448 31068
rect 119344 31016 119396 31068
rect 121000 31016 121052 31068
rect 175924 31016 175976 31068
rect 180524 31016 180576 31068
rect 185492 31016 185544 31068
rect 228916 31016 228968 31068
rect 373264 31016 373316 31068
rect 23388 30948 23440 31000
rect 38660 30948 38712 31000
rect 39948 30948 40000 31000
rect 46296 30948 46348 31000
rect 119252 30948 119304 31000
rect 177396 30948 177448 31000
rect 192300 30948 192352 31000
rect 202328 30948 202380 31000
rect 344284 30948 344336 31000
rect 20628 30880 20680 30932
rect 36820 30880 36872 30932
rect 92296 30880 92348 30932
rect 135444 30880 135496 30932
rect 179972 30880 180024 30932
rect 195612 30880 195664 30932
rect 337384 30880 337436 30932
rect 22008 30812 22060 30864
rect 37924 30812 37976 30864
rect 90916 30812 90968 30864
rect 139952 30812 140004 30864
rect 181444 30812 181496 30864
rect 188436 30812 188488 30864
rect 188988 30812 189040 30864
rect 195060 30812 195112 30864
rect 195796 30812 195848 30864
rect 333244 30812 333296 30864
rect 24768 30744 24820 30796
rect 39120 30744 39172 30796
rect 102048 30744 102100 30796
rect 28816 30676 28868 30728
rect 41420 30676 41472 30728
rect 89628 30676 89680 30728
rect 129740 30676 129792 30728
rect 173164 30744 173216 30796
rect 185584 30744 185636 30796
rect 323676 30744 323728 30796
rect 142804 30676 142856 30728
rect 175188 30676 175240 30728
rect 301504 30676 301556 30728
rect 27528 30608 27580 30660
rect 40224 30608 40276 30660
rect 88156 30608 88208 30660
rect 127164 30608 127216 30660
rect 132500 30608 132552 30660
rect 136548 30608 136600 30660
rect 26148 30540 26200 30592
rect 39672 30540 39724 30592
rect 117688 30540 117740 30592
rect 128268 30540 128320 30592
rect 137928 30608 137980 30660
rect 177212 30608 177264 30660
rect 178960 30608 179012 30660
rect 181168 30540 181220 30592
rect 182088 30540 182140 30592
rect 183928 30540 183980 30592
rect 184848 30540 184900 30592
rect 187332 30540 187384 30592
rect 187608 30540 187660 30592
rect 203432 30540 203484 30592
rect 204076 30540 204128 30592
rect 210700 30540 210752 30592
rect 211068 30540 211120 30592
rect 224040 30540 224092 30592
rect 224868 30540 224920 30592
rect 227352 30540 227404 30592
rect 227628 30540 227680 30592
rect 232412 30540 232464 30592
rect 28908 30472 28960 30524
rect 40776 30472 40828 30524
rect 49608 30472 49660 30524
rect 51080 30472 51132 30524
rect 172244 30472 172296 30524
rect 244924 30472 244976 30524
rect 37096 30404 37148 30456
rect 45192 30404 45244 30456
rect 46848 30404 46900 30456
rect 49700 30404 49752 30456
rect 63132 30404 63184 30456
rect 63408 30404 63460 30456
rect 65892 30404 65944 30456
rect 66168 30404 66220 30456
rect 88708 30404 88760 30456
rect 93124 30404 93176 30456
rect 97080 30404 97132 30456
rect 97908 30404 97960 30456
rect 100300 30404 100352 30456
rect 100668 30404 100720 30456
rect 123852 30404 123904 30456
rect 124128 30404 124180 30456
rect 128820 30404 128872 30456
rect 129648 30404 129700 30456
rect 132132 30404 132184 30456
rect 132408 30404 132460 30456
rect 149428 30404 149480 30456
rect 150348 30404 150400 30456
rect 152740 30404 152792 30456
rect 153108 30404 153160 30456
rect 158352 30404 158404 30456
rect 158628 30404 158680 30456
rect 161112 30404 161164 30456
rect 161388 30404 161440 30456
rect 163320 30404 163372 30456
rect 164148 30404 164200 30456
rect 170588 30404 170640 30456
rect 242164 30404 242216 30456
rect 242440 30404 242492 30456
rect 250168 30472 250220 30524
rect 250996 30472 251048 30524
rect 251916 30472 251968 30524
rect 252468 30472 252520 30524
rect 253020 30472 253072 30524
rect 253572 30472 253624 30524
rect 254676 30472 254728 30524
rect 255136 30472 255188 30524
rect 255780 30472 255832 30524
rect 256516 30472 256568 30524
rect 257436 30472 257488 30524
rect 257988 30472 258040 30524
rect 259092 30472 259144 30524
rect 259276 30472 259328 30524
rect 260196 30472 260248 30524
rect 260748 30472 260800 30524
rect 261392 30472 261444 30524
rect 261944 30472 261996 30524
rect 263048 30472 263100 30524
rect 263508 30472 263560 30524
rect 264152 30472 264204 30524
rect 264704 30472 264756 30524
rect 266912 30472 266964 30524
rect 267556 30472 267608 30524
rect 268568 30472 268620 30524
rect 269028 30472 269080 30524
rect 269672 30608 269724 30660
rect 270500 30608 270552 30660
rect 276296 30608 276348 30660
rect 276388 30608 276440 30660
rect 277308 30608 277360 30660
rect 279700 30608 279752 30660
rect 280068 30608 280120 30660
rect 284760 30608 284812 30660
rect 285588 30608 285640 30660
rect 288072 30608 288124 30660
rect 288348 30608 288400 30660
rect 293132 30608 293184 30660
rect 293960 30608 294012 30660
rect 301412 30608 301464 30660
rect 308404 30608 308456 30660
rect 309784 30540 309836 30592
rect 270224 30472 270276 30524
rect 270408 30472 270460 30524
rect 271328 30472 271380 30524
rect 271788 30472 271840 30524
rect 272524 30472 272576 30524
rect 273076 30472 273128 30524
rect 273628 30472 273680 30524
rect 274456 30472 274508 30524
rect 275284 30472 275336 30524
rect 275928 30472 275980 30524
rect 276940 30472 276992 30524
rect 277216 30472 277268 30524
rect 278044 30472 278096 30524
rect 278688 30472 278740 30524
rect 279148 30472 279200 30524
rect 279884 30472 279936 30524
rect 280804 30472 280856 30524
rect 281356 30472 281408 30524
rect 281908 30472 281960 30524
rect 282736 30472 282788 30524
rect 283656 30472 283708 30524
rect 284208 30472 284260 30524
rect 285312 30472 285364 30524
rect 285496 30472 285548 30524
rect 286416 30472 286468 30524
rect 286968 30472 287020 30524
rect 287520 30472 287572 30524
rect 288164 30472 288216 30524
rect 289176 30472 289228 30524
rect 289636 30472 289688 30524
rect 290280 30472 290332 30524
rect 291016 30472 291068 30524
rect 291936 30472 291988 30524
rect 292396 30472 292448 30524
rect 293684 30472 293736 30524
rect 293868 30472 293920 30524
rect 294788 30472 294840 30524
rect 295248 30472 295300 30524
rect 295892 30472 295944 30524
rect 296444 30472 296496 30524
rect 298652 30472 298704 30524
rect 299296 30472 299348 30524
rect 301964 30472 302016 30524
rect 304264 30472 304316 30524
rect 245476 30404 245528 30456
rect 315396 30404 315448 30456
rect 37188 30336 37240 30388
rect 44640 30336 44692 30388
rect 48228 30336 48280 30388
rect 50252 30336 50304 30388
rect 52460 30336 52512 30388
rect 53012 30336 53064 30388
rect 54760 30336 54812 30388
rect 55128 30336 55180 30388
rect 55864 30336 55916 30388
rect 56416 30336 56468 30388
rect 56968 30336 57020 30388
rect 57796 30336 57848 30388
rect 58624 30336 58676 30388
rect 59176 30336 59228 30388
rect 59728 30336 59780 30388
rect 60648 30336 60700 30388
rect 61476 30336 61528 30388
rect 62028 30336 62080 30388
rect 62580 30336 62632 30388
rect 63224 30336 63276 30388
rect 64236 30336 64288 30388
rect 64696 30336 64748 30388
rect 65340 30336 65392 30388
rect 65984 30336 66036 30388
rect 66996 30336 67048 30388
rect 67548 30336 67600 30388
rect 68100 30336 68152 30388
rect 68928 30336 68980 30388
rect 69756 30336 69808 30388
rect 70308 30336 70360 30388
rect 71504 30336 71556 30388
rect 71688 30336 71740 30388
rect 73712 30336 73764 30388
rect 74356 30336 74408 30388
rect 76472 30336 76524 30388
rect 77116 30336 77168 30388
rect 78128 30336 78180 30388
rect 78588 30336 78640 30388
rect 79232 30336 79284 30388
rect 79876 30336 79928 30388
rect 80888 30336 80940 30388
rect 81348 30336 81400 30388
rect 85948 30336 86000 30388
rect 86776 30336 86828 30388
rect 87604 30336 87656 30388
rect 88248 30336 88300 30388
rect 91468 30336 91520 30388
rect 92296 30336 92348 30388
rect 93216 30336 93268 30388
rect 93768 30336 93820 30388
rect 94320 30336 94372 30388
rect 94872 30336 94924 30388
rect 95976 30336 96028 30388
rect 96436 30336 96488 30388
rect 97632 30336 97684 30388
rect 97816 30336 97868 30388
rect 98736 30336 98788 30388
rect 99288 30336 99340 30388
rect 99840 30336 99892 30388
rect 100576 30336 100628 30388
rect 101496 30336 101548 30388
rect 102048 30336 102100 30388
rect 102692 30336 102744 30388
rect 103244 30336 103296 30388
rect 105452 30336 105504 30388
rect 106188 30336 106240 30388
rect 107108 30336 107160 30388
rect 107568 30336 107620 30388
rect 108212 30336 108264 30388
rect 108764 30336 108816 30388
rect 113824 30336 113876 30388
rect 114468 30336 114520 30388
rect 114928 30336 114980 30388
rect 115756 30336 115808 30388
rect 116584 30336 116636 30388
rect 117136 30336 117188 30388
rect 120448 30336 120500 30388
rect 121368 30336 121420 30388
rect 122104 30336 122156 30388
rect 122748 30336 122800 30388
rect 123208 30336 123260 30388
rect 123944 30336 123996 30388
rect 124956 30336 125008 30388
rect 125416 30336 125468 30388
rect 126060 30336 126112 30388
rect 126796 30336 126848 30388
rect 127716 30336 127768 30388
rect 128268 30336 128320 30388
rect 129372 30336 129424 30388
rect 129556 30336 129608 30388
rect 130476 30336 130528 30388
rect 131028 30336 131080 30388
rect 131580 30336 131632 30388
rect 132224 30336 132276 30388
rect 133236 30336 133288 30388
rect 133696 30336 133748 30388
rect 134432 30336 134484 30388
rect 135076 30336 135128 30388
rect 136088 30336 136140 30388
rect 136548 30336 136600 30388
rect 137192 30336 137244 30388
rect 137928 30336 137980 30388
rect 140504 30336 140556 30388
rect 140688 30336 140740 30388
rect 141608 30336 141660 30388
rect 142068 30336 142120 30388
rect 142712 30336 142764 30388
rect 143264 30336 143316 30388
rect 143448 30336 143500 30388
rect 144368 30336 144420 30388
rect 144828 30336 144880 30388
rect 145564 30336 145616 30388
rect 146116 30336 146168 30388
rect 146668 30336 146720 30388
rect 147496 30336 147548 30388
rect 148324 30336 148376 30388
rect 148968 30336 149020 30388
rect 149980 30336 150032 30388
rect 150256 30336 150308 30388
rect 151084 30336 151136 30388
rect 151728 30336 151780 30388
rect 152188 30336 152240 30388
rect 152924 30336 152976 30388
rect 153844 30336 153896 30388
rect 154396 30336 154448 30388
rect 154948 30336 155000 30388
rect 155776 30336 155828 30388
rect 156696 30336 156748 30388
rect 157248 30336 157300 30388
rect 157800 30336 157852 30388
rect 158444 30336 158496 30388
rect 159456 30336 159508 30388
rect 159916 30336 159968 30388
rect 160560 30336 160612 30388
rect 161204 30336 161256 30388
rect 163872 30336 163924 30388
rect 164056 30336 164108 30388
rect 164976 30336 165028 30388
rect 165528 30336 165580 30388
rect 166172 30336 166224 30388
rect 166908 30336 166960 30388
rect 171692 30336 171744 30388
rect 172428 30336 172480 30388
rect 173348 30336 173400 30388
rect 173808 30336 173860 30388
rect 174452 30336 174504 30388
rect 175004 30336 175056 30388
rect 177304 30336 177356 30388
rect 177856 30336 177908 30388
rect 178408 30336 178460 30388
rect 179236 30336 179288 30388
rect 180064 30336 180116 30388
rect 180708 30336 180760 30388
rect 181720 30336 181772 30388
rect 181996 30336 182048 30388
rect 182824 30336 182876 30388
rect 183468 30336 183520 30388
rect 184480 30336 184532 30388
rect 184756 30336 184808 30388
rect 186688 30336 186740 30388
rect 187424 30336 187476 30388
rect 189540 30336 189592 30388
rect 190276 30336 190328 30388
rect 191196 30336 191248 30388
rect 191748 30336 191800 30388
rect 192852 30336 192904 30388
rect 193128 30336 193180 30388
rect 193956 30336 194008 30388
rect 194508 30336 194560 30388
rect 196716 30336 196768 30388
rect 197176 30336 197228 30388
rect 197912 30336 197964 30388
rect 198648 30336 198700 30388
rect 199568 30336 199620 30388
rect 200028 30336 200080 30388
rect 200672 30336 200724 30388
rect 143448 30200 143500 30252
rect 201224 30336 201276 30388
rect 201408 30336 201460 30388
rect 203892 30336 203944 30388
rect 204168 30336 204220 30388
rect 205088 30336 205140 30388
rect 205548 30336 205600 30388
rect 206192 30336 206244 30388
rect 206744 30336 206796 30388
rect 210148 30336 210200 30388
rect 210884 30336 210936 30388
rect 211804 30336 211856 30388
rect 212448 30336 212500 30388
rect 212908 30336 212960 30388
rect 213736 30336 213788 30388
rect 214564 30336 214616 30388
rect 215208 30336 215260 30388
rect 216220 30336 216272 30388
rect 216588 30336 216640 30388
rect 217324 30336 217376 30388
rect 217968 30336 218020 30388
rect 218428 30336 218480 30388
rect 219256 30336 219308 30388
rect 220176 30336 220228 30388
rect 220636 30336 220688 30388
rect 221280 30336 221332 30388
rect 222108 30336 222160 30388
rect 222936 30336 222988 30388
rect 223488 30336 223540 30388
rect 224592 30336 224644 30388
rect 224776 30336 224828 30388
rect 226800 30336 226852 30388
rect 227444 30336 227496 30388
rect 228456 30336 228508 30388
rect 229008 30336 229060 30388
rect 229652 30336 229704 30388
rect 230296 30336 230348 30388
rect 231308 30336 231360 30388
rect 231768 30336 231820 30388
rect 232964 30336 233016 30388
rect 233148 30336 233200 30388
rect 235172 30336 235224 30388
rect 235816 30336 235868 30388
rect 235724 30268 235776 30320
rect 239588 30336 239640 30388
rect 240048 30336 240100 30388
rect 240784 30336 240836 30388
rect 241336 30336 241388 30388
rect 241888 30336 241940 30388
rect 242716 30336 242768 30388
rect 243544 30336 243596 30388
rect 244188 30336 244240 30388
rect 244648 30336 244700 30388
rect 245568 30336 245620 30388
rect 246304 30336 246356 30388
rect 246948 30336 247000 30388
rect 247408 30336 247460 30388
rect 248144 30336 248196 30388
rect 312544 30336 312596 30388
rect 201408 30200 201460 30252
rect 296628 30200 296680 30252
rect 296536 29996 296588 30048
rect 258540 27276 258592 27328
rect 259368 27276 259420 27328
rect 302884 20612 302936 20664
rect 579988 20612 580040 20664
rect 234436 16056 234488 16108
rect 436744 16056 436796 16108
rect 241336 15988 241388 16040
rect 450912 15988 450964 16040
rect 244096 15920 244148 15972
rect 456800 15920 456852 15972
rect 248144 15852 248196 15904
rect 465172 15852 465224 15904
rect 227444 15104 227496 15156
rect 420920 15104 420972 15156
rect 229008 15036 229060 15088
rect 423680 15036 423732 15088
rect 230204 14968 230256 15020
rect 428464 14968 428516 15020
rect 231676 14900 231728 14952
rect 432052 14900 432104 14952
rect 233056 14832 233108 14884
rect 435088 14832 435140 14884
rect 248236 14764 248288 14816
rect 465816 14764 465868 14816
rect 249708 14696 249760 14748
rect 469864 14696 469916 14748
rect 253664 14628 253716 14680
rect 476488 14628 476540 14680
rect 250904 14560 250956 14612
rect 473452 14560 473504 14612
rect 290924 14492 290976 14544
rect 556896 14492 556948 14544
rect 292396 14424 292448 14476
rect 559288 14424 559340 14476
rect 208216 14356 208268 14408
rect 381176 14356 381228 14408
rect 206744 14288 206796 14340
rect 377680 14288 377732 14340
rect 184664 14220 184716 14272
rect 332692 14220 332744 14272
rect 187424 14152 187476 14204
rect 336280 14152 336332 14204
rect 183376 14084 183428 14136
rect 328736 14084 328788 14136
rect 181904 14016 181956 14068
rect 326344 14016 326396 14068
rect 181996 13948 182048 14000
rect 324320 13948 324372 14000
rect 177856 13880 177908 13932
rect 316040 13880 316092 13932
rect 173716 13812 173768 13864
rect 307760 13812 307812 13864
rect 257896 13744 257948 13796
rect 487160 13744 487212 13796
rect 259184 13676 259236 13728
rect 489920 13676 489972 13728
rect 261944 13608 261996 13660
rect 494704 13608 494756 13660
rect 275836 13540 275888 13592
rect 525432 13540 525484 13592
rect 277124 13472 277176 13524
rect 528560 13472 528612 13524
rect 158444 13404 158496 13456
rect 274824 13404 274876 13456
rect 279884 13404 279936 13456
rect 532056 13404 532108 13456
rect 159916 13336 159968 13388
rect 278320 13336 278372 13388
rect 281356 13336 281408 13388
rect 536104 13336 536156 13388
rect 162768 13268 162820 13320
rect 284944 13268 284996 13320
rect 285404 13268 285456 13320
rect 546684 13268 546736 13320
rect 163964 13200 164016 13252
rect 288992 13200 289044 13252
rect 289636 13200 289688 13252
rect 553768 13200 553820 13252
rect 169576 13132 169628 13184
rect 299664 13132 299716 13184
rect 300676 13132 300728 13184
rect 576952 13132 577004 13184
rect 171048 13064 171100 13116
rect 303160 13064 303212 13116
rect 304264 13064 304316 13116
rect 581736 13064 581788 13116
rect 256424 12996 256476 13048
rect 484032 12996 484084 13048
rect 255136 12928 255188 12980
rect 480536 12928 480588 12980
rect 203984 12860 204036 12912
rect 374092 12860 374144 12912
rect 202788 12792 202840 12844
rect 370136 12792 370188 12844
rect 177948 12724 178000 12776
rect 317328 12724 317380 12776
rect 176476 12656 176528 12708
rect 313832 12656 313884 12708
rect 172336 12588 172388 12640
rect 306380 12588 306432 12640
rect 175096 12520 175148 12572
rect 309692 12520 309744 12572
rect 168196 12452 168248 12504
rect 295616 12452 295668 12504
rect 296444 12452 296496 12504
rect 418804 12452 418856 12504
rect 250996 12384 251048 12436
rect 470600 12384 470652 12436
rect 252468 12316 252520 12368
rect 474096 12316 474148 12368
rect 253756 12248 253808 12300
rect 478144 12248 478196 12300
rect 256516 12180 256568 12232
rect 482376 12180 482428 12232
rect 257988 12112 258040 12164
rect 486424 12112 486476 12164
rect 259276 12044 259328 12096
rect 490012 12044 490064 12096
rect 260656 11976 260708 12028
rect 493048 11976 493100 12028
rect 262036 11908 262088 11960
rect 497096 11908 497148 11960
rect 264704 11840 264756 11892
rect 500592 11840 500644 11892
rect 266176 11772 266228 11824
rect 503720 11772 503772 11824
rect 267464 11704 267516 11756
rect 507216 11704 507268 11756
rect 248328 11636 248380 11688
rect 467472 11636 467524 11688
rect 246856 11568 246908 11620
rect 463976 11568 464028 11620
rect 245476 11500 245528 11552
rect 459928 11500 459980 11552
rect 244188 11432 244240 11484
rect 456892 11432 456944 11484
rect 242716 11364 242768 11416
rect 453304 11364 453356 11416
rect 239956 11296 240008 11348
rect 448520 11296 448572 11348
rect 238576 11228 238628 11280
rect 445760 11228 445812 11280
rect 235816 11160 235868 11212
rect 439136 11160 439188 11212
rect 164056 11092 164108 11144
rect 287336 11092 287388 11144
rect 201224 10956 201276 11008
rect 367744 10956 367796 11008
rect 204076 10888 204128 10940
rect 371240 10888 371292 10940
rect 205548 10820 205600 10872
rect 375288 10820 375340 10872
rect 206836 10752 206888 10804
rect 378416 10752 378468 10804
rect 208308 10684 208360 10736
rect 382372 10684 382424 10736
rect 210884 10616 210936 10668
rect 385960 10616 386012 10668
rect 212448 10548 212500 10600
rect 389456 10548 389508 10600
rect 213644 10480 213696 10532
rect 392584 10480 392636 10532
rect 215116 10412 215168 10464
rect 396080 10412 396132 10464
rect 216496 10344 216548 10396
rect 398840 10344 398892 10396
rect 219256 10276 219308 10328
rect 403624 10276 403676 10328
rect 199936 10208 199988 10260
rect 364616 10208 364668 10260
rect 198556 10140 198608 10192
rect 361120 10140 361172 10192
rect 197176 10072 197228 10124
rect 357532 10072 357584 10124
rect 195796 10004 195848 10056
rect 353576 10004 353628 10056
rect 193036 9936 193088 9988
rect 349160 9936 349212 9988
rect 191656 9868 191708 9920
rect 346952 9868 347004 9920
rect 190184 9800 190236 9852
rect 342904 9800 342956 9852
rect 188988 9732 189040 9784
rect 339500 9732 339552 9784
rect 244924 9664 244976 9716
rect 305552 9664 305604 9716
rect 157156 9596 157208 9648
rect 273628 9596 273680 9648
rect 274456 9596 274508 9648
rect 520740 9596 520792 9648
rect 158536 9528 158588 9580
rect 277124 9528 277176 9580
rect 277216 9528 277268 9580
rect 527824 9528 527876 9580
rect 160008 9460 160060 9512
rect 279516 9460 279568 9512
rect 161204 9392 161256 9444
rect 280712 9460 280764 9512
rect 282736 9460 282788 9512
rect 279976 9392 280028 9444
rect 164148 9324 164200 9376
rect 161296 9256 161348 9308
rect 283104 9256 283156 9308
rect 284208 9392 284260 9444
rect 534908 9460 534960 9512
rect 286600 9324 286652 9376
rect 538404 9392 538456 9444
rect 541992 9324 542044 9376
rect 286876 9256 286928 9308
rect 549076 9256 549128 9308
rect 165528 9188 165580 9240
rect 290188 9188 290240 9240
rect 293776 9188 293828 9240
rect 563244 9188 563296 9240
rect 166816 9120 166868 9172
rect 293684 9120 293736 9172
rect 295156 9120 295208 9172
rect 566832 9120 566884 9172
rect 173808 9052 173860 9104
rect 307944 9052 307996 9104
rect 308404 9052 308456 9104
rect 581000 9052 581052 9104
rect 168288 8984 168340 9036
rect 297272 8984 297324 9036
rect 299296 8984 299348 9036
rect 300676 8984 300728 9036
rect 169668 8916 169720 8968
rect 300768 8916 300820 8968
rect 573916 8984 573968 9036
rect 578608 8916 578660 8968
rect 155684 8848 155736 8900
rect 270040 8848 270092 8900
rect 270316 8848 270368 8900
rect 513564 8848 513616 8900
rect 154396 8780 154448 8832
rect 266544 8780 266596 8832
rect 267556 8780 267608 8832
rect 506480 8780 506532 8832
rect 150164 8712 150216 8764
rect 259460 8712 259512 8764
rect 262128 8712 262180 8764
rect 152924 8644 152976 8696
rect 262956 8644 263008 8696
rect 263416 8712 263468 8764
rect 499396 8712 499448 8764
rect 495900 8644 495952 8696
rect 148876 8576 148928 8628
rect 255872 8576 255924 8628
rect 259368 8576 259420 8628
rect 488816 8576 488868 8628
rect 147404 8508 147456 8560
rect 252376 8508 252428 8560
rect 256608 8508 256660 8560
rect 485228 8508 485280 8560
rect 146116 8440 146168 8492
rect 248788 8440 248840 8492
rect 255228 8440 255280 8492
rect 481732 8440 481784 8492
rect 175188 8372 175240 8424
rect 311440 8372 311492 8424
rect 172428 8304 172480 8356
rect 304356 8304 304408 8356
rect 223488 8236 223540 8288
rect 413100 8236 413152 8288
rect 123944 8168 123996 8220
rect 201500 8168 201552 8220
rect 224776 8168 224828 8220
rect 416688 8168 416740 8220
rect 125416 8100 125468 8152
rect 205088 8100 205140 8152
rect 226248 8100 226300 8152
rect 420184 8100 420236 8152
rect 126704 8032 126756 8084
rect 208584 8032 208636 8084
rect 230296 8032 230348 8084
rect 427268 8032 427320 8084
rect 132224 7964 132276 8016
rect 219256 7964 219308 8016
rect 227536 7964 227588 8016
rect 423772 7964 423824 8016
rect 129464 7896 129516 7948
rect 215668 7896 215720 7948
rect 231768 7896 231820 7948
rect 430856 7896 430908 7948
rect 133696 7828 133748 7880
rect 222752 7828 222804 7880
rect 233148 7828 233200 7880
rect 434444 7828 434496 7880
rect 134984 7760 135036 7812
rect 226340 7760 226392 7812
rect 234528 7760 234580 7812
rect 437940 7760 437992 7812
rect 139216 7692 139268 7744
rect 234620 7692 234672 7744
rect 235908 7692 235960 7744
rect 441528 7692 441580 7744
rect 141976 7624 142028 7676
rect 241704 7624 241756 7676
rect 242808 7624 242860 7676
rect 455696 7624 455748 7676
rect 143264 7556 143316 7608
rect 245200 7556 245252 7608
rect 245568 7556 245620 7608
rect 459192 7556 459244 7608
rect 222108 7488 222160 7540
rect 409604 7488 409656 7540
rect 219348 7420 219400 7472
rect 406016 7420 406068 7472
rect 217876 7352 217928 7404
rect 402520 7352 402572 7404
rect 216588 7284 216640 7336
rect 398932 7284 398984 7336
rect 215208 7216 215260 7268
rect 395344 7216 395396 7268
rect 213736 7148 213788 7200
rect 391848 7148 391900 7200
rect 210976 7080 211028 7132
rect 388260 7080 388312 7132
rect 209688 7012 209740 7064
rect 384764 7012 384816 7064
rect 158628 6944 158680 6996
rect 276020 6944 276072 6996
rect 276664 6944 276716 6996
rect 319720 6944 319772 6996
rect 142068 6808 142120 6860
rect 240508 6808 240560 6860
rect 242164 6808 242216 6860
rect 301412 6808 301464 6860
rect 301504 6808 301556 6860
rect 312636 6808 312688 6860
rect 315304 6808 315356 6860
rect 580172 6808 580224 6860
rect 117136 6740 117188 6792
rect 187332 6740 187384 6792
rect 198648 6740 198700 6792
rect 359924 6740 359976 6792
rect 118516 6672 118568 6724
rect 190828 6672 190880 6724
rect 200028 6672 200080 6724
rect 363512 6672 363564 6724
rect 119988 6604 120040 6656
rect 194324 6604 194376 6656
rect 201316 6604 201368 6656
rect 367008 6604 367060 6656
rect 121276 6536 121328 6588
rect 197912 6536 197964 6588
rect 237196 6536 237248 6588
rect 442632 6536 442684 6588
rect 143356 6468 143408 6520
rect 244096 6468 244148 6520
rect 260748 6468 260800 6520
rect 492312 6468 492364 6520
rect 144736 6400 144788 6452
rect 247592 6400 247644 6452
rect 264796 6400 264848 6452
rect 502984 6400 503036 6452
rect 147496 6332 147548 6384
rect 251180 6332 251232 6384
rect 269028 6332 269080 6384
rect 510068 6332 510120 6384
rect 99196 6264 99248 6316
rect 150624 6264 150676 6316
rect 151636 6264 151688 6316
rect 261760 6264 261812 6316
rect 271696 6264 271748 6316
rect 517152 6264 517204 6316
rect 100484 6196 100536 6248
rect 154212 6196 154264 6248
rect 155776 6196 155828 6248
rect 268844 6196 268896 6248
rect 275928 6196 275980 6248
rect 524236 6196 524288 6248
rect 111616 6128 111668 6180
rect 176660 6128 176712 6180
rect 179328 6128 179380 6180
rect 320916 6128 320968 6180
rect 322204 6128 322256 6180
rect 115756 6060 115808 6112
rect 183744 6060 183796 6112
rect 194416 6060 194468 6112
rect 352840 6060 352892 6112
rect 113088 5992 113140 6044
rect 180248 5992 180300 6044
rect 193128 5992 193180 6044
rect 349252 5992 349304 6044
rect 114468 5924 114520 5976
rect 181444 5924 181496 5976
rect 191748 5924 191800 5976
rect 345756 5924 345808 5976
rect 110236 5856 110288 5908
rect 173164 5856 173216 5908
rect 190276 5856 190328 5908
rect 342168 5856 342220 5908
rect 108948 5788 109000 5840
rect 170772 5788 170824 5840
rect 187516 5788 187568 5840
rect 338672 5788 338724 5840
rect 108856 5720 108908 5772
rect 169576 5720 169628 5772
rect 186228 5720 186280 5772
rect 335084 5720 335136 5772
rect 106096 5652 106148 5704
rect 166080 5652 166132 5704
rect 184756 5652 184808 5704
rect 331588 5652 331640 5704
rect 104808 5584 104860 5636
rect 162492 5584 162544 5636
rect 183468 5584 183520 5636
rect 328000 5584 328052 5636
rect 103244 5516 103296 5568
rect 157800 5516 157852 5568
rect 182088 5516 182140 5568
rect 324412 5516 324464 5568
rect 93768 5448 93820 5500
rect 137652 5448 137704 5500
rect 137836 5448 137888 5500
rect 232228 5448 232280 5500
rect 278688 5448 278740 5500
rect 530124 5448 530176 5500
rect 94964 5380 95016 5432
rect 140044 5380 140096 5432
rect 140596 5380 140648 5432
rect 239312 5380 239364 5432
rect 274548 5380 274600 5432
rect 280068 5380 280120 5432
rect 533712 5380 533764 5432
rect 95056 5312 95108 5364
rect 141240 5312 141292 5364
rect 143448 5312 143500 5364
rect 242900 5312 242952 5364
rect 277308 5312 277360 5364
rect 282828 5312 282880 5364
rect 96528 5244 96580 5296
rect 144736 5244 144788 5296
rect 144828 5244 144880 5296
rect 246396 5244 246448 5296
rect 284300 5244 284352 5296
rect 285588 5244 285640 5296
rect 537208 5312 537260 5364
rect 96436 5176 96488 5228
rect 143540 5176 143592 5228
rect 146208 5176 146260 5228
rect 249984 5176 250036 5228
rect 281908 5176 281960 5228
rect 288348 5176 288400 5228
rect 291660 5176 291712 5228
rect 540796 5244 540848 5296
rect 544384 5176 544436 5228
rect 97816 5108 97868 5160
rect 147128 5108 147180 5160
rect 147588 5108 147640 5160
rect 253480 5108 253532 5160
rect 271788 5108 271840 5160
rect 286968 5108 287020 5160
rect 547880 5108 547932 5160
rect 97724 5040 97776 5092
rect 148324 5040 148376 5092
rect 150348 5040 150400 5092
rect 257068 5040 257120 5092
rect 264888 5040 264940 5092
rect 273168 5040 273220 5092
rect 100576 4972 100628 5024
rect 151820 4972 151872 5024
rect 153108 4972 153160 5024
rect 264152 4972 264204 5024
rect 266268 4972 266320 5024
rect 281448 4972 281500 5024
rect 102048 4904 102100 4956
rect 155408 4904 155460 4956
rect 155868 4904 155920 4956
rect 271236 4904 271288 4956
rect 291936 5040 291988 5092
rect 551468 5040 551520 5092
rect 295248 4972 295300 5024
rect 103336 4836 103388 4888
rect 158904 4836 158956 4888
rect 161388 4836 161440 4888
rect 291384 4836 291436 4888
rect 298468 4904 298520 4956
rect 299388 4904 299440 4956
rect 562048 4972 562100 5024
rect 565636 4904 565688 4956
rect 294880 4836 294932 4888
rect 296628 4836 296680 4888
rect 569132 4836 569184 4888
rect 106188 4768 106240 4820
rect 163688 4768 163740 4820
rect 166908 4768 166960 4820
rect 92296 4700 92348 4752
rect 134156 4700 134208 4752
rect 136548 4700 136600 4752
rect 228732 4700 228784 4752
rect 292580 4768 292632 4820
rect 293868 4768 293920 4820
rect 576308 4768 576360 4820
rect 523040 4700 523092 4752
rect 89628 4632 89680 4684
rect 129372 4632 129424 4684
rect 135076 4632 135128 4684
rect 225144 4632 225196 4684
rect 263508 4632 263560 4684
rect 526628 4632 526680 4684
rect 88248 4564 88300 4616
rect 125876 4564 125928 4616
rect 132316 4564 132368 4616
rect 221556 4564 221608 4616
rect 130936 4496 130988 4548
rect 218060 4496 218112 4548
rect 124036 4428 124088 4480
rect 203892 4428 203944 4480
rect 204904 4428 204956 4480
rect 519544 4564 519596 4616
rect 515956 4496 516008 4548
rect 267648 4428 267700 4480
rect 128268 4360 128320 4412
rect 210976 4360 211028 4412
rect 213184 4360 213236 4412
rect 270408 4428 270460 4480
rect 512460 4428 512512 4480
rect 508872 4360 508924 4412
rect 126796 4292 126848 4344
rect 207388 4292 207440 4344
rect 209044 4292 209096 4344
rect 505376 4292 505428 4344
rect 129556 4224 129608 4276
rect 214472 4224 214524 4276
rect 63316 4088 63368 4140
rect 75000 4088 75052 4140
rect 77208 4088 77260 4140
rect 104532 4088 104584 4140
rect 110328 4156 110380 4208
rect 122656 4156 122708 4208
rect 200304 4156 200356 4208
rect 200764 4156 200816 4208
rect 501788 4224 501840 4276
rect 498200 4156 498252 4208
rect 65984 4020 66036 4072
rect 78588 4020 78640 4072
rect 79876 4020 79928 4072
rect 108120 4020 108172 4072
rect 29092 3952 29144 4004
rect 60648 3952 60700 4004
rect 66720 3952 66772 4004
rect 67548 3952 67600 4004
rect 81348 3952 81400 4004
rect 111616 4088 111668 4140
rect 117964 4088 118016 4140
rect 115204 4020 115256 4072
rect 115848 4020 115900 4072
rect 184940 4088 184992 4140
rect 185584 4088 185636 4140
rect 201408 4088 201460 4140
rect 365812 4088 365864 4140
rect 366364 4088 366416 4140
rect 121368 4020 121420 4072
rect 114008 3952 114060 4004
rect 117228 3952 117280 4004
rect 117964 3952 118016 4004
rect 123484 3952 123536 4004
rect 124128 3952 124180 4004
rect 127440 3952 127492 4004
rect 188528 4020 188580 4072
rect 204168 4020 204220 4072
rect 372896 4020 372948 4072
rect 383476 4088 383528 4140
rect 433248 4088 433300 4140
rect 376484 4020 376536 4072
rect 376576 4020 376628 4072
rect 195612 3952 195664 4004
rect 206192 3952 206244 4004
rect 206928 3952 206980 4004
rect 379980 3952 380032 4004
rect 380164 4020 380216 4072
rect 447416 4020 447468 4072
rect 382924 3952 382976 4004
rect 475752 3952 475804 4004
rect 30564 3884 30616 3936
rect 64788 3884 64840 3936
rect 77392 3884 77444 3936
rect 79784 3884 79836 3936
rect 109316 3884 109368 3936
rect 119896 3884 119948 3936
rect 122748 3884 122800 3936
rect 17040 3816 17092 3868
rect 19432 3748 19484 3800
rect 20536 3748 20588 3800
rect 66168 3816 66220 3868
rect 79692 3816 79744 3868
rect 81256 3816 81308 3868
rect 112812 3816 112864 3868
rect 118608 3816 118660 3868
rect 192024 3884 192076 3936
rect 194508 3884 194560 3936
rect 211068 3884 211120 3936
rect 387156 3884 387208 3936
rect 36084 3748 36136 3800
rect 70216 3748 70268 3800
rect 12256 3680 12308 3732
rect 33324 3680 33376 3732
rect 62028 3680 62080 3732
rect 70308 3680 70360 3732
rect 80888 3748 80940 3800
rect 82084 3748 82136 3800
rect 82728 3748 82780 3800
rect 108396 3748 108448 3800
rect 124680 3748 124732 3800
rect 125508 3748 125560 3800
rect 199108 3816 199160 3868
rect 127808 3748 127860 3800
rect 202696 3816 202748 3868
rect 213828 3816 213880 3868
rect 394240 3816 394292 3868
rect 89168 3680 89220 3732
rect 7656 3612 7708 3664
rect 2872 3544 2924 3596
rect 1676 3476 1728 3528
rect 27804 3612 27856 3664
rect 60464 3612 60516 3664
rect 68928 3612 68980 3664
rect 84476 3612 84528 3664
rect 86868 3612 86920 3664
rect 87604 3612 87656 3664
rect 93124 3680 93176 3732
rect 128176 3680 128228 3732
rect 27712 3544 27764 3596
rect 28816 3544 28868 3596
rect 35992 3544 36044 3596
rect 37096 3544 37148 3596
rect 44272 3544 44324 3596
rect 45376 3544 45428 3596
rect 60556 3544 60608 3596
rect 69112 3544 69164 3596
rect 71596 3544 71648 3596
rect 92756 3544 92808 3596
rect 122288 3612 122340 3664
rect 126888 3612 126940 3664
rect 129648 3612 129700 3664
rect 209780 3748 209832 3800
rect 217968 3748 218020 3800
rect 401324 3816 401376 3868
rect 398840 3748 398892 3800
rect 400128 3748 400180 3800
rect 220728 3680 220780 3732
rect 408408 3680 408460 3732
rect 93952 3544 94004 3596
rect 94504 3544 94556 3596
rect 131764 3544 131816 3596
rect 212172 3612 212224 3664
rect 224868 3612 224920 3664
rect 415492 3612 415544 3664
rect 418804 3612 418856 3664
rect 568028 3612 568080 3664
rect 213368 3544 213420 3596
rect 227628 3544 227680 3596
rect 422576 3544 422628 3596
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 52460 3476 52512 3528
rect 53748 3476 53800 3528
rect 54024 3476 54076 3528
rect 54944 3476 54996 3528
rect 56416 3476 56468 3528
rect 58440 3476 58492 3528
rect 59176 3476 59228 3528
rect 64328 3476 64380 3528
rect 67916 3476 67968 3528
rect 70400 3476 70452 3528
rect 85672 3476 85724 3528
rect 86776 3476 86828 3528
rect 88984 3476 89036 3528
rect 90364 3476 90416 3528
rect 119344 3476 119396 3528
rect 121092 3476 121144 3528
rect 132408 3476 132460 3528
rect 220452 3476 220504 3528
rect 230388 3476 230440 3528
rect 429660 3544 429712 3596
rect 489920 3544 489972 3596
rect 491116 3544 491168 3596
rect 423680 3476 423732 3528
rect 424968 3476 425020 3528
rect 448520 3476 448572 3528
rect 449808 3476 449860 3528
rect 456800 3476 456852 3528
rect 458088 3476 458140 3528
rect 572 3408 624 3460
rect 27620 3408 27672 3460
rect 57796 3408 57848 3460
rect 60832 3408 60884 3460
rect 61936 3408 61988 3460
rect 71504 3408 71556 3460
rect 71688 3408 71740 3460
rect 91560 3408 91612 3460
rect 92388 3408 92440 3460
rect 135260 3408 135312 3460
rect 137928 3408 137980 3460
rect 231032 3408 231084 3460
rect 237288 3408 237340 3460
rect 443828 3408 443880 3460
rect 8760 3340 8812 3392
rect 9588 3340 9640 3392
rect 9956 3340 10008 3392
rect 10968 3340 11020 3392
rect 11152 3340 11204 3392
rect 12348 3340 12400 3392
rect 15936 3340 15988 3392
rect 16488 3340 16540 3392
rect 18236 3340 18288 3392
rect 19248 3340 19300 3392
rect 24216 3340 24268 3392
rect 24768 3340 24820 3392
rect 25320 3340 25372 3392
rect 26148 3340 26200 3392
rect 57888 3340 57940 3392
rect 63224 3340 63276 3392
rect 64696 3340 64748 3392
rect 76196 3340 76248 3392
rect 78496 3340 78548 3392
rect 55128 3272 55180 3324
rect 56048 3272 56100 3324
rect 66076 3272 66128 3324
rect 87972 3272 88024 3324
rect 90456 3272 90508 3324
rect 57704 3204 57756 3256
rect 62028 3204 62080 3256
rect 63408 3204 63460 3256
rect 73804 3204 73856 3256
rect 77116 3204 77168 3256
rect 102232 3204 102284 3256
rect 104164 3340 104216 3392
rect 106924 3340 106976 3392
rect 105728 3204 105780 3256
rect 105820 3204 105872 3256
rect 111708 3340 111760 3392
rect 177856 3340 177908 3392
rect 116400 3272 116452 3324
rect 107568 3204 107620 3256
rect 174268 3272 174320 3324
rect 177396 3272 177448 3324
rect 193220 3272 193272 3324
rect 167184 3204 167236 3256
rect 175924 3204 175976 3256
rect 55036 3136 55088 3188
rect 57244 3136 57296 3188
rect 63316 3136 63368 3188
rect 72608 3136 72660 3188
rect 75828 3136 75880 3188
rect 101036 3136 101088 3188
rect 101404 3136 101456 3188
rect 103612 3136 103664 3188
rect 160100 3136 160152 3188
rect 160744 3136 160796 3188
rect 56508 3068 56560 3120
rect 59636 3068 59688 3120
rect 68836 3068 68888 3120
rect 75736 3068 75788 3120
rect 99840 3068 99892 3120
rect 74448 3000 74500 3052
rect 98644 3000 98696 3052
rect 74264 2932 74316 2984
rect 97448 2932 97500 2984
rect 100668 3000 100720 3052
rect 153016 3068 153068 3120
rect 155224 3068 155276 3120
rect 161296 3068 161348 3120
rect 170404 3136 170456 3188
rect 189724 3136 189776 3188
rect 190368 3136 190420 3188
rect 197268 3272 197320 3324
rect 355968 3340 356020 3392
rect 349160 3272 349212 3324
rect 350448 3272 350500 3324
rect 351184 3272 351236 3324
rect 344560 3204 344612 3256
rect 351644 3204 351696 3256
rect 351828 3272 351880 3324
rect 358084 3340 358136 3392
rect 369492 3340 369544 3392
rect 373264 3340 373316 3392
rect 426164 3340 426216 3392
rect 355876 3204 355928 3256
rect 383476 3272 383528 3324
rect 383568 3272 383620 3324
rect 418988 3272 419040 3324
rect 337476 3136 337528 3188
rect 337568 3136 337620 3188
rect 344284 3136 344336 3188
rect 369400 3204 369452 3256
rect 411904 3204 411956 3256
rect 404820 3136 404872 3188
rect 175464 3068 175516 3120
rect 177304 3068 177356 3120
rect 181536 3068 181588 3120
rect 237012 3068 237064 3120
rect 307760 3068 307812 3120
rect 309048 3068 309100 3120
rect 309784 3068 309836 3120
rect 461584 3068 461636 3120
rect 583392 3111 583444 3120
rect 583392 3077 583401 3111
rect 583401 3077 583435 3111
rect 583435 3077 583444 3111
rect 583392 3068 583444 3077
rect 59268 2864 59320 2916
rect 65524 2864 65576 2916
rect 73068 2864 73120 2916
rect 95148 2864 95200 2916
rect 95884 2864 95936 2916
rect 74356 2796 74408 2848
rect 96252 2796 96304 2848
rect 99288 2932 99340 2984
rect 149520 3000 149572 3052
rect 156604 3000 156656 3052
rect 164884 3000 164936 3052
rect 167644 3000 167696 3052
rect 182548 3000 182600 3052
rect 184848 3000 184900 3052
rect 145932 2932 145984 2984
rect 166264 2932 166316 2984
rect 179052 2932 179104 2984
rect 180064 2932 180116 2984
rect 142436 2864 142488 2916
rect 142804 2864 142856 2916
rect 156604 2864 156656 2916
rect 157984 2864 158036 2916
rect 168380 2864 168432 2916
rect 169024 2864 169076 2916
rect 186136 2864 186188 2916
rect 187608 3000 187660 3052
rect 330392 3000 330444 3052
rect 330484 3000 330536 3052
rect 333244 3000 333296 3052
rect 348056 3000 348108 3052
rect 362316 3000 362368 3052
rect 362408 3000 362460 3052
rect 397736 3000 397788 3052
rect 233424 2932 233476 2984
rect 315396 2932 315448 2984
rect 454500 2932 454552 2984
rect 196808 2864 196860 2916
rect 323308 2864 323360 2916
rect 323676 2864 323728 2916
rect 333888 2864 333940 2916
rect 95240 2728 95292 2780
rect 97908 2796 97960 2848
rect 138848 2796 138900 2848
rect 159364 2796 159416 2848
rect 171968 2796 172020 2848
rect 173256 2796 173308 2848
rect 229836 2796 229888 2848
rect 312544 2796 312596 2848
rect 324320 2728 324372 2780
rect 325608 2728 325660 2780
rect 340972 2864 341024 2916
rect 341524 2864 341576 2916
rect 355232 2864 355284 2916
rect 355324 2864 355376 2916
rect 358728 2864 358780 2916
rect 390652 2864 390704 2916
rect 440332 2796 440384 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3148 593360 3200 593366
rect 3148 593302 3200 593308
rect 3160 593065 3188 593302
rect 3146 593056 3202 593065
rect 3146 592991 3202 593000
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3332 540932 3384 540938
rect 3332 540874 3384 540880
rect 3344 540841 3372 540874
rect 3330 540832 3386 540841
rect 3330 540767 3386 540776
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3148 489864 3200 489870
rect 3148 489806 3200 489812
rect 3160 488753 3188 489806
rect 3146 488744 3202 488753
rect 3146 488679 3202 488688
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 3332 437436 3384 437442
rect 3332 437378 3384 437384
rect 3344 436665 3372 437378
rect 3330 436656 3386 436665
rect 3330 436591 3386 436600
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422346 3188 423535
rect 3148 422340 3200 422346
rect 3148 422282 3200 422288
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3436 314498 3464 658135
rect 4804 650072 4856 650078
rect 4804 650014 4856 650020
rect 3792 644496 3844 644502
rect 3792 644438 3844 644444
rect 3698 644328 3754 644337
rect 3698 644263 3754 644272
rect 3608 643272 3660 643278
rect 3608 643214 3660 643220
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3424 314492 3476 314498
rect 3424 314434 3476 314440
rect 3528 314430 3556 632023
rect 3620 514865 3648 643214
rect 3712 566953 3740 644263
rect 3804 619177 3832 644438
rect 3790 619168 3846 619177
rect 3790 619103 3846 619112
rect 3698 566944 3754 566953
rect 3698 566879 3754 566888
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3882 358456 3938 358465
rect 3882 358391 3938 358400
rect 3606 319288 3662 319297
rect 3606 319223 3662 319232
rect 3620 318850 3648 319223
rect 3608 318844 3660 318850
rect 3608 318786 3660 318792
rect 3516 314424 3568 314430
rect 3516 314366 3568 314372
rect 3896 312934 3924 358391
rect 3884 312928 3936 312934
rect 3884 312870 3936 312876
rect 3332 312656 3384 312662
rect 3332 312598 3384 312604
rect 2964 306264 3016 306270
rect 2962 306232 2964 306241
rect 3016 306232 3018 306241
rect 2962 306167 3018 306176
rect 2780 293276 2832 293282
rect 2780 293218 2832 293224
rect 2792 293185 2820 293218
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2780 267232 2832 267238
rect 2778 267200 2780 267209
rect 2832 267200 2834 267209
rect 2778 267135 2834 267144
rect 3344 254153 3372 312598
rect 3976 312588 4028 312594
rect 3976 312530 4028 312536
rect 3700 312452 3752 312458
rect 3700 312394 3752 312400
rect 3608 311976 3660 311982
rect 3514 311944 3570 311953
rect 3608 311918 3660 311924
rect 3514 311879 3570 311888
rect 3424 309664 3476 309670
rect 3424 309606 3476 309612
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 2780 215008 2832 215014
rect 2778 214976 2780 214985
rect 2832 214976 2834 214985
rect 2778 214911 2834 214920
rect 2780 163396 2832 163402
rect 2780 163338 2832 163344
rect 2792 162897 2820 163338
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 2780 123888 2832 123894
rect 2780 123830 2832 123836
rect 2792 123729 2820 123830
rect 2778 123720 2834 123729
rect 2778 123655 2834 123664
rect 2780 110764 2832 110770
rect 2780 110706 2832 110712
rect 2792 110673 2820 110706
rect 2778 110664 2834 110673
rect 2778 110599 2834 110608
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 2780 85196 2832 85202
rect 2780 85138 2832 85144
rect 2792 84697 2820 85138
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 2780 71664 2832 71670
rect 2778 71632 2780 71641
rect 2832 71632 2834 71641
rect 2778 71567 2834 71576
rect 3148 45552 3200 45558
rect 3146 45520 3148 45529
rect 3200 45520 3202 45529
rect 3146 45455 3202 45464
rect 2780 32904 2832 32910
rect 2780 32846 2832 32852
rect 2792 32473 2820 32846
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 3436 6497 3464 309606
rect 3528 19417 3556 311879
rect 3620 58585 3648 311918
rect 3712 136785 3740 312394
rect 3792 312384 3844 312390
rect 3792 312326 3844 312332
rect 3804 149841 3832 312326
rect 3884 309868 3936 309874
rect 3884 309810 3936 309816
rect 3896 188873 3924 309810
rect 3988 201929 4016 312530
rect 4712 310072 4764 310078
rect 4712 310014 4764 310020
rect 4068 310004 4120 310010
rect 4068 309946 4120 309952
rect 4080 241097 4108 309946
rect 4724 293282 4752 310014
rect 4712 293276 4764 293282
rect 4712 293218 4764 293224
rect 4066 241088 4122 241097
rect 4066 241023 4122 241032
rect 3974 201920 4030 201929
rect 3974 201855 4030 201864
rect 3882 188864 3938 188873
rect 3882 188799 3938 188808
rect 3790 149832 3846 149841
rect 3790 149767 3846 149776
rect 3698 136776 3754 136785
rect 3698 136711 3754 136720
rect 4816 123894 4844 650014
rect 8220 314566 8248 702406
rect 24320 700942 24348 703520
rect 24308 700936 24360 700942
rect 24308 700878 24360 700884
rect 40512 700738 40540 703520
rect 40500 700732 40552 700738
rect 40500 700674 40552 700680
rect 72988 700398 73016 703520
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 89180 700330 89208 703520
rect 105464 700466 105492 703520
rect 105452 700460 105504 700466
rect 105452 700402 105504 700408
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 137848 700058 137876 703520
rect 147588 700528 147640 700534
rect 147588 700470 147640 700476
rect 147312 700460 147364 700466
rect 147312 700402 147364 700408
rect 147128 700392 147180 700398
rect 147128 700334 147180 700340
rect 147220 700392 147272 700398
rect 147220 700334 147272 700340
rect 146944 700324 146996 700330
rect 146944 700266 146996 700272
rect 147036 700324 147088 700330
rect 147036 700266 147088 700272
rect 137836 700052 137888 700058
rect 137836 699994 137888 700000
rect 40130 650176 40186 650185
rect 40130 650111 40186 650120
rect 40144 650078 40172 650111
rect 40132 650072 40184 650078
rect 40132 650014 40184 650020
rect 104714 645416 104770 645425
rect 104714 645351 104770 645360
rect 104728 644502 104756 645351
rect 104716 644496 104768 644502
rect 104716 644438 104768 644444
rect 98642 644328 98698 644337
rect 98642 644263 98644 644272
rect 98696 644263 98698 644272
rect 104254 644328 104310 644337
rect 104254 644263 104256 644272
rect 98644 644234 98696 644240
rect 104308 644263 104310 644272
rect 104256 644234 104308 644240
rect 133878 643648 133934 643657
rect 133800 643606 133878 643634
rect 133800 643278 133828 643606
rect 133878 643583 133934 643592
rect 133788 643272 133840 643278
rect 133788 643214 133840 643220
rect 40130 625696 40186 625705
rect 40130 625631 40186 625640
rect 40038 623520 40094 623529
rect 40038 623455 40094 623464
rect 40052 593366 40080 623455
rect 40040 593360 40092 593366
rect 40040 593302 40092 593308
rect 40038 582176 40094 582185
rect 40038 582111 40094 582120
rect 40052 437442 40080 582111
rect 40144 489870 40172 625631
rect 40222 606792 40278 606801
rect 40222 606727 40278 606736
rect 40236 540938 40264 606727
rect 114468 606416 114520 606422
rect 114468 606358 114520 606364
rect 118976 606416 119028 606422
rect 119988 606416 120040 606422
rect 119028 606364 119988 606370
rect 118976 606358 120040 606364
rect 114480 606121 114508 606358
rect 118988 606342 120028 606358
rect 114466 606112 114522 606121
rect 114466 606047 114522 606056
rect 118606 590744 118662 590753
rect 118606 590679 118662 590688
rect 92388 558952 92440 558958
rect 92388 558894 92440 558900
rect 40224 540932 40276 540938
rect 40224 540874 40276 540880
rect 40132 489864 40184 489870
rect 40132 489806 40184 489812
rect 40040 437436 40092 437442
rect 40040 437378 40092 437384
rect 89628 378208 89680 378214
rect 89628 378150 89680 378156
rect 88248 351960 88300 351966
rect 88248 351902 88300 351908
rect 82544 324352 82596 324358
rect 82544 324294 82596 324300
rect 8208 314560 8260 314566
rect 8208 314502 8260 314508
rect 77668 312996 77720 313002
rect 77668 312938 77720 312944
rect 6368 312860 6420 312866
rect 6368 312802 6420 312808
rect 5448 312792 5500 312798
rect 5448 312734 5500 312740
rect 5356 312724 5408 312730
rect 5356 312666 5408 312672
rect 5264 312520 5316 312526
rect 5264 312462 5316 312468
rect 5172 312316 5224 312322
rect 5172 312258 5224 312264
rect 5080 312248 5132 312254
rect 5080 312190 5132 312196
rect 4988 312112 5040 312118
rect 4988 312054 5040 312060
rect 4896 309732 4948 309738
rect 4896 309674 4948 309680
rect 4804 123888 4856 123894
rect 4804 123830 4856 123836
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 4908 32910 4936 309674
rect 5000 71670 5028 312054
rect 5092 85202 5120 312190
rect 5184 110770 5212 312258
rect 5276 163402 5304 312462
rect 5368 215014 5396 312666
rect 5460 267238 5488 312734
rect 6276 312180 6328 312186
rect 6276 312122 6328 312128
rect 6184 312044 6236 312050
rect 6184 311986 6236 311992
rect 5448 267232 5500 267238
rect 5448 267174 5500 267180
rect 5356 215008 5408 215014
rect 5356 214950 5408 214956
rect 5264 163396 5316 163402
rect 5264 163338 5316 163344
rect 5172 110764 5224 110770
rect 5172 110706 5224 110712
rect 5080 85196 5132 85202
rect 5080 85138 5132 85144
rect 4988 71664 5040 71670
rect 4988 71606 5040 71612
rect 6196 45558 6224 311986
rect 6288 97782 6316 312122
rect 6380 306270 6408 312802
rect 68006 312488 68062 312497
rect 68006 312423 68062 312432
rect 50986 312352 51042 312361
rect 50986 312287 51042 312296
rect 43994 312216 44050 312225
rect 43994 312151 44050 312160
rect 34334 312080 34390 312089
rect 34334 312015 34390 312024
rect 34348 310706 34376 312015
rect 44008 310706 44036 312151
rect 51000 310706 51028 312287
rect 68020 310706 68048 312423
rect 77680 310706 77708 312938
rect 82556 310706 82584 324294
rect 88260 313070 88288 351902
rect 87328 313064 87380 313070
rect 87328 313006 87380 313012
rect 88248 313064 88300 313070
rect 88248 313006 88300 313012
rect 84936 311908 84988 311914
rect 84936 311850 84988 311856
rect 84948 310706 84976 311850
rect 87340 310706 87368 313006
rect 89640 310706 89668 378150
rect 92400 316034 92428 558894
rect 99288 542428 99340 542434
rect 99288 542370 99340 542376
rect 96528 430636 96580 430642
rect 96528 430578 96580 430584
rect 95148 404388 95200 404394
rect 95148 404330 95200 404336
rect 92216 316006 92428 316034
rect 92216 310706 92244 316006
rect 95160 313070 95188 404330
rect 94504 313064 94556 313070
rect 94504 313006 94556 313012
rect 95148 313064 95200 313070
rect 95148 313006 95200 313012
rect 94516 310706 94544 313006
rect 34040 310678 34376 310706
rect 43700 310678 44036 310706
rect 50876 310678 51028 310706
rect 67712 310678 68048 310706
rect 77372 310678 77708 310706
rect 82156 310678 82584 310706
rect 84640 310678 84976 310706
rect 87032 310678 87368 310706
rect 89424 310678 89668 310706
rect 91816 310678 92244 310706
rect 94208 310678 94544 310706
rect 96540 310706 96568 430578
rect 99300 310706 99328 542370
rect 111708 536852 111760 536858
rect 111708 536794 111760 536800
rect 108948 510672 109000 510678
rect 108948 510614 109000 510620
rect 104808 484424 104860 484430
rect 104808 484366 104860 484372
rect 100760 457496 100812 457502
rect 100760 457438 100812 457444
rect 100772 325694 100800 457438
rect 100772 325666 101076 325694
rect 96540 310678 96600 310706
rect 99084 310678 99328 310706
rect 101048 310706 101076 325666
rect 104820 313070 104848 484366
rect 106188 470620 106240 470626
rect 106188 470562 106240 470568
rect 104164 313064 104216 313070
rect 104164 313006 104216 313012
rect 104808 313064 104860 313070
rect 104808 313006 104860 313012
rect 104176 310706 104204 313006
rect 101048 310678 101476 310706
rect 103868 310678 104204 310706
rect 106200 310706 106228 470562
rect 108960 310706 108988 510614
rect 111720 316034 111748 536794
rect 115848 533384 115900 533390
rect 115848 533326 115900 533332
rect 114468 524476 114520 524482
rect 114468 524418 114520 524424
rect 111444 316006 111748 316034
rect 111444 310706 111472 316006
rect 114480 313070 114508 524418
rect 113824 313064 113876 313070
rect 113824 313006 113876 313012
rect 114468 313064 114520 313070
rect 114468 313006 114520 313012
rect 113836 310706 113864 313006
rect 106200 310678 106260 310706
rect 108652 310678 108988 310706
rect 111044 310678 111472 310706
rect 113528 310678 113864 310706
rect 115860 310706 115888 533326
rect 118620 310706 118648 590679
rect 121366 576872 121422 576881
rect 121366 576807 121422 576816
rect 121380 316034 121408 576807
rect 143448 533452 143500 533458
rect 143448 533394 143500 533400
rect 121104 316006 121408 316034
rect 121104 310706 121132 316006
rect 135076 314356 135128 314362
rect 135076 314298 135128 314304
rect 133052 314220 133104 314226
rect 133052 314162 133104 314168
rect 130660 314152 130712 314158
rect 130660 314094 130712 314100
rect 128268 314084 128320 314090
rect 128268 314026 128320 314032
rect 125508 314016 125560 314022
rect 125508 313958 125560 313964
rect 123392 313948 123444 313954
rect 123392 313890 123444 313896
rect 123404 310706 123432 313890
rect 115860 310678 115920 310706
rect 118312 310678 118648 310706
rect 120704 310678 121132 310706
rect 123096 310678 123432 310706
rect 125520 310706 125548 313958
rect 128280 310706 128308 314026
rect 130672 310706 130700 314094
rect 133064 310706 133092 314162
rect 125520 310678 125580 310706
rect 127972 310678 128308 310706
rect 130364 310678 130700 310706
rect 132756 310678 133092 310706
rect 135088 310570 135116 314298
rect 137836 314288 137888 314294
rect 137836 314230 137888 314236
rect 137848 310706 137876 314230
rect 140320 313132 140372 313138
rect 140320 313074 140372 313080
rect 140332 310706 140360 313074
rect 143460 313070 143488 533394
rect 144736 313336 144788 313342
rect 144736 313278 144788 313284
rect 142712 313064 142764 313070
rect 142712 313006 142764 313012
rect 143448 313064 143500 313070
rect 143448 313006 143500 313012
rect 142724 310706 142752 313006
rect 137540 310678 137876 310706
rect 140024 310678 140360 310706
rect 142416 310678 142752 310706
rect 144748 310570 144776 313278
rect 146956 313206 146984 700266
rect 146944 313200 146996 313206
rect 146944 313142 146996 313148
rect 147048 313138 147076 700266
rect 147140 314634 147168 700334
rect 147128 314628 147180 314634
rect 147128 314570 147180 314576
rect 147232 313342 147260 700334
rect 147324 313886 147352 700402
rect 147312 313880 147364 313886
rect 147312 313822 147364 313828
rect 147220 313336 147272 313342
rect 147220 313278 147272 313284
rect 147036 313132 147088 313138
rect 147036 313074 147088 313080
rect 147600 310706 147628 700470
rect 150348 700460 150400 700466
rect 150348 700402 150400 700408
rect 150360 313070 150388 700402
rect 154132 699922 154160 703520
rect 166908 701004 166960 701010
rect 166908 700946 166960 700952
rect 162768 700868 162820 700874
rect 162768 700810 162820 700816
rect 154488 700664 154540 700670
rect 154488 700606 154540 700612
rect 154120 699916 154172 699922
rect 154120 699858 154172 699864
rect 153106 643920 153162 643929
rect 153106 643855 153162 643864
rect 153120 313138 153148 643855
rect 154500 625154 154528 700606
rect 157248 700596 157300 700602
rect 157248 700538 157300 700544
rect 154408 625126 154528 625154
rect 154408 615494 154436 625126
rect 154408 615466 154528 615494
rect 152280 313132 152332 313138
rect 152280 313074 152332 313080
rect 153108 313132 153160 313138
rect 153108 313074 153160 313080
rect 149888 313064 149940 313070
rect 149888 313006 149940 313012
rect 150348 313064 150400 313070
rect 150348 313006 150400 313012
rect 149900 310706 149928 313006
rect 152292 310706 152320 313074
rect 154500 310978 154528 615466
rect 147200 310678 147628 310706
rect 149592 310678 149928 310706
rect 151984 310678 152320 310706
rect 154454 310950 154528 310978
rect 154454 310692 154482 310950
rect 157260 310706 157288 700538
rect 160008 642932 160060 642938
rect 160008 642874 160060 642880
rect 160020 313138 160048 642874
rect 162780 313138 162808 700810
rect 164148 700800 164200 700806
rect 164148 700742 164200 700748
rect 159548 313132 159600 313138
rect 159548 313074 159600 313080
rect 160008 313132 160060 313138
rect 160008 313074 160060 313080
rect 161940 313132 161992 313138
rect 161940 313074 161992 313080
rect 162768 313132 162820 313138
rect 162768 313074 162820 313080
rect 159560 310706 159588 313074
rect 161952 310706 161980 313074
rect 164160 310706 164188 700742
rect 166920 310706 166948 700946
rect 169668 700188 169720 700194
rect 169668 700130 169720 700136
rect 167460 591320 167512 591326
rect 167460 591262 167512 591268
rect 167472 590753 167500 591262
rect 167458 590744 167514 590753
rect 167458 590679 167514 590688
rect 167458 580272 167514 580281
rect 167458 580207 167514 580216
rect 167472 579698 167500 580207
rect 167460 579692 167512 579698
rect 167460 579634 167512 579640
rect 167460 577516 167512 577522
rect 167460 577458 167512 577464
rect 167472 576881 167500 577458
rect 167458 576872 167514 576881
rect 167458 576807 167514 576816
rect 169680 313138 169708 700130
rect 170324 699786 170352 703520
rect 185124 700936 185176 700942
rect 185124 700878 185176 700884
rect 172428 700256 172480 700262
rect 172428 700198 172480 700204
rect 170312 699780 170364 699786
rect 170312 699722 170364 699728
rect 172440 313138 172468 700198
rect 173808 700120 173860 700126
rect 173808 700062 173860 700068
rect 169208 313132 169260 313138
rect 169208 313074 169260 313080
rect 169668 313132 169720 313138
rect 169668 313074 169720 313080
rect 171600 313132 171652 313138
rect 171600 313074 171652 313080
rect 172428 313132 172480 313138
rect 172428 313074 172480 313080
rect 169220 310706 169248 313074
rect 171612 310706 171640 313074
rect 173820 310706 173848 700062
rect 182180 700052 182232 700058
rect 182180 699994 182232 700000
rect 179328 699984 179380 699990
rect 179328 699926 179380 699932
rect 176568 699848 176620 699854
rect 176568 699790 176620 699796
rect 176580 316034 176608 699790
rect 176488 316006 176608 316034
rect 176488 310706 176516 316006
rect 179340 313138 179368 699926
rect 180064 699916 180116 699922
rect 180064 699858 180116 699864
rect 180076 313138 180104 699858
rect 180800 699780 180852 699786
rect 180800 699722 180852 699728
rect 178776 313132 178828 313138
rect 178776 313074 178828 313080
rect 179328 313132 179380 313138
rect 179328 313074 179380 313080
rect 180064 313132 180116 313138
rect 180064 313074 180116 313080
rect 178788 310706 178816 313074
rect 156860 310678 157288 310706
rect 159252 310678 159588 310706
rect 161644 310678 161980 310706
rect 164036 310678 164188 310706
rect 166520 310678 166948 310706
rect 168912 310678 169248 310706
rect 171304 310678 171640 310706
rect 173696 310678 173848 310706
rect 176088 310678 176516 310706
rect 178480 310678 178816 310706
rect 180812 310706 180840 699722
rect 182192 325694 182220 699994
rect 185136 643618 185164 700878
rect 202800 699854 202828 703520
rect 218992 699990 219020 703520
rect 235184 700126 235212 703520
rect 236000 700732 236052 700738
rect 236000 700674 236052 700680
rect 235172 700120 235224 700126
rect 235172 700062 235224 700068
rect 218980 699984 219032 699990
rect 218980 699926 219032 699932
rect 202788 699848 202840 699854
rect 202788 699790 202840 699796
rect 230480 683188 230532 683194
rect 230480 683130 230532 683136
rect 193128 670744 193180 670750
rect 193128 670686 193180 670692
rect 192390 645416 192446 645425
rect 192758 645416 192814 645425
rect 192446 645374 192758 645402
rect 192390 645351 192446 645360
rect 192758 645351 192814 645360
rect 193140 644722 193168 670686
rect 196992 650412 197044 650418
rect 196992 650354 197044 650360
rect 193140 644694 193214 644722
rect 192206 644328 192262 644337
rect 193186 644314 193214 644694
rect 196898 644328 196954 644337
rect 192206 644263 192262 644272
rect 193140 644286 193214 644314
rect 196544 644286 196898 644314
rect 189722 644056 189778 644065
rect 192220 644042 192248 644263
rect 192758 644056 192814 644065
rect 192220 644014 192758 644042
rect 189722 643991 189778 644000
rect 192758 643991 192814 644000
rect 189736 643793 189764 643991
rect 189722 643784 189778 643793
rect 189722 643719 189778 643728
rect 193140 643686 193168 644286
rect 196544 644065 196572 644286
rect 196898 644263 196954 644272
rect 196530 644056 196586 644065
rect 196530 643991 196586 644000
rect 193128 643680 193180 643686
rect 192206 643648 192262 643657
rect 185124 643612 185176 643618
rect 192758 643648 192814 643657
rect 192262 643606 192758 643634
rect 192206 643583 192262 643592
rect 193128 643622 193180 643628
rect 196622 643648 196678 643657
rect 192758 643583 192814 643592
rect 196622 643583 196624 643592
rect 185124 643554 185176 643560
rect 196676 643583 196678 643592
rect 196624 643554 196676 643560
rect 192206 643376 192262 643385
rect 185124 643340 185176 643346
rect 192206 643311 192262 643320
rect 185124 643282 185176 643288
rect 185136 640014 185164 643282
rect 192220 643142 192248 643311
rect 193128 643272 193180 643278
rect 193128 643214 193180 643220
rect 192208 643136 192260 643142
rect 192208 643078 192260 643084
rect 190918 642968 190974 642977
rect 190918 642903 190920 642912
rect 190972 642903 190974 642912
rect 190920 642874 190972 642880
rect 192208 642184 192260 642190
rect 192206 642152 192208 642161
rect 192260 642152 192262 642161
rect 192206 642087 192262 642096
rect 193140 640014 193168 643214
rect 197004 642870 197032 650354
rect 230492 646134 230520 683130
rect 236012 650622 236040 700674
rect 251468 699718 251496 703520
rect 267660 700194 267688 703520
rect 283852 700262 283880 703520
rect 300136 701010 300164 703520
rect 300124 701004 300176 701010
rect 300124 700946 300176 700952
rect 332520 700874 332548 703520
rect 332508 700868 332560 700874
rect 332508 700810 332560 700816
rect 348804 700806 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700800 348844 700806
rect 348792 700742 348844 700748
rect 283840 700256 283892 700262
rect 283840 700198 283892 700204
rect 267648 700188 267700 700194
rect 267648 700130 267700 700136
rect 251456 699712 251508 699718
rect 251456 699654 251508 699660
rect 252468 699712 252520 699718
rect 252468 699654 252520 699660
rect 252480 666534 252508 699654
rect 252468 666528 252520 666534
rect 252468 666470 252520 666476
rect 300768 666528 300820 666534
rect 300768 666470 300820 666476
rect 300780 665281 300808 666470
rect 300766 665272 300822 665281
rect 300766 665207 300822 665216
rect 236000 650616 236052 650622
rect 236000 650558 236052 650564
rect 230480 646128 230532 646134
rect 230480 646070 230532 646076
rect 230480 645516 230532 645522
rect 230480 645458 230532 645464
rect 202696 645448 202748 645454
rect 202694 645416 202696 645425
rect 202748 645416 202750 645425
rect 202694 645351 202750 645360
rect 201774 644872 201830 644881
rect 201774 644807 201830 644816
rect 199014 644328 199070 644337
rect 199290 644328 199346 644337
rect 199070 644286 199290 644314
rect 199014 644263 199070 644272
rect 199290 644263 199346 644272
rect 199384 643680 199436 643686
rect 198094 643648 198150 643657
rect 198016 643618 198094 643634
rect 198004 643612 198094 643618
rect 198056 643606 198094 643612
rect 198094 643583 198150 643592
rect 199290 643648 199346 643657
rect 199346 643628 199384 643634
rect 199346 643622 199436 643628
rect 199568 643680 199620 643686
rect 199658 643648 199714 643657
rect 199620 643628 199658 643634
rect 199568 643622 199658 643628
rect 199346 643606 199424 643622
rect 199580 643606 199658 643622
rect 199290 643583 199346 643592
rect 199658 643583 199714 643592
rect 198004 643554 198056 643560
rect 196992 642864 197044 642870
rect 196992 642806 197044 642812
rect 201788 642462 201816 644807
rect 204536 644292 204588 644298
rect 204536 644234 204588 644240
rect 202510 643784 202566 643793
rect 202786 643784 202842 643793
rect 202566 643742 202786 643770
rect 202510 643719 202566 643728
rect 202786 643719 202842 643728
rect 202234 643648 202290 643657
rect 204548 643618 204576 644234
rect 208398 643648 208454 643657
rect 202234 643583 202290 643592
rect 204536 643612 204588 643618
rect 202248 643249 202276 643583
rect 208398 643583 208454 643592
rect 204536 643554 204588 643560
rect 202234 643240 202290 643249
rect 202234 643175 202290 643184
rect 206558 643240 206614 643249
rect 208412 643210 208440 643583
rect 206558 643175 206614 643184
rect 208400 643204 208452 643210
rect 206572 643142 206600 643175
rect 208400 643146 208452 643152
rect 220176 643204 220228 643210
rect 220176 643146 220228 643152
rect 206560 643136 206612 643142
rect 206560 643078 206612 643084
rect 209688 643136 209740 643142
rect 209688 643078 209740 643084
rect 220084 643136 220136 643142
rect 220084 643078 220136 643084
rect 201776 642456 201828 642462
rect 201776 642398 201828 642404
rect 201776 642252 201828 642258
rect 201776 642194 201828 642200
rect 196900 640212 196952 640218
rect 196900 640154 196952 640160
rect 185124 640008 185176 640014
rect 185124 639950 185176 639956
rect 193128 640008 193180 640014
rect 193128 639950 193180 639956
rect 185124 639736 185176 639742
rect 185124 639678 185176 639684
rect 185136 636138 185164 639678
rect 193128 639600 193180 639606
rect 193128 639542 193180 639548
rect 193140 636206 193168 639542
rect 193128 636200 193180 636206
rect 193128 636142 193180 636148
rect 185124 636132 185176 636138
rect 185124 636074 185176 636080
rect 185124 635860 185176 635866
rect 185124 635802 185176 635808
rect 185136 632466 185164 635802
rect 193128 635792 193180 635798
rect 193128 635734 193180 635740
rect 193140 632534 193168 635734
rect 193128 632528 193180 632534
rect 193128 632470 193180 632476
rect 185124 632460 185176 632466
rect 185124 632402 185176 632408
rect 185124 632188 185176 632194
rect 185124 632130 185176 632136
rect 185136 628930 185164 632130
rect 193128 632120 193180 632126
rect 193128 632062 193180 632068
rect 193140 628998 193168 632062
rect 193128 628992 193180 628998
rect 193128 628934 193180 628940
rect 185124 628924 185176 628930
rect 185124 628866 185176 628872
rect 196912 628726 196940 640154
rect 196900 628720 196952 628726
rect 196900 628662 196952 628668
rect 185124 628652 185176 628658
rect 185124 628594 185176 628600
rect 182192 325666 182956 325694
rect 182928 310706 182956 325666
rect 185136 313274 185164 628594
rect 193128 628516 193180 628522
rect 193128 628458 193180 628464
rect 190460 314628 190512 314634
rect 190460 314570 190512 314576
rect 187792 313880 187844 313886
rect 187792 313822 187844 313828
rect 185124 313268 185176 313274
rect 185124 313210 185176 313216
rect 185676 313268 185728 313274
rect 185676 313210 185728 313216
rect 185688 313138 185716 313210
rect 185400 313132 185452 313138
rect 185400 313074 185452 313080
rect 185676 313132 185728 313138
rect 185676 313074 185728 313080
rect 185412 310706 185440 313074
rect 187804 310706 187832 313822
rect 190472 310706 190500 314570
rect 193140 313206 193168 628458
rect 196992 628380 197044 628386
rect 196992 628322 197044 628328
rect 197004 313342 197032 628322
rect 200764 462392 200816 462398
rect 200764 462334 200816 462340
rect 197452 314560 197504 314566
rect 197452 314502 197504 314508
rect 195704 313336 195756 313342
rect 195704 313278 195756 313284
rect 196992 313336 197044 313342
rect 196992 313278 197044 313284
rect 192576 313200 192628 313206
rect 192576 313142 192628 313148
rect 193128 313200 193180 313206
rect 193128 313142 193180 313148
rect 192588 310706 192616 313142
rect 195716 310706 195744 313278
rect 180812 310678 180964 310706
rect 182928 310678 183356 310706
rect 185412 310678 185748 310706
rect 187804 310678 188140 310706
rect 190472 310678 190532 310706
rect 192588 310678 192924 310706
rect 195408 310678 195744 310706
rect 197464 310706 197492 314502
rect 200120 313132 200172 313138
rect 200120 313074 200172 313080
rect 200132 310706 200160 313074
rect 200776 313070 200804 462334
rect 201788 313206 201816 642194
rect 209700 640492 209728 643078
rect 202236 639260 202288 639266
rect 202236 639202 202288 639208
rect 202248 634814 202276 639202
rect 201880 634786 202276 634814
rect 201880 325694 201908 634786
rect 220096 634710 220124 643078
rect 220188 640334 220216 643146
rect 220188 640306 220308 640334
rect 220280 634710 220308 640306
rect 230492 639985 230520 645458
rect 236182 644328 236238 644337
rect 236182 644263 236184 644272
rect 236236 644263 236238 644272
rect 240690 644328 240746 644337
rect 240690 644263 240692 644272
rect 236184 644234 236236 644240
rect 240744 644263 240746 644272
rect 240692 644234 240744 644240
rect 364352 642326 364380 702406
rect 381188 699718 381216 703520
rect 397472 700670 397500 703520
rect 397460 700664 397512 700670
rect 397460 700606 397512 700612
rect 413664 700602 413692 703520
rect 413652 700596 413704 700602
rect 413652 700538 413704 700544
rect 381176 699712 381228 699718
rect 381176 699654 381228 699660
rect 382188 699712 382240 699718
rect 382188 699654 382240 699660
rect 236184 642320 236236 642326
rect 236182 642288 236184 642297
rect 241612 642320 241664 642326
rect 236236 642288 236238 642297
rect 236182 642223 236238 642232
rect 241610 642288 241612 642297
rect 364340 642320 364392 642326
rect 241664 642288 241666 642297
rect 364340 642262 364392 642268
rect 241610 642223 241666 642232
rect 230478 639976 230534 639985
rect 230478 639911 230534 639920
rect 230478 639704 230534 639713
rect 230478 639639 230534 639648
rect 230492 639606 230520 639639
rect 224868 639600 224920 639606
rect 224866 639568 224868 639577
rect 230480 639600 230532 639606
rect 224920 639568 224922 639577
rect 230480 639542 230532 639548
rect 224866 639503 224922 639512
rect 220084 634704 220136 634710
rect 220084 634646 220136 634652
rect 220268 634704 220320 634710
rect 220268 634646 220320 634652
rect 219900 631984 219952 631990
rect 219900 631926 219952 631932
rect 220360 631984 220412 631990
rect 220360 631926 220412 631932
rect 219912 625154 219940 631926
rect 220372 625154 220400 631926
rect 219912 625126 220124 625154
rect 211160 606416 211212 606422
rect 211160 606358 211212 606364
rect 210424 579692 210476 579698
rect 210424 579634 210476 579640
rect 201880 325666 202184 325694
rect 201776 313200 201828 313206
rect 201776 313142 201828 313148
rect 200764 313064 200816 313070
rect 200764 313006 200816 313012
rect 202156 310706 202184 325666
rect 204628 314492 204680 314498
rect 204628 314434 204680 314440
rect 204640 310706 204668 314434
rect 209780 314424 209832 314430
rect 209780 314366 209832 314372
rect 207020 313132 207072 313138
rect 207020 313074 207072 313080
rect 207032 310706 207060 313074
rect 209792 310706 209820 314366
rect 210436 313138 210464 579634
rect 211172 325694 211200 606358
rect 218060 553444 218112 553450
rect 218060 553386 218112 553392
rect 217324 409896 217376 409902
rect 217324 409838 217376 409844
rect 211172 325666 211844 325694
rect 210424 313132 210476 313138
rect 210424 313074 210476 313080
rect 211816 310706 211844 325666
rect 214288 313200 214340 313206
rect 214288 313142 214340 313148
rect 214300 310706 214328 313142
rect 217336 313138 217364 409838
rect 218072 325694 218100 553386
rect 218072 325666 219020 325694
rect 216680 313132 216732 313138
rect 216680 313074 216732 313080
rect 217324 313132 217376 313138
rect 217324 313074 217376 313080
rect 216692 310706 216720 313074
rect 218992 310706 219020 325666
rect 220096 313410 220124 625126
rect 220188 625126 220400 625154
rect 220084 313404 220136 313410
rect 220084 313346 220136 313352
rect 220188 313342 220216 625126
rect 382200 615534 382228 699654
rect 429212 644366 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700534 462360 703520
rect 462320 700528 462372 700534
rect 462320 700470 462372 700476
rect 478524 700466 478552 703520
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 542372 702406 543504 702434
rect 558932 702406 559696 702434
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 443736 688696 443788 688702
rect 463332 688696 463384 688702
rect 443736 688638 443788 688644
rect 463330 688664 463332 688673
rect 463384 688664 463386 688673
rect 443748 654134 443776 688638
rect 463330 688599 463386 688608
rect 465538 688664 465594 688673
rect 465594 688622 465750 688650
rect 465538 688599 465594 688608
rect 542372 666466 542400 702406
rect 542360 666460 542412 666466
rect 542360 666402 542412 666408
rect 542360 661768 542412 661774
rect 542360 661710 542412 661716
rect 443748 654106 443868 654134
rect 443840 644842 443868 654106
rect 443828 644836 443880 644842
rect 443828 644778 443880 644784
rect 443736 644632 443788 644638
rect 443736 644574 443788 644580
rect 429200 644360 429252 644366
rect 429200 644302 429252 644308
rect 443748 639674 443776 644574
rect 471796 640892 471848 640898
rect 471796 640834 471848 640840
rect 471808 640529 471836 640834
rect 459558 640520 459614 640529
rect 459558 640455 459614 640464
rect 468666 640520 468722 640529
rect 469034 640520 469090 640529
rect 468722 640478 469034 640506
rect 468666 640455 468722 640464
rect 469034 640455 469090 640464
rect 471794 640520 471850 640529
rect 471794 640455 471850 640464
rect 459572 640354 459600 640455
rect 459560 640348 459612 640354
rect 459560 640290 459612 640296
rect 443736 639668 443788 639674
rect 443736 639610 443788 639616
rect 443644 639192 443696 639198
rect 443644 639134 443696 639140
rect 443736 639192 443788 639198
rect 443736 639134 443788 639140
rect 404266 628144 404322 628153
rect 404266 628079 404322 628088
rect 382188 615528 382240 615534
rect 382188 615470 382240 615476
rect 404280 566914 404308 628079
rect 424968 570648 425020 570654
rect 424968 570590 425020 570596
rect 424980 569974 425008 570590
rect 410340 569968 410392 569974
rect 410340 569910 410392 569916
rect 424324 569968 424376 569974
rect 424324 569910 424376 569916
rect 424968 569968 425020 569974
rect 424968 569910 425020 569916
rect 410352 567610 410380 569910
rect 410044 567582 410380 567610
rect 404268 566908 404320 566914
rect 404268 566850 404320 566856
rect 391846 559464 391902 559473
rect 391846 559399 391902 559408
rect 391860 558958 391888 559399
rect 391848 558952 391900 558958
rect 391848 558894 391900 558900
rect 391386 543552 391442 543561
rect 391386 543487 391442 543496
rect 391400 542434 391428 543487
rect 391388 542428 391440 542434
rect 391388 542370 391440 542376
rect 391756 542428 391808 542434
rect 391756 542370 391808 542376
rect 223580 527196 223632 527202
rect 223580 527138 223632 527144
rect 223592 325694 223620 527138
rect 226340 501016 226392 501022
rect 226340 500958 226392 500964
rect 223592 325666 223896 325694
rect 220176 313336 220228 313342
rect 220176 313278 220228 313284
rect 221556 313336 221608 313342
rect 221556 313278 221608 313284
rect 221568 310706 221596 313278
rect 223868 310706 223896 325666
rect 226352 310706 226380 500958
rect 230480 474768 230532 474774
rect 230480 474710 230532 474716
rect 230492 325694 230520 474710
rect 233240 448588 233292 448594
rect 233240 448530 233292 448536
rect 233252 325694 233280 448530
rect 237380 422340 237432 422346
rect 237380 422282 237432 422288
rect 237392 325694 237420 422282
rect 391768 419490 391796 542370
rect 391756 419484 391808 419490
rect 391756 419426 391808 419432
rect 240140 397520 240192 397526
rect 240140 397462 240192 397468
rect 240152 325694 240180 397462
rect 245660 371272 245712 371278
rect 245660 371214 245712 371220
rect 230492 325666 231072 325694
rect 233252 325666 233464 325694
rect 237392 325666 238340 325694
rect 240152 325666 240732 325694
rect 228732 313404 228784 313410
rect 228732 313346 228784 313352
rect 228744 310706 228772 313346
rect 231044 310706 231072 325666
rect 233436 310706 233464 325666
rect 236000 313064 236052 313070
rect 236000 313006 236052 313012
rect 236012 310706 236040 313006
rect 238312 310706 238340 325666
rect 240704 310706 240732 325666
rect 243176 313132 243228 313138
rect 243176 313074 243228 313080
rect 243188 310706 243216 313074
rect 245672 310706 245700 371214
rect 391860 365702 391888 558894
rect 402040 535758 402100 535786
rect 402072 534002 402100 535758
rect 417712 535622 418048 535650
rect 417712 534070 417740 535622
rect 417700 534064 417752 534070
rect 417700 534006 417752 534012
rect 401600 533996 401652 534002
rect 401600 533938 401652 533944
rect 402060 533996 402112 534002
rect 402060 533938 402112 533944
rect 401612 533458 401640 533938
rect 401600 533452 401652 533458
rect 401600 533394 401652 533400
rect 417712 533390 417740 534006
rect 417700 533384 417752 533390
rect 417700 533326 417752 533332
rect 424336 458182 424364 569910
rect 427820 566500 427872 566506
rect 427820 566442 427872 566448
rect 427832 551585 427860 566442
rect 427818 551576 427874 551585
rect 427818 551511 427874 551520
rect 424324 458176 424376 458182
rect 424324 458118 424376 458124
rect 424968 458176 425020 458182
rect 424968 458118 425020 458124
rect 424980 457502 425008 458118
rect 424968 457496 425020 457502
rect 424968 457438 425020 457444
rect 391848 365696 391900 365702
rect 391848 365638 391900 365644
rect 247040 345092 247092 345098
rect 247040 345034 247092 345040
rect 247052 325694 247080 345034
rect 247052 325666 247908 325694
rect 247880 310706 247908 325666
rect 252744 318844 252796 318850
rect 252744 318786 252796 318792
rect 250444 312928 250496 312934
rect 250444 312870 250496 312876
rect 250456 310706 250484 312870
rect 252756 310706 252784 318786
rect 443656 314362 443684 639134
rect 443748 570654 443776 639134
rect 542372 617914 542400 661710
rect 542360 617908 542412 617914
rect 542360 617850 542412 617856
rect 542360 613420 542412 613426
rect 542360 613362 542412 613368
rect 443736 570648 443788 570654
rect 443736 570590 443788 570596
rect 542372 534002 542400 613362
rect 542360 533996 542412 534002
rect 542360 533938 542412 533944
rect 443644 314356 443696 314362
rect 443644 314298 443696 314304
rect 558932 314294 558960 702406
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 580172 591320 580224 591326
rect 580172 591262 580224 591268
rect 580184 591025 580212 591262
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 577522 580212 577623
rect 580172 577516 580224 577522
rect 580172 577458 580224 577464
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 579618 484664 579674 484673
rect 579618 484599 579674 484608
rect 579632 484430 579660 484599
rect 579620 484424 579672 484430
rect 579620 484366 579672 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 579620 419484 579672 419490
rect 579620 419426 579672 419432
rect 579632 418305 579660 419426
rect 579618 418296 579674 418305
rect 579618 418231 579674 418240
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 579618 378448 579674 378457
rect 579618 378383 579674 378392
rect 579632 378214 579660 378383
rect 579620 378208 579672 378214
rect 579620 378150 579672 378156
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 580000 324358 580028 325207
rect 579988 324352 580040 324358
rect 579988 324294 580040 324300
rect 558920 314288 558972 314294
rect 558920 314230 558972 314236
rect 580276 314226 580304 697167
rect 580538 683904 580594 683913
rect 580538 683839 580594 683848
rect 580354 670712 580410 670721
rect 580354 670647 580410 670656
rect 580264 314220 580316 314226
rect 580264 314162 580316 314168
rect 580368 314158 580396 670647
rect 580446 644056 580502 644065
rect 580446 643991 580502 644000
rect 580356 314152 580408 314158
rect 580356 314094 580408 314100
rect 580460 314022 580488 643991
rect 580552 641714 580580 683839
rect 580540 641708 580592 641714
rect 580540 641650 580592 641656
rect 580538 630864 580594 630873
rect 580538 630799 580594 630808
rect 580552 314090 580580 630799
rect 580630 617536 580686 617545
rect 580630 617471 580686 617480
rect 580540 314084 580592 314090
rect 580540 314026 580592 314032
rect 580448 314016 580500 314022
rect 580448 313958 580500 313964
rect 580644 313954 580672 617471
rect 580722 564360 580778 564369
rect 580722 564295 580778 564304
rect 580736 534070 580764 564295
rect 580724 534064 580776 534070
rect 580724 534006 580776 534012
rect 580632 313948 580684 313954
rect 580632 313890 580684 313896
rect 304632 312996 304684 313002
rect 304632 312938 304684 312944
rect 257620 312860 257672 312866
rect 257620 312802 257672 312808
rect 257632 310706 257660 312802
rect 260012 312792 260064 312798
rect 260012 312734 260064 312740
rect 260024 310706 260052 312734
rect 267280 312724 267332 312730
rect 267280 312666 267332 312672
rect 264980 312656 265032 312662
rect 264980 312598 265032 312604
rect 264992 310706 265020 312598
rect 267292 310706 267320 312666
rect 272064 312588 272116 312594
rect 272064 312530 272116 312536
rect 272076 310706 272104 312530
rect 274640 312520 274692 312526
rect 274640 312462 274692 312468
rect 304446 312488 304502 312497
rect 274652 310706 274680 312462
rect 276940 312452 276992 312458
rect 304446 312423 304502 312432
rect 276940 312394 276992 312400
rect 276952 310706 276980 312394
rect 279332 312384 279384 312390
rect 279332 312326 279384 312332
rect 303342 312352 303398 312361
rect 279344 310706 279372 312326
rect 281724 312316 281776 312322
rect 303342 312287 303398 312296
rect 281724 312258 281776 312264
rect 281736 310706 281764 312258
rect 284300 312248 284352 312254
rect 284300 312190 284352 312196
rect 303158 312216 303214 312225
rect 284312 310706 284340 312190
rect 286508 312180 286560 312186
rect 303158 312151 303214 312160
rect 286508 312122 286560 312128
rect 286520 310706 286548 312122
rect 288900 312112 288952 312118
rect 288900 312054 288952 312060
rect 302882 312080 302938 312089
rect 288912 310706 288940 312054
rect 291384 312044 291436 312050
rect 302882 312015 302938 312024
rect 291384 311986 291436 311992
rect 291396 310706 291424 311986
rect 293960 311976 294012 311982
rect 293960 311918 294012 311924
rect 300950 311944 301006 311953
rect 293972 310706 294000 311918
rect 300950 311879 301006 311888
rect 300964 310706 300992 311879
rect 197464 310678 197800 310706
rect 200132 310678 200192 310706
rect 202156 310678 202584 310706
rect 204640 310678 204976 310706
rect 207032 310678 207368 310706
rect 209792 310678 209852 310706
rect 211816 310678 212244 310706
rect 214300 310678 214636 310706
rect 216692 310678 217028 310706
rect 218992 310678 219420 310706
rect 221568 310678 221904 310706
rect 223868 310678 224296 310706
rect 226352 310678 226688 310706
rect 228744 310678 229080 310706
rect 231044 310678 231472 310706
rect 233436 310678 233864 310706
rect 236012 310678 236348 310706
rect 238312 310678 238740 310706
rect 240704 310678 241132 310706
rect 243188 310678 243524 310706
rect 245672 310678 245916 310706
rect 247880 310678 248308 310706
rect 250456 310678 250792 310706
rect 252756 310678 253184 310706
rect 257632 310678 257968 310706
rect 260024 310678 260360 310706
rect 264992 310678 265236 310706
rect 267292 310678 267628 310706
rect 272076 310678 272412 310706
rect 274652 310678 274804 310706
rect 276952 310678 277288 310706
rect 279344 310678 279680 310706
rect 281736 310678 282072 310706
rect 284312 310678 284464 310706
rect 286520 310678 286856 310706
rect 288912 310678 289248 310706
rect 291396 310678 291732 310706
rect 293972 310678 294124 310706
rect 300964 310678 301300 310706
rect 135088 310542 135148 310570
rect 144748 310542 144808 310570
rect 79968 310480 80020 310486
rect 74980 310418 75316 310434
rect 79764 310428 79968 310434
rect 79764 310422 80020 310428
rect 74980 310412 75328 310418
rect 74980 310406 75276 310412
rect 79764 310406 80008 310422
rect 75276 310354 75328 310360
rect 70308 310344 70360 310350
rect 60536 310282 60688 310298
rect 62928 310282 63264 310298
rect 65320 310282 65656 310298
rect 70104 310292 70308 310298
rect 72884 310344 72936 310350
rect 70104 310286 70360 310292
rect 72588 310292 72884 310298
rect 72588 310286 72936 310292
rect 60536 310276 60700 310282
rect 60536 310270 60648 310276
rect 62928 310276 63276 310282
rect 62928 310270 63224 310276
rect 60648 310218 60700 310224
rect 65320 310276 65668 310282
rect 65320 310270 65616 310276
rect 63224 310218 63276 310224
rect 70104 310270 70348 310286
rect 72588 310270 72924 310286
rect 65616 310218 65668 310224
rect 55956 310208 56008 310214
rect 36432 310146 36768 310162
rect 38824 310146 39160 310162
rect 41216 310146 41368 310162
rect 46092 310146 46428 310162
rect 48484 310146 48820 310162
rect 53268 310146 53604 310162
rect 55660 310156 55956 310162
rect 58440 310208 58492 310214
rect 55660 310150 56008 310156
rect 58144 310156 58440 310162
rect 58144 310150 58492 310156
rect 36432 310140 36780 310146
rect 36432 310134 36728 310140
rect 38824 310140 39172 310146
rect 38824 310134 39120 310140
rect 36728 310082 36780 310088
rect 41216 310140 41380 310146
rect 41216 310134 41328 310140
rect 39120 310082 39172 310088
rect 46092 310140 46440 310146
rect 46092 310134 46388 310140
rect 41328 310082 41380 310088
rect 48484 310140 48832 310146
rect 48484 310134 48780 310140
rect 46388 310082 46440 310088
rect 53268 310140 53616 310146
rect 53268 310134 53564 310140
rect 48780 310082 48832 310088
rect 55660 310134 55996 310150
rect 58144 310134 58480 310150
rect 53564 310082 53616 310088
rect 255320 310072 255372 310078
rect 29550 310040 29606 310049
rect 29256 309998 29550 310026
rect 31758 310040 31814 310049
rect 31648 309998 31758 310026
rect 29550 309975 29606 309984
rect 255372 310020 255576 310026
rect 255320 310014 255576 310020
rect 255332 309998 255576 310014
rect 262508 310010 262844 310026
rect 269684 310010 270020 310026
rect 296180 310010 296516 310026
rect 298572 310010 298908 310026
rect 262496 310004 262844 310010
rect 31758 309975 31814 309984
rect 262548 309998 262844 310004
rect 269672 310004 270020 310010
rect 262496 309946 262548 309952
rect 269724 309998 270020 310004
rect 296168 310004 296516 310010
rect 269672 309946 269724 309952
rect 296220 309998 296516 310004
rect 298560 310004 298908 310010
rect 296168 309946 296220 309952
rect 298612 309998 298908 310004
rect 298560 309946 298612 309952
rect 6368 306264 6420 306270
rect 6368 306206 6420 306212
rect 6276 97776 6328 97782
rect 6276 97718 6328 97724
rect 6184 45552 6236 45558
rect 6184 45494 6236 45500
rect 27632 34054 28336 34082
rect 28552 34054 28888 34082
rect 29104 34054 29440 34082
rect 29656 34054 29992 34082
rect 30392 34054 30544 34082
rect 30760 34054 31096 34082
rect 31312 34054 31648 34082
rect 31864 34054 32200 34082
rect 32416 34054 32752 34082
rect 33152 34054 33304 34082
rect 33520 34054 33856 34082
rect 34072 34054 34408 34082
rect 34624 34054 34960 34082
rect 35176 34054 35512 34082
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 19248 31748 19300 31754
rect 19248 31690 19300 31696
rect 16488 31680 16540 31686
rect 16488 31622 16540 31628
rect 15108 31544 15160 31550
rect 15108 31486 15160 31492
rect 13728 31476 13780 31482
rect 13728 31418 13780 31424
rect 10968 31408 11020 31414
rect 10968 31350 11020 31356
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 6828 31204 6880 31210
rect 6828 31146 6880 31152
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 4068 31068 4120 31074
rect 4068 31010 4120 31016
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 2884 480 2912 3538
rect 4080 480 4108 31010
rect 5460 6914 5488 31078
rect 6840 6914 6868 31146
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7668 480 7696 3606
rect 9600 3398 9628 31214
rect 10980 3398 11008 31350
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 8772 480 8800 3334
rect 9968 480 9996 3334
rect 11164 480 11192 3334
rect 12268 1850 12296 3674
rect 12360 3398 12388 31282
rect 13740 6914 13768 31418
rect 15120 6914 15148 31486
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12268 1822 12388 1850
rect 12360 480 12388 1822
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3398 16528 31622
rect 17040 3868 17092 3874
rect 17040 3810 17092 3816
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 15948 480 15976 3334
rect 17052 480 17080 3810
rect 19260 3398 19288 31690
rect 20536 31612 20588 31618
rect 20536 31554 20588 31560
rect 20548 16574 20576 31554
rect 23388 31000 23440 31006
rect 23388 30942 23440 30948
rect 20628 30932 20680 30938
rect 20628 30874 20680 30880
rect 20456 16546 20576 16574
rect 19432 3800 19484 3806
rect 19432 3742 19484 3748
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 18248 480 18276 3334
rect 19444 480 19472 3742
rect 20456 3482 20484 16546
rect 20640 6914 20668 30874
rect 22008 30864 22060 30870
rect 22008 30806 22060 30812
rect 22020 6914 22048 30806
rect 23400 6914 23428 30942
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 20548 6886 20668 6914
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20548 3806 20576 6886
rect 20536 3800 20588 3806
rect 20536 3742 20588 3748
rect 20456 3454 20668 3482
rect 20640 480 20668 3454
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3398 24808 30738
rect 27528 30660 27580 30666
rect 27528 30602 27580 30608
rect 26148 30592 26200 30598
rect 26148 30534 26200 30540
rect 26160 3398 26188 30534
rect 27540 3534 27568 30602
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 24228 480 24256 3334
rect 25332 480 25360 3334
rect 26528 480 26556 3470
rect 27632 3466 27660 34054
rect 28552 26234 28580 34054
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 27816 26206 28580 26234
rect 27816 3670 27844 26206
rect 28828 16574 28856 30670
rect 28908 30524 28960 30530
rect 28908 30466 28960 30472
rect 28736 16546 28856 16574
rect 27804 3664 27856 3670
rect 27804 3606 27856 3612
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27620 3460 27672 3466
rect 27620 3402 27672 3408
rect 27724 480 27752 3538
rect 28736 3482 28764 16546
rect 28920 6914 28948 30466
rect 28828 6886 28948 6914
rect 28828 3602 28856 6886
rect 29104 4010 29132 34054
rect 29656 31074 29684 34054
rect 30392 31142 30420 34054
rect 30760 31210 30788 34054
rect 30748 31204 30800 31210
rect 30748 31146 30800 31152
rect 30380 31136 30432 31142
rect 30380 31078 30432 31084
rect 29644 31068 29696 31074
rect 29644 31010 29696 31016
rect 30288 31068 30340 31074
rect 30288 31010 30340 31016
rect 30300 6914 30328 31010
rect 31312 26234 31340 34054
rect 31864 31278 31892 34054
rect 32416 31414 32444 34054
rect 32404 31408 32456 31414
rect 32404 31350 32456 31356
rect 33152 31346 33180 34054
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 31852 31272 31904 31278
rect 31852 31214 31904 31220
rect 33048 31204 33100 31210
rect 33048 31146 33100 31152
rect 31668 31136 31720 31142
rect 31668 31078 31720 31084
rect 30116 6886 30328 6914
rect 30576 26206 31340 26234
rect 29092 4004 29144 4010
rect 29092 3946 29144 3952
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 28736 3454 28948 3482
rect 28920 480 28948 3454
rect 30116 480 30144 6886
rect 30576 3942 30604 26206
rect 31680 6914 31708 31078
rect 31312 6886 31708 6914
rect 30564 3936 30616 3942
rect 30564 3878 30616 3884
rect 31312 480 31340 6886
rect 33060 3534 33088 31146
rect 33520 26234 33548 34054
rect 34072 31482 34100 34054
rect 34624 31550 34652 34054
rect 35176 31686 35204 34054
rect 36050 33810 36078 34068
rect 36280 34054 36616 34082
rect 36832 34054 37168 34082
rect 37384 34054 37720 34082
rect 37936 34054 38272 34082
rect 38672 34054 38916 34082
rect 39132 34054 39468 34082
rect 39684 34054 40020 34082
rect 40236 34054 40572 34082
rect 40788 34054 41124 34082
rect 41432 34054 41676 34082
rect 41892 34054 42228 34082
rect 42444 34054 42780 34082
rect 42996 34054 43332 34082
rect 43548 34054 43884 34082
rect 44192 34054 44436 34082
rect 44652 34054 44988 34082
rect 45204 34054 45540 34082
rect 45756 34054 46092 34082
rect 46308 34054 46644 34082
rect 46952 34054 47196 34082
rect 47412 34054 47748 34082
rect 47964 34054 48300 34082
rect 48516 34054 48852 34082
rect 49160 34054 49496 34082
rect 49712 34054 50048 34082
rect 50264 34054 50600 34082
rect 51092 34054 51152 34082
rect 51276 34054 51704 34082
rect 51828 34054 52256 34082
rect 52564 34054 52808 34082
rect 53024 34054 53360 34082
rect 53912 34054 54064 34082
rect 54464 34054 54800 34082
rect 36050 33782 36124 33810
rect 35164 31680 35216 31686
rect 35164 31622 35216 31628
rect 34612 31544 34664 31550
rect 34612 31486 34664 31492
rect 34060 31476 34112 31482
rect 34060 31418 34112 31424
rect 34428 31340 34480 31346
rect 34428 31282 34480 31288
rect 33336 26206 33548 26234
rect 33336 3738 33364 26206
rect 33324 3732 33376 3738
rect 33324 3674 33376 3680
rect 34440 3534 34468 31282
rect 35808 31272 35860 31278
rect 35808 31214 35860 31220
rect 35820 3534 35848 31214
rect 36096 3806 36124 33782
rect 36280 31754 36308 34054
rect 36268 31748 36320 31754
rect 36268 31690 36320 31696
rect 36832 30938 36860 34054
rect 37384 31618 37412 34054
rect 37372 31612 37424 31618
rect 37372 31554 37424 31560
rect 36820 30932 36872 30938
rect 36820 30874 36872 30880
rect 37936 30870 37964 34054
rect 38568 31544 38620 31550
rect 38568 31486 38620 31492
rect 37924 30864 37976 30870
rect 37924 30806 37976 30812
rect 37096 30456 37148 30462
rect 37096 30398 37148 30404
rect 37108 16574 37136 30398
rect 37188 30388 37240 30394
rect 37188 30330 37240 30336
rect 37016 16546 37136 16574
rect 36084 3800 36136 3806
rect 36084 3742 36136 3748
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34808 480 34836 3470
rect 36004 480 36032 3538
rect 37016 3482 37044 16546
rect 37200 6914 37228 30330
rect 38580 6914 38608 31486
rect 38672 31006 38700 34054
rect 38660 31000 38712 31006
rect 38660 30942 38712 30948
rect 39132 30802 39160 34054
rect 39120 30796 39172 30802
rect 39120 30738 39172 30744
rect 39684 30598 39712 34054
rect 39948 31000 40000 31006
rect 39948 30942 40000 30948
rect 39672 30592 39724 30598
rect 39672 30534 39724 30540
rect 39960 6914 39988 30942
rect 40236 30666 40264 34054
rect 40224 30660 40276 30666
rect 40224 30602 40276 30608
rect 40788 30530 40816 34054
rect 41328 31748 41380 31754
rect 41328 31690 41380 31696
rect 40776 30524 40828 30530
rect 40776 30466 40828 30472
rect 37108 6886 37228 6914
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 37108 3602 37136 6886
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 37016 3454 37228 3482
rect 37200 480 37228 3454
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3534 41368 31690
rect 41432 30734 41460 34054
rect 41892 31074 41920 34054
rect 42444 31142 42472 34054
rect 42708 31612 42760 31618
rect 42708 31554 42760 31560
rect 42432 31136 42484 31142
rect 42432 31078 42484 31084
rect 41880 31068 41932 31074
rect 41880 31010 41932 31016
rect 41420 30728 41472 30734
rect 41420 30670 41472 30676
rect 42720 3534 42748 31554
rect 42996 31210 43024 34054
rect 43548 31346 43576 34054
rect 44088 31680 44140 31686
rect 44088 31622 44140 31628
rect 43536 31340 43588 31346
rect 43536 31282 43588 31288
rect 42984 31204 43036 31210
rect 42984 31146 43036 31152
rect 44100 3534 44128 31622
rect 44192 31278 44220 34054
rect 44180 31272 44232 31278
rect 44180 31214 44232 31220
rect 44652 30394 44680 34054
rect 45204 30462 45232 34054
rect 45756 31550 45784 34054
rect 45744 31544 45796 31550
rect 45744 31486 45796 31492
rect 45468 31340 45520 31346
rect 45468 31282 45520 31288
rect 45376 31204 45428 31210
rect 45376 31146 45428 31152
rect 45192 30456 45244 30462
rect 45192 30398 45244 30404
rect 44640 30388 44692 30394
rect 44640 30330 44692 30336
rect 45388 16574 45416 31146
rect 45296 16546 45416 16574
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3538
rect 45296 3482 45324 16546
rect 45480 6914 45508 31282
rect 46308 31006 46336 34054
rect 46952 31754 46980 34054
rect 46940 31748 46992 31754
rect 46940 31690 46992 31696
rect 47412 31618 47440 34054
rect 47964 31686 47992 34054
rect 47952 31680 48004 31686
rect 47952 31622 48004 31628
rect 47400 31612 47452 31618
rect 47400 31554 47452 31560
rect 48516 31346 48544 34054
rect 48504 31340 48556 31346
rect 48504 31282 48556 31288
rect 49160 31210 49188 34054
rect 49148 31204 49200 31210
rect 49148 31146 49200 31152
rect 46296 31000 46348 31006
rect 46296 30942 46348 30948
rect 49608 30524 49660 30530
rect 49608 30466 49660 30472
rect 46848 30456 46900 30462
rect 46848 30398 46900 30404
rect 46860 6914 46888 30398
rect 48228 30388 48280 30394
rect 48228 30330 48280 30336
rect 48240 6914 48268 30330
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 45388 3602 45416 6886
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45296 3454 45508 3482
rect 45480 480 45508 3454
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3534 49648 30466
rect 49712 30462 49740 34054
rect 49700 30456 49752 30462
rect 49700 30398 49752 30404
rect 50264 30394 50292 34054
rect 51092 30530 51120 34054
rect 51080 30524 51132 30530
rect 51080 30466 51132 30472
rect 51276 30410 51304 34054
rect 50252 30388 50304 30394
rect 50252 30330 50304 30336
rect 51000 30382 51304 30410
rect 51000 3534 51028 30382
rect 51828 26234 51856 34054
rect 52460 30388 52512 30394
rect 52460 30330 52512 30336
rect 51276 26206 51856 26234
rect 51276 16574 51304 26206
rect 51276 16546 51396 16574
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51368 480 51396 16546
rect 52472 3534 52500 30330
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 34054
rect 53024 30394 53052 34054
rect 53012 30388 53064 30394
rect 53012 30330 53064 30336
rect 54036 3534 54064 34054
rect 54772 30394 54800 34054
rect 55002 33810 55030 34068
rect 55568 34054 55904 34082
rect 56120 34054 56548 34082
rect 56672 34054 57008 34082
rect 57224 34054 57560 34082
rect 57776 34054 57928 34082
rect 58328 34054 58664 34082
rect 58880 34054 59308 34082
rect 59432 34054 59768 34082
rect 60076 34054 60504 34082
rect 55002 33782 55076 33810
rect 54760 30388 54812 30394
rect 54760 30330 54812 30336
rect 53748 3528 53800 3534
rect 53748 3470 53800 3476
rect 54024 3528 54076 3534
rect 54024 3470 54076 3476
rect 54944 3528 54996 3534
rect 54944 3470 54996 3476
rect 53760 480 53788 3470
rect 54956 480 54984 3470
rect 55048 3194 55076 33782
rect 55876 30394 55904 34054
rect 55128 30388 55180 30394
rect 55128 30330 55180 30336
rect 55864 30388 55916 30394
rect 55864 30330 55916 30336
rect 56416 30388 56468 30394
rect 56416 30330 56468 30336
rect 55140 3330 55168 30330
rect 56428 3534 56456 30330
rect 56416 3528 56468 3534
rect 56416 3470 56468 3476
rect 55128 3324 55180 3330
rect 55128 3266 55180 3272
rect 56048 3324 56100 3330
rect 56048 3266 56100 3272
rect 55036 3188 55088 3194
rect 55036 3130 55088 3136
rect 56060 480 56088 3266
rect 56520 3126 56548 34054
rect 56980 30394 57008 34054
rect 56968 30388 57020 30394
rect 56968 30330 57020 30336
rect 57532 26234 57560 34054
rect 57796 30388 57848 30394
rect 57796 30330 57848 30336
rect 57532 26206 57744 26234
rect 57716 3262 57744 26206
rect 57808 3466 57836 30330
rect 57796 3460 57848 3466
rect 57796 3402 57848 3408
rect 57900 3398 57928 34054
rect 58636 30394 58664 34054
rect 58624 30388 58676 30394
rect 58624 30330 58676 30336
rect 59176 30388 59228 30394
rect 59176 30330 59228 30336
rect 59188 3534 59216 30330
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59176 3528 59228 3534
rect 59176 3470 59228 3476
rect 57888 3392 57940 3398
rect 57888 3334 57940 3340
rect 57704 3256 57756 3262
rect 57704 3198 57756 3204
rect 57244 3188 57296 3194
rect 57244 3130 57296 3136
rect 56508 3120 56560 3126
rect 56508 3062 56560 3068
rect 57256 480 57284 3130
rect 58452 480 58480 3470
rect 59280 2922 59308 34054
rect 59740 30394 59768 34054
rect 59728 30388 59780 30394
rect 59728 30330 59780 30336
rect 60476 3670 60504 34054
rect 60568 34054 60628 34082
rect 61180 34054 61516 34082
rect 61732 34054 61976 34082
rect 62284 34054 62620 34082
rect 62836 34054 63172 34082
rect 60464 3664 60516 3670
rect 60464 3606 60516 3612
rect 60568 3602 60596 34054
rect 61488 30394 61516 34054
rect 60648 30388 60700 30394
rect 60648 30330 60700 30336
rect 61476 30388 61528 30394
rect 61476 30330 61528 30336
rect 60660 4010 60688 30330
rect 60648 4004 60700 4010
rect 60648 3946 60700 3952
rect 60556 3596 60608 3602
rect 60556 3538 60608 3544
rect 61948 3466 61976 34054
rect 62592 30394 62620 34054
rect 63144 30462 63172 34054
rect 63328 34054 63388 34082
rect 63940 34054 64276 34082
rect 64492 34054 64828 34082
rect 65044 34054 65380 34082
rect 65596 34054 65932 34082
rect 63132 30456 63184 30462
rect 63132 30398 63184 30404
rect 62028 30388 62080 30394
rect 62028 30330 62080 30336
rect 62580 30388 62632 30394
rect 62580 30330 62632 30336
rect 63224 30388 63276 30394
rect 63224 30330 63276 30336
rect 62040 3738 62068 30330
rect 63236 4026 63264 30330
rect 63328 4146 63356 34054
rect 63408 30456 63460 30462
rect 63408 30398 63460 30404
rect 63316 4140 63368 4146
rect 63316 4082 63368 4088
rect 63236 3998 63356 4026
rect 62028 3732 62080 3738
rect 62028 3674 62080 3680
rect 60832 3460 60884 3466
rect 60832 3402 60884 3408
rect 61936 3460 61988 3466
rect 61936 3402 61988 3408
rect 59636 3120 59688 3126
rect 59636 3062 59688 3068
rect 59268 2916 59320 2922
rect 59268 2858 59320 2864
rect 59648 480 59676 3062
rect 60844 480 60872 3402
rect 63224 3392 63276 3398
rect 63224 3334 63276 3340
rect 62028 3256 62080 3262
rect 62028 3198 62080 3204
rect 62040 480 62068 3198
rect 63236 480 63264 3334
rect 63328 3194 63356 3998
rect 63420 3262 63448 30398
rect 64248 30394 64276 34054
rect 64236 30388 64288 30394
rect 64236 30330 64288 30336
rect 64696 30388 64748 30394
rect 64696 30330 64748 30336
rect 64328 3528 64380 3534
rect 64328 3470 64380 3476
rect 63408 3256 63460 3262
rect 63408 3198 63460 3204
rect 63316 3188 63368 3194
rect 63316 3130 63368 3136
rect 64340 480 64368 3470
rect 64708 3398 64736 30330
rect 64800 3942 64828 34054
rect 65352 30394 65380 34054
rect 65904 30462 65932 34054
rect 66088 34054 66148 34082
rect 66700 34054 67036 34082
rect 67252 34054 67588 34082
rect 67804 34054 68140 34082
rect 68356 34054 68784 34082
rect 65892 30456 65944 30462
rect 65892 30398 65944 30404
rect 65340 30388 65392 30394
rect 65340 30330 65392 30336
rect 65984 30388 66036 30394
rect 65984 30330 66036 30336
rect 65996 4078 66024 30330
rect 65984 4072 66036 4078
rect 65984 4014 66036 4020
rect 64788 3936 64840 3942
rect 64788 3878 64840 3884
rect 64696 3392 64748 3398
rect 64696 3334 64748 3340
rect 66088 3330 66116 34054
rect 66168 30456 66220 30462
rect 66168 30398 66220 30404
rect 66180 3874 66208 30398
rect 67008 30394 67036 34054
rect 67560 31074 67588 34054
rect 67548 31068 67600 31074
rect 67548 31010 67600 31016
rect 68112 30394 68140 34054
rect 66996 30388 67048 30394
rect 66996 30330 67048 30336
rect 67548 30388 67600 30394
rect 67548 30330 67600 30336
rect 68100 30388 68152 30394
rect 68100 30330 68152 30336
rect 67560 4010 67588 30330
rect 68756 26234 68784 34054
rect 68848 34054 68908 34082
rect 69460 34054 69796 34082
rect 70012 34054 70256 34082
rect 70656 34054 70992 34082
rect 71208 34054 71544 34082
rect 68848 31686 68876 34054
rect 68836 31680 68888 31686
rect 68836 31622 68888 31628
rect 69768 30394 69796 34054
rect 68928 30388 68980 30394
rect 68928 30330 68980 30336
rect 69756 30388 69808 30394
rect 69756 30330 69808 30336
rect 68756 26206 68876 26234
rect 66720 4004 66772 4010
rect 66720 3946 66772 3952
rect 67548 4004 67600 4010
rect 67548 3946 67600 3952
rect 66168 3868 66220 3874
rect 66168 3810 66220 3816
rect 66076 3324 66128 3330
rect 66076 3266 66128 3272
rect 65524 2916 65576 2922
rect 65524 2858 65576 2864
rect 65536 480 65564 2858
rect 66732 480 66760 3946
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 67928 480 67956 3470
rect 68848 3126 68876 26206
rect 68940 3670 68968 30330
rect 70228 3806 70256 34054
rect 70964 31414 70992 34054
rect 70952 31408 71004 31414
rect 70952 31350 71004 31356
rect 71516 30394 71544 34054
rect 71608 34054 71760 34082
rect 72312 34054 72648 34082
rect 72864 34054 73108 34082
rect 73416 34054 73752 34082
rect 73968 34054 74304 34082
rect 70308 30388 70360 30394
rect 70308 30330 70360 30336
rect 71504 30388 71556 30394
rect 71504 30330 71556 30336
rect 70320 3890 70348 30330
rect 70320 3862 70440 3890
rect 70216 3800 70268 3806
rect 70216 3742 70268 3748
rect 70308 3732 70360 3738
rect 70308 3674 70360 3680
rect 68928 3664 68980 3670
rect 68928 3606 68980 3612
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 68836 3120 68888 3126
rect 68836 3062 68888 3068
rect 69124 480 69152 3538
rect 70320 480 70348 3674
rect 70412 3534 70440 3862
rect 71608 3602 71636 34054
rect 72620 31550 72648 34054
rect 72608 31544 72660 31550
rect 72608 31486 72660 31492
rect 71688 30388 71740 30394
rect 71688 30330 71740 30336
rect 71596 3596 71648 3602
rect 71596 3538 71648 3544
rect 70400 3528 70452 3534
rect 70400 3470 70452 3476
rect 71700 3466 71728 30330
rect 71504 3460 71556 3466
rect 71504 3402 71556 3408
rect 71688 3460 71740 3466
rect 71688 3402 71740 3408
rect 71516 480 71544 3402
rect 72608 3188 72660 3194
rect 72608 3130 72660 3136
rect 72620 480 72648 3130
rect 73080 2922 73108 34054
rect 73724 30394 73752 34054
rect 73712 30388 73764 30394
rect 73712 30330 73764 30336
rect 73804 3256 73856 3262
rect 73804 3198 73856 3204
rect 73068 2916 73120 2922
rect 73068 2858 73120 2864
rect 73816 480 73844 3198
rect 74276 2990 74304 34054
rect 74460 34054 74520 34082
rect 75072 34054 75500 34082
rect 75624 34054 75868 34082
rect 76176 34054 76512 34082
rect 76728 34054 77064 34082
rect 74356 30388 74408 30394
rect 74356 30330 74408 30336
rect 74264 2984 74316 2990
rect 74264 2926 74316 2932
rect 74368 2854 74396 30330
rect 74460 3058 74488 34054
rect 75472 26234 75500 34054
rect 75472 26206 75776 26234
rect 75000 4140 75052 4146
rect 75000 4082 75052 4088
rect 74448 3052 74500 3058
rect 74448 2994 74500 3000
rect 74356 2848 74408 2854
rect 74356 2790 74408 2796
rect 75012 480 75040 4082
rect 75748 3126 75776 26206
rect 75840 3194 75868 34054
rect 76484 30394 76512 34054
rect 77036 31278 77064 34054
rect 77220 34054 77280 34082
rect 77832 34054 78168 34082
rect 78384 34054 78628 34082
rect 78936 34054 79272 34082
rect 79488 34054 79824 34082
rect 77024 31272 77076 31278
rect 77024 31214 77076 31220
rect 76472 30388 76524 30394
rect 76472 30330 76524 30336
rect 77116 30388 77168 30394
rect 77116 30330 77168 30336
rect 76196 3392 76248 3398
rect 76196 3334 76248 3340
rect 75828 3188 75880 3194
rect 75828 3130 75880 3136
rect 75736 3120 75788 3126
rect 75736 3062 75788 3068
rect 76208 480 76236 3334
rect 77128 3262 77156 30330
rect 77220 4146 77248 34054
rect 78140 30394 78168 34054
rect 78600 31210 78628 34054
rect 78588 31204 78640 31210
rect 78588 31146 78640 31152
rect 79244 30394 79272 34054
rect 78128 30388 78180 30394
rect 78128 30330 78180 30336
rect 78588 30388 78640 30394
rect 78588 30330 78640 30336
rect 79232 30388 79284 30394
rect 79232 30330 79284 30336
rect 78600 6914 78628 30330
rect 78508 6886 78628 6914
rect 77208 4140 77260 4146
rect 77208 4082 77260 4088
rect 77392 3936 77444 3942
rect 77392 3878 77444 3884
rect 77116 3256 77168 3262
rect 77116 3198 77168 3204
rect 77404 480 77432 3878
rect 78508 3398 78536 6886
rect 78588 4072 78640 4078
rect 78588 4014 78640 4020
rect 78496 3392 78548 3398
rect 78496 3334 78548 3340
rect 78600 480 78628 4014
rect 79796 3942 79824 34054
rect 79980 34054 80040 34082
rect 80592 34054 80928 34082
rect 79876 30388 79928 30394
rect 79876 30330 79928 30336
rect 79888 4078 79916 30330
rect 79876 4072 79928 4078
rect 79876 4014 79928 4020
rect 79784 3936 79836 3942
rect 79784 3878 79836 3884
rect 79692 3868 79744 3874
rect 79692 3810 79744 3816
rect 79704 480 79732 3810
rect 79980 3641 80008 34054
rect 80900 30394 80928 34054
rect 81222 33810 81250 34068
rect 81788 34054 82124 34082
rect 82340 34054 82768 34082
rect 82892 34054 83228 34082
rect 83444 34054 83872 34082
rect 83996 34054 84148 34082
rect 84548 34054 84884 34082
rect 85100 34054 85436 34082
rect 85652 34054 85988 34082
rect 86204 34054 86540 34082
rect 86756 34054 86908 34082
rect 87308 34054 87644 34082
rect 87860 34054 88196 34082
rect 88412 34054 88748 34082
rect 88964 34054 89300 34082
rect 89516 34054 89668 34082
rect 90068 34054 90404 34082
rect 90620 34054 90956 34082
rect 91172 34054 91508 34082
rect 91816 34054 92244 34082
rect 81222 33782 81296 33810
rect 80888 30388 80940 30394
rect 80888 30330 80940 30336
rect 81268 3874 81296 33782
rect 82096 31142 82124 34054
rect 82084 31136 82136 31142
rect 82084 31078 82136 31084
rect 81348 30388 81400 30394
rect 81348 30330 81400 30336
rect 81360 4010 81388 30330
rect 81348 4004 81400 4010
rect 81348 3946 81400 3952
rect 81256 3868 81308 3874
rect 81256 3810 81308 3816
rect 82740 3806 82768 34054
rect 83200 31686 83228 34054
rect 83188 31680 83240 31686
rect 83188 31622 83240 31628
rect 83004 31068 83056 31074
rect 83004 31010 83056 31016
rect 83016 16574 83044 31010
rect 83844 26234 83872 34054
rect 83844 26206 84056 26234
rect 83016 16546 83320 16574
rect 80888 3800 80940 3806
rect 80888 3742 80940 3748
rect 82084 3800 82136 3806
rect 82084 3742 82136 3748
rect 82728 3800 82780 3806
rect 82728 3742 82780 3748
rect 79966 3632 80022 3641
rect 79966 3567 80022 3576
rect 80900 480 80928 3742
rect 82096 480 82124 3742
rect 83292 480 83320 16546
rect 84028 3505 84056 26206
rect 84014 3496 84070 3505
rect 84014 3431 84070 3440
rect 84120 3369 84148 34054
rect 84856 31346 84884 34054
rect 84844 31340 84896 31346
rect 84844 31282 84896 31288
rect 85408 31074 85436 34054
rect 85764 31612 85816 31618
rect 85764 31554 85816 31560
rect 85396 31068 85448 31074
rect 85396 31010 85448 31016
rect 85776 16574 85804 31554
rect 85960 30394 85988 34054
rect 86512 31482 86540 34054
rect 86500 31476 86552 31482
rect 86500 31418 86552 31424
rect 85948 30388 86000 30394
rect 85948 30330 86000 30336
rect 86776 30388 86828 30394
rect 86776 30330 86828 30336
rect 85776 16546 86448 16574
rect 84476 3664 84528 3670
rect 84476 3606 84528 3612
rect 84106 3360 84162 3369
rect 84106 3295 84162 3304
rect 84488 480 84516 3606
rect 85672 3528 85724 3534
rect 85672 3470 85724 3476
rect 85684 480 85712 3470
rect 86420 490 86448 16546
rect 86788 3534 86816 30330
rect 86880 3670 86908 34054
rect 87512 31544 87564 31550
rect 87512 31486 87564 31492
rect 87524 26234 87552 31486
rect 87616 30394 87644 34054
rect 88168 30666 88196 34054
rect 88156 30660 88208 30666
rect 88156 30602 88208 30608
rect 88720 30462 88748 34054
rect 88984 31408 89036 31414
rect 88984 31350 89036 31356
rect 88708 30456 88760 30462
rect 88708 30398 88760 30404
rect 87604 30388 87656 30394
rect 87604 30330 87656 30336
rect 88248 30388 88300 30394
rect 88248 30330 88300 30336
rect 87524 26206 87644 26234
rect 87616 3670 87644 26206
rect 88260 4622 88288 30330
rect 88248 4616 88300 4622
rect 88248 4558 88300 4564
rect 86868 3664 86920 3670
rect 86868 3606 86920 3612
rect 87604 3664 87656 3670
rect 87604 3606 87656 3612
rect 88996 3534 89024 31350
rect 89272 26234 89300 34054
rect 89640 30734 89668 34054
rect 90376 31686 90404 34054
rect 90272 31680 90324 31686
rect 90272 31622 90324 31628
rect 90364 31680 90416 31686
rect 90364 31622 90416 31628
rect 89628 30728 89680 30734
rect 89628 30670 89680 30676
rect 90284 26234 90312 31622
rect 90928 30870 90956 34054
rect 90916 30864 90968 30870
rect 90916 30806 90968 30812
rect 91480 30394 91508 34054
rect 92216 30546 92244 34054
rect 92308 34054 92368 34082
rect 92920 34054 93256 34082
rect 93472 34054 93716 34082
rect 94024 34054 94360 34082
rect 94576 34054 95004 34082
rect 92308 30938 92336 34054
rect 92296 30932 92348 30938
rect 92296 30874 92348 30880
rect 92216 30518 92428 30546
rect 91468 30388 91520 30394
rect 91468 30330 91520 30336
rect 92296 30388 92348 30394
rect 92296 30330 92348 30336
rect 89272 26206 89668 26234
rect 90284 26206 90404 26234
rect 89640 4690 89668 26206
rect 90376 16574 90404 26206
rect 90376 16546 90496 16574
rect 89628 4684 89680 4690
rect 89628 4626 89680 4632
rect 89168 3732 89220 3738
rect 89168 3674 89220 3680
rect 86776 3528 86828 3534
rect 86776 3470 86828 3476
rect 88984 3528 89036 3534
rect 88984 3470 89036 3476
rect 87972 3324 88024 3330
rect 87972 3266 88024 3272
rect 86696 598 86908 626
rect 86696 490 86724 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 462 86724 490
rect 86880 480 86908 598
rect 87984 480 88012 3266
rect 89180 480 89208 3674
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 90376 480 90404 3470
rect 90468 3330 90496 16546
rect 92308 4758 92336 30330
rect 92296 4752 92348 4758
rect 92296 4694 92348 4700
rect 92400 3466 92428 30518
rect 93124 30456 93176 30462
rect 93124 30398 93176 30404
rect 93136 3738 93164 30398
rect 93228 30394 93256 34054
rect 93688 31618 93716 34054
rect 93676 31612 93728 31618
rect 93676 31554 93728 31560
rect 94332 30394 94360 34054
rect 94504 31680 94556 31686
rect 94504 31622 94556 31628
rect 93216 30388 93268 30394
rect 93216 30330 93268 30336
rect 93768 30388 93820 30394
rect 93768 30330 93820 30336
rect 94320 30388 94372 30394
rect 94320 30330 94372 30336
rect 93780 5506 93808 30330
rect 93768 5500 93820 5506
rect 93768 5442 93820 5448
rect 93124 3732 93176 3738
rect 93124 3674 93176 3680
rect 94516 3602 94544 31622
rect 94872 30388 94924 30394
rect 94872 30330 94924 30336
rect 94884 26234 94912 30330
rect 94976 30138 95004 34054
rect 95114 33810 95142 34068
rect 95680 34054 96016 34082
rect 96232 34054 96568 34082
rect 96784 34054 97120 34082
rect 97336 34054 97672 34082
rect 95114 33782 95188 33810
rect 94976 30110 95096 30138
rect 94884 26206 95004 26234
rect 94976 5438 95004 26206
rect 94964 5432 95016 5438
rect 94964 5374 95016 5380
rect 95068 5370 95096 30110
rect 95056 5364 95108 5370
rect 95056 5306 95108 5312
rect 92756 3596 92808 3602
rect 92756 3538 92808 3544
rect 93952 3596 94004 3602
rect 93952 3538 94004 3544
rect 94504 3596 94556 3602
rect 94504 3538 94556 3544
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 92388 3460 92440 3466
rect 92388 3402 92440 3408
rect 90456 3324 90508 3330
rect 90456 3266 90508 3272
rect 91572 480 91600 3402
rect 92768 480 92796 3538
rect 93964 480 93992 3538
rect 95160 3074 95188 33782
rect 95884 31612 95936 31618
rect 95884 31554 95936 31560
rect 95160 3046 95280 3074
rect 95148 2916 95200 2922
rect 95148 2858 95200 2864
rect 95160 480 95188 2858
rect 95252 2786 95280 3046
rect 95896 2922 95924 31554
rect 95988 30394 96016 34054
rect 95976 30388 96028 30394
rect 95976 30330 96028 30336
rect 96436 30388 96488 30394
rect 96436 30330 96488 30336
rect 96448 5234 96476 30330
rect 96540 5302 96568 34054
rect 97092 30462 97120 34054
rect 97080 30456 97132 30462
rect 97080 30398 97132 30404
rect 97644 30394 97672 34054
rect 97736 34054 97888 34082
rect 98440 34054 98776 34082
rect 98992 34054 99236 34082
rect 99544 34054 99880 34082
rect 100096 34054 100340 34082
rect 97632 30388 97684 30394
rect 97632 30330 97684 30336
rect 96528 5296 96580 5302
rect 96528 5238 96580 5244
rect 96436 5228 96488 5234
rect 96436 5170 96488 5176
rect 97736 5098 97764 34054
rect 97908 30456 97960 30462
rect 97908 30398 97960 30404
rect 97816 30388 97868 30394
rect 97816 30330 97868 30336
rect 97828 5166 97856 30330
rect 97816 5160 97868 5166
rect 97816 5102 97868 5108
rect 97724 5092 97776 5098
rect 97724 5034 97776 5040
rect 97448 2984 97500 2990
rect 97448 2926 97500 2932
rect 95884 2916 95936 2922
rect 95884 2858 95936 2864
rect 96252 2848 96304 2854
rect 96252 2790 96304 2796
rect 95240 2780 95292 2786
rect 95240 2722 95292 2728
rect 96264 480 96292 2790
rect 97460 480 97488 2926
rect 97920 2854 97948 30398
rect 98748 30394 98776 34054
rect 98736 30388 98788 30394
rect 98736 30330 98788 30336
rect 99208 6322 99236 34054
rect 99852 30394 99880 34054
rect 100312 30462 100340 34054
rect 100496 34054 100648 34082
rect 101200 34054 101536 34082
rect 101752 34054 102088 34082
rect 102396 34054 102732 34082
rect 102948 34054 103376 34082
rect 100300 30456 100352 30462
rect 100300 30398 100352 30404
rect 99288 30388 99340 30394
rect 99288 30330 99340 30336
rect 99840 30388 99892 30394
rect 99840 30330 99892 30336
rect 99196 6316 99248 6322
rect 99196 6258 99248 6264
rect 98644 3052 98696 3058
rect 98644 2994 98696 3000
rect 97908 2848 97960 2854
rect 97908 2790 97960 2796
rect 98656 480 98684 2994
rect 99300 2990 99328 30330
rect 100496 6254 100524 34054
rect 101404 31476 101456 31482
rect 101404 31418 101456 31424
rect 100668 30456 100720 30462
rect 100668 30398 100720 30404
rect 100576 30388 100628 30394
rect 100576 30330 100628 30336
rect 100484 6248 100536 6254
rect 100484 6190 100536 6196
rect 100588 5030 100616 30330
rect 100576 5024 100628 5030
rect 100576 4966 100628 4972
rect 99840 3120 99892 3126
rect 99840 3062 99892 3068
rect 99288 2984 99340 2990
rect 99288 2926 99340 2932
rect 99852 480 99880 3062
rect 100680 3058 100708 30398
rect 101416 3194 101444 31418
rect 101508 30394 101536 34054
rect 102060 30802 102088 34054
rect 102324 31272 102376 31278
rect 102324 31214 102376 31220
rect 102048 30796 102100 30802
rect 102048 30738 102100 30744
rect 101496 30388 101548 30394
rect 101496 30330 101548 30336
rect 102048 30388 102100 30394
rect 102048 30330 102100 30336
rect 102060 4962 102088 30330
rect 102336 16574 102364 31214
rect 102704 30394 102732 34054
rect 102692 30388 102744 30394
rect 102692 30330 102744 30336
rect 103244 30388 103296 30394
rect 103244 30330 103296 30336
rect 102336 16546 103192 16574
rect 102048 4956 102100 4962
rect 102048 4898 102100 4904
rect 103164 3482 103192 16546
rect 103256 5574 103284 30330
rect 103244 5568 103296 5574
rect 103244 5510 103296 5516
rect 103348 4894 103376 34054
rect 103440 34054 103500 34082
rect 104052 34054 104388 34082
rect 104604 34054 104848 34082
rect 105156 34054 105492 34082
rect 105708 34054 106044 34082
rect 103336 4888 103388 4894
rect 103336 4830 103388 4836
rect 103164 3454 103376 3482
rect 102232 3256 102284 3262
rect 102232 3198 102284 3204
rect 101036 3188 101088 3194
rect 101036 3130 101088 3136
rect 101404 3188 101456 3194
rect 101404 3130 101456 3136
rect 100668 3052 100720 3058
rect 100668 2994 100720 3000
rect 101048 480 101076 3130
rect 102244 480 102272 3198
rect 103348 480 103376 3454
rect 103440 3074 103468 34054
rect 104360 31618 104388 34054
rect 104348 31612 104400 31618
rect 104348 31554 104400 31560
rect 104164 31204 104216 31210
rect 104164 31146 104216 31152
rect 104176 3398 104204 31146
rect 104820 5642 104848 34054
rect 105464 30394 105492 34054
rect 106016 31686 106044 34054
rect 106108 34054 106260 34082
rect 106812 34054 107148 34082
rect 106004 31680 106056 31686
rect 106004 31622 106056 31628
rect 105544 31408 105596 31414
rect 105544 31350 105596 31356
rect 105452 30388 105504 30394
rect 105452 30330 105504 30336
rect 105556 16574 105584 31350
rect 105556 16546 105860 16574
rect 104808 5636 104860 5642
rect 104808 5578 104860 5584
rect 104532 4140 104584 4146
rect 104532 4082 104584 4088
rect 104164 3392 104216 3398
rect 104164 3334 104216 3340
rect 103612 3188 103664 3194
rect 103612 3130 103664 3136
rect 103624 3074 103652 3130
rect 103440 3046 103652 3074
rect 104544 480 104572 4082
rect 105832 3262 105860 16546
rect 106108 5710 106136 34054
rect 107120 30394 107148 34054
rect 107350 33862 107378 34068
rect 107916 34054 108252 34082
rect 108468 34054 108896 34082
rect 109020 34054 109356 34082
rect 109572 34054 110000 34082
rect 110124 34054 110368 34082
rect 110676 34054 111012 34082
rect 111228 34054 111656 34082
rect 107338 33856 107390 33862
rect 107338 33798 107390 33804
rect 108224 30394 108252 34054
rect 108304 31136 108356 31142
rect 108304 31078 108356 31084
rect 106188 30388 106240 30394
rect 106188 30330 106240 30336
rect 107108 30388 107160 30394
rect 107108 30330 107160 30336
rect 107568 30388 107620 30394
rect 107568 30330 107620 30336
rect 108212 30388 108264 30394
rect 108212 30330 108264 30336
rect 106096 5704 106148 5710
rect 106096 5646 106148 5652
rect 106200 4826 106228 30330
rect 106188 4820 106240 4826
rect 106188 4762 106240 4768
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 105728 3256 105780 3262
rect 105728 3198 105780 3204
rect 105820 3256 105872 3262
rect 105820 3198 105872 3204
rect 105740 480 105768 3198
rect 106936 480 106964 3334
rect 107580 3262 107608 30330
rect 108316 16574 108344 31078
rect 108764 30388 108816 30394
rect 108764 30330 108816 30336
rect 108776 26234 108804 30330
rect 108868 30138 108896 34054
rect 109328 31414 109356 34054
rect 109972 31754 110000 34054
rect 109972 31726 110276 31754
rect 109316 31408 109368 31414
rect 109316 31350 109368 31356
rect 108868 30110 108988 30138
rect 108776 26206 108896 26234
rect 108316 16546 108436 16574
rect 108120 4072 108172 4078
rect 108120 4014 108172 4020
rect 107568 3256 107620 3262
rect 107568 3198 107620 3204
rect 108132 480 108160 4014
rect 108408 3806 108436 16546
rect 108868 5778 108896 26206
rect 108960 5846 108988 30110
rect 110248 5914 110276 31726
rect 110236 5908 110288 5914
rect 110236 5850 110288 5856
rect 108948 5840 109000 5846
rect 108948 5782 109000 5788
rect 108856 5772 108908 5778
rect 108856 5714 108908 5720
rect 110340 4214 110368 34054
rect 110984 31754 111012 34054
rect 110972 31748 111024 31754
rect 110972 31690 111024 31696
rect 111628 6186 111656 34054
rect 111720 34054 111780 34082
rect 112332 34054 112668 34082
rect 112976 34054 113128 34082
rect 113528 34054 113864 34082
rect 114080 34054 114416 34082
rect 114632 34054 114968 34082
rect 115184 34054 115612 34082
rect 115736 34054 115888 34082
rect 116288 34054 116624 34082
rect 116840 34054 117268 34082
rect 117392 34054 117728 34082
rect 117944 34054 118280 34082
rect 118496 34054 118648 34082
rect 119048 34054 119292 34082
rect 119600 34054 120028 34082
rect 120152 34054 120488 34082
rect 120704 34054 121040 34082
rect 111616 6180 111668 6186
rect 111616 6122 111668 6128
rect 110328 4208 110380 4214
rect 110328 4150 110380 4156
rect 111616 4140 111668 4146
rect 111616 4082 111668 4088
rect 109316 3936 109368 3942
rect 109316 3878 109368 3884
rect 108396 3800 108448 3806
rect 108396 3742 108448 3748
rect 109328 480 109356 3878
rect 110510 3632 110566 3641
rect 110510 3567 110566 3576
rect 110524 480 110552 3567
rect 111628 480 111656 4082
rect 111720 3398 111748 34054
rect 112640 31142 112668 34054
rect 112628 31136 112680 31142
rect 112628 31078 112680 31084
rect 113100 6050 113128 34054
rect 113836 30394 113864 34054
rect 114388 31210 114416 34054
rect 114376 31204 114428 31210
rect 114376 31146 114428 31152
rect 114940 30394 114968 34054
rect 115584 30546 115612 34054
rect 115860 31346 115888 34054
rect 115848 31340 115900 31346
rect 115848 31282 115900 31288
rect 115584 30518 115888 30546
rect 113824 30388 113876 30394
rect 113824 30330 113876 30336
rect 114468 30388 114520 30394
rect 114468 30330 114520 30336
rect 114928 30388 114980 30394
rect 114928 30330 114980 30336
rect 115756 30388 115808 30394
rect 115756 30330 115808 30336
rect 113088 6044 113140 6050
rect 113088 5986 113140 5992
rect 114480 5982 114508 30330
rect 115768 6118 115796 30330
rect 115756 6112 115808 6118
rect 115756 6054 115808 6060
rect 114468 5976 114520 5982
rect 114468 5918 114520 5924
rect 115860 4078 115888 30518
rect 116596 30394 116624 34054
rect 116584 30388 116636 30394
rect 116584 30330 116636 30336
rect 117136 30388 117188 30394
rect 117136 30330 117188 30336
rect 117148 6798 117176 30330
rect 117136 6792 117188 6798
rect 117136 6734 117188 6740
rect 115204 4072 115256 4078
rect 115204 4014 115256 4020
rect 115848 4072 115900 4078
rect 115848 4014 115900 4020
rect 114008 4004 114060 4010
rect 114008 3946 114060 3952
rect 112812 3868 112864 3874
rect 112812 3810 112864 3816
rect 111708 3392 111760 3398
rect 111708 3334 111760 3340
rect 112824 480 112852 3810
rect 114020 480 114048 3946
rect 115216 480 115244 4014
rect 117240 4010 117268 34054
rect 117700 30598 117728 34054
rect 118252 31754 118280 34054
rect 118252 31726 118556 31754
rect 117688 30592 117740 30598
rect 117688 30534 117740 30540
rect 118528 6730 118556 31726
rect 118516 6724 118568 6730
rect 118516 6666 118568 6672
rect 117964 4140 118016 4146
rect 117964 4082 118016 4088
rect 117976 4010 118004 4082
rect 117228 4004 117280 4010
rect 117228 3946 117280 3952
rect 117964 4004 118016 4010
rect 117964 3946 118016 3952
rect 118620 3874 118648 34054
rect 119264 31006 119292 34054
rect 119344 31068 119396 31074
rect 119344 31010 119396 31016
rect 119252 31000 119304 31006
rect 119252 30942 119304 30948
rect 118608 3868 118660 3874
rect 118608 3810 118660 3816
rect 119356 3534 119384 31010
rect 120000 6662 120028 34054
rect 120460 30394 120488 34054
rect 121012 31074 121040 34054
rect 121242 33810 121270 34068
rect 121808 34054 122144 34082
rect 122360 34054 122696 34082
rect 122912 34054 123248 34082
rect 123556 34054 123892 34082
rect 121242 33782 121316 33810
rect 121000 31068 121052 31074
rect 121000 31010 121052 31016
rect 120448 30388 120500 30394
rect 120448 30330 120500 30336
rect 119988 6656 120040 6662
rect 119988 6598 120040 6604
rect 121288 6594 121316 33782
rect 122116 30394 122144 34054
rect 121368 30388 121420 30394
rect 121368 30330 121420 30336
rect 122104 30388 122156 30394
rect 122104 30330 122156 30336
rect 121276 6588 121328 6594
rect 121276 6530 121328 6536
rect 121380 4078 121408 30330
rect 122668 4214 122696 34054
rect 123220 30394 123248 34054
rect 123864 30462 123892 34054
rect 124048 34054 124108 34082
rect 124660 34054 124996 34082
rect 125212 34054 125548 34082
rect 125764 34054 126100 34082
rect 126316 34054 126744 34082
rect 123852 30456 123904 30462
rect 123852 30398 123904 30404
rect 122748 30388 122800 30394
rect 122748 30330 122800 30336
rect 123208 30388 123260 30394
rect 123208 30330 123260 30336
rect 123944 30388 123996 30394
rect 123944 30330 123996 30336
rect 122656 4208 122708 4214
rect 122656 4150 122708 4156
rect 121368 4072 121420 4078
rect 121368 4014 121420 4020
rect 122760 3942 122788 30330
rect 123956 8226 123984 30330
rect 123944 8220 123996 8226
rect 123944 8162 123996 8168
rect 124048 4486 124076 34054
rect 124128 30456 124180 30462
rect 124128 30398 124180 30404
rect 124036 4480 124088 4486
rect 124036 4422 124088 4428
rect 124140 4010 124168 30398
rect 124968 30394 124996 34054
rect 124956 30388 125008 30394
rect 124956 30330 125008 30336
rect 125416 30388 125468 30394
rect 125416 30330 125468 30336
rect 125428 8158 125456 30330
rect 125416 8152 125468 8158
rect 125416 8094 125468 8100
rect 123484 4004 123536 4010
rect 123484 3946 123536 3952
rect 124128 4004 124180 4010
rect 124128 3946 124180 3952
rect 119896 3936 119948 3942
rect 119896 3878 119948 3884
rect 122748 3936 122800 3942
rect 122748 3878 122800 3884
rect 119344 3528 119396 3534
rect 117594 3496 117650 3505
rect 119344 3470 119396 3476
rect 117594 3431 117650 3440
rect 116400 3324 116452 3330
rect 116400 3266 116452 3272
rect 116412 480 116440 3266
rect 117608 480 117636 3431
rect 118790 3360 118846 3369
rect 118790 3295 118846 3304
rect 118804 480 118832 3295
rect 119908 480 119936 3878
rect 122288 3664 122340 3670
rect 122288 3606 122340 3612
rect 121092 3528 121144 3534
rect 121092 3470 121144 3476
rect 121104 480 121132 3470
rect 122300 480 122328 3606
rect 123496 480 123524 3946
rect 125520 3806 125548 34054
rect 126072 30394 126100 34054
rect 126060 30388 126112 30394
rect 126060 30330 126112 30336
rect 126716 8090 126744 34054
rect 126854 33810 126882 34068
rect 127420 34054 127756 34082
rect 127972 34054 128308 34082
rect 128524 34054 128860 34082
rect 129076 34054 129412 34082
rect 126854 33782 126928 33810
rect 126796 30388 126848 30394
rect 126796 30330 126848 30336
rect 126704 8084 126756 8090
rect 126704 8026 126756 8032
rect 125876 4616 125928 4622
rect 125876 4558 125928 4564
rect 124680 3800 124732 3806
rect 124680 3742 124732 3748
rect 125508 3800 125560 3806
rect 125508 3742 125560 3748
rect 124692 480 124720 3742
rect 125888 480 125916 4558
rect 126808 4350 126836 30330
rect 126796 4344 126848 4350
rect 126796 4286 126848 4292
rect 126900 3670 126928 33782
rect 127164 30660 127216 30666
rect 127164 30602 127216 30608
rect 127176 6914 127204 30602
rect 127728 30394 127756 34054
rect 128280 30598 128308 34054
rect 128268 30592 128320 30598
rect 128268 30534 128320 30540
rect 128832 30462 128860 34054
rect 128820 30456 128872 30462
rect 128820 30398 128872 30404
rect 129384 30394 129412 34054
rect 129476 34054 129628 34082
rect 130180 34054 130516 34082
rect 130732 34054 130976 34082
rect 131284 34054 131620 34082
rect 131836 34054 132172 34082
rect 127716 30388 127768 30394
rect 127716 30330 127768 30336
rect 128268 30388 128320 30394
rect 128268 30330 128320 30336
rect 129372 30388 129424 30394
rect 129372 30330 129424 30336
rect 126992 6886 127204 6914
rect 126888 3664 126940 3670
rect 126888 3606 126940 3612
rect 126992 480 127020 6886
rect 128280 4418 128308 30330
rect 129476 7954 129504 34054
rect 129740 30728 129792 30734
rect 129740 30670 129792 30676
rect 129648 30456 129700 30462
rect 129648 30398 129700 30404
rect 129556 30388 129608 30394
rect 129556 30330 129608 30336
rect 129464 7948 129516 7954
rect 129464 7890 129516 7896
rect 129372 4684 129424 4690
rect 129372 4626 129424 4632
rect 128268 4412 128320 4418
rect 128268 4354 128320 4360
rect 127440 4004 127492 4010
rect 127440 3946 127492 3952
rect 127452 3890 127480 3946
rect 127452 3862 127848 3890
rect 127820 3806 127848 3862
rect 127808 3800 127860 3806
rect 127808 3742 127860 3748
rect 128176 3732 128228 3738
rect 128176 3674 128228 3680
rect 128188 480 128216 3674
rect 129384 480 129412 4626
rect 129568 4282 129596 30330
rect 129556 4276 129608 4282
rect 129556 4218 129608 4224
rect 129660 3670 129688 30398
rect 129752 16574 129780 30670
rect 130488 30394 130516 34054
rect 130476 30388 130528 30394
rect 130476 30330 130528 30336
rect 129752 16546 130608 16574
rect 129648 3664 129700 3670
rect 129648 3606 129700 3612
rect 130580 480 130608 16546
rect 130948 4554 130976 34054
rect 131592 30394 131620 34054
rect 132144 30462 132172 34054
rect 132328 34054 132388 34082
rect 132940 34054 133276 34082
rect 133492 34054 133828 34082
rect 134136 34054 134472 34082
rect 134688 34054 135024 34082
rect 132132 30456 132184 30462
rect 132132 30398 132184 30404
rect 131028 30388 131080 30394
rect 131028 30330 131080 30336
rect 131580 30388 131632 30394
rect 131580 30330 131632 30336
rect 132224 30388 132276 30394
rect 132224 30330 132276 30336
rect 130936 4548 130988 4554
rect 130936 4490 130988 4496
rect 131040 3777 131068 30330
rect 132236 8022 132264 30330
rect 132224 8016 132276 8022
rect 132224 7958 132276 7964
rect 132328 4622 132356 34054
rect 132500 30660 132552 30666
rect 132500 30602 132552 30608
rect 132408 30456 132460 30462
rect 132408 30398 132460 30404
rect 132316 4616 132368 4622
rect 132316 4558 132368 4564
rect 131026 3768 131082 3777
rect 131026 3703 131082 3712
rect 131764 3596 131816 3602
rect 131764 3538 131816 3544
rect 131776 480 131804 3538
rect 132420 3534 132448 30398
rect 132512 16574 132540 30602
rect 133248 30394 133276 34054
rect 133236 30388 133288 30394
rect 133236 30330 133288 30336
rect 133696 30388 133748 30394
rect 133696 30330 133748 30336
rect 132512 16546 133000 16574
rect 132408 3528 132460 3534
rect 132408 3470 132460 3476
rect 132972 480 133000 16546
rect 133708 7886 133736 30330
rect 133696 7880 133748 7886
rect 133696 7822 133748 7828
rect 133800 3641 133828 34054
rect 134444 30394 134472 34054
rect 134432 30388 134484 30394
rect 134432 30330 134484 30336
rect 134996 7818 135024 34054
rect 135180 34054 135240 34082
rect 135792 34054 136128 34082
rect 136344 34054 136588 34082
rect 136896 34054 137232 34082
rect 137448 34054 137876 34082
rect 135076 30388 135128 30394
rect 135076 30330 135128 30336
rect 134984 7812 135036 7818
rect 134984 7754 135036 7760
rect 134156 4752 134208 4758
rect 134156 4694 134208 4700
rect 133786 3632 133842 3641
rect 133786 3567 133842 3576
rect 134168 480 134196 4694
rect 135088 4690 135116 30330
rect 135076 4684 135128 4690
rect 135076 4626 135128 4632
rect 135180 3505 135208 34054
rect 135444 30932 135496 30938
rect 135444 30874 135496 30880
rect 135456 16574 135484 30874
rect 136100 30394 136128 34054
rect 136560 30666 136588 34054
rect 136548 30660 136600 30666
rect 136548 30602 136600 30608
rect 137204 30394 137232 34054
rect 136088 30388 136140 30394
rect 136088 30330 136140 30336
rect 136548 30388 136600 30394
rect 136548 30330 136600 30336
rect 137192 30388 137244 30394
rect 137192 30330 137244 30336
rect 135456 16546 136496 16574
rect 135166 3496 135222 3505
rect 135166 3431 135222 3440
rect 135260 3460 135312 3466
rect 135260 3402 135312 3408
rect 135272 480 135300 3402
rect 136468 480 136496 16546
rect 136560 4758 136588 30330
rect 137848 5506 137876 34054
rect 137940 34054 138000 34082
rect 138552 34054 138980 34082
rect 139104 34054 139348 34082
rect 139656 34054 139992 34082
rect 140208 34054 140544 34082
rect 137940 30666 137968 34054
rect 137928 30660 137980 30666
rect 137928 30602 137980 30608
rect 137928 30388 137980 30394
rect 137928 30330 137980 30336
rect 137652 5500 137704 5506
rect 137652 5442 137704 5448
rect 137836 5500 137888 5506
rect 137836 5442 137888 5448
rect 136548 4752 136600 4758
rect 136548 4694 136600 4700
rect 137664 480 137692 5442
rect 137940 3466 137968 30330
rect 138952 26234 138980 34054
rect 138952 26206 139256 26234
rect 139228 7750 139256 26206
rect 139216 7744 139268 7750
rect 139216 7686 139268 7692
rect 139320 5137 139348 34054
rect 139964 30870 139992 34054
rect 139952 30864 140004 30870
rect 139952 30806 140004 30812
rect 140516 30394 140544 34054
rect 140608 34054 140760 34082
rect 141312 34054 141648 34082
rect 141864 34054 142016 34082
rect 142416 34054 142752 34082
rect 142968 34054 143396 34082
rect 140504 30388 140556 30394
rect 140504 30330 140556 30336
rect 140608 5438 140636 34054
rect 141620 30394 141648 34054
rect 140688 30388 140740 30394
rect 140688 30330 140740 30336
rect 141608 30388 141660 30394
rect 141608 30330 141660 30336
rect 140044 5432 140096 5438
rect 140044 5374 140096 5380
rect 140596 5432 140648 5438
rect 140596 5374 140648 5380
rect 139306 5128 139362 5137
rect 139306 5063 139362 5072
rect 137928 3460 137980 3466
rect 137928 3402 137980 3408
rect 138848 2848 138900 2854
rect 138848 2790 138900 2796
rect 138860 480 138888 2790
rect 140056 480 140084 5374
rect 140700 3369 140728 30330
rect 141988 7682 142016 34054
rect 142724 30394 142752 34054
rect 142804 30728 142856 30734
rect 142804 30670 142856 30676
rect 142068 30388 142120 30394
rect 142068 30330 142120 30336
rect 142712 30388 142764 30394
rect 142712 30330 142764 30336
rect 141976 7676 142028 7682
rect 141976 7618 142028 7624
rect 142080 6866 142108 30330
rect 142068 6860 142120 6866
rect 142068 6802 142120 6808
rect 141240 5364 141292 5370
rect 141240 5306 141292 5312
rect 140686 3360 140742 3369
rect 140686 3295 140742 3304
rect 141252 480 141280 5306
rect 142816 2922 142844 30670
rect 143264 30388 143316 30394
rect 143264 30330 143316 30336
rect 143276 7614 143304 30330
rect 143264 7608 143316 7614
rect 143264 7550 143316 7556
rect 143368 6526 143396 34054
rect 143460 34054 143520 34082
rect 144072 34054 144408 34082
rect 143460 30394 143488 34054
rect 144380 30394 144408 34054
rect 144702 33810 144730 34068
rect 145268 34054 145604 34082
rect 145820 34054 146248 34082
rect 146372 34054 146708 34082
rect 146924 34054 147352 34082
rect 147476 34054 147628 34082
rect 148028 34054 148364 34082
rect 148580 34054 148916 34082
rect 149132 34054 149468 34082
rect 149684 34054 150020 34082
rect 144702 33782 144776 33810
rect 143448 30388 143500 30394
rect 143448 30330 143500 30336
rect 144368 30388 144420 30394
rect 144368 30330 144420 30336
rect 143448 30252 143500 30258
rect 143448 30194 143500 30200
rect 143356 6520 143408 6526
rect 143356 6462 143408 6468
rect 143460 5370 143488 30194
rect 144748 6458 144776 33782
rect 145576 30394 145604 34054
rect 144828 30388 144880 30394
rect 144828 30330 144880 30336
rect 145564 30388 145616 30394
rect 145564 30330 145616 30336
rect 146116 30388 146168 30394
rect 146116 30330 146168 30336
rect 144736 6452 144788 6458
rect 144736 6394 144788 6400
rect 143448 5364 143500 5370
rect 143448 5306 143500 5312
rect 144840 5302 144868 30330
rect 146128 8498 146156 30330
rect 146116 8492 146168 8498
rect 146116 8434 146168 8440
rect 144736 5296 144788 5302
rect 144736 5238 144788 5244
rect 144828 5296 144880 5302
rect 144828 5238 144880 5244
rect 143540 5228 143592 5234
rect 143540 5170 143592 5176
rect 142436 2916 142488 2922
rect 142436 2858 142488 2864
rect 142804 2916 142856 2922
rect 142804 2858 142856 2864
rect 142448 480 142476 2858
rect 143552 480 143580 5170
rect 144748 480 144776 5238
rect 146220 5234 146248 34054
rect 146680 30394 146708 34054
rect 146668 30388 146720 30394
rect 146668 30330 146720 30336
rect 147324 26234 147352 34054
rect 147496 30388 147548 30394
rect 147496 30330 147548 30336
rect 147324 26206 147444 26234
rect 147416 8566 147444 26206
rect 147404 8560 147456 8566
rect 147404 8502 147456 8508
rect 147508 6390 147536 30330
rect 147496 6384 147548 6390
rect 147496 6326 147548 6332
rect 146208 5228 146260 5234
rect 146208 5170 146260 5176
rect 147600 5166 147628 34054
rect 148336 30394 148364 34054
rect 148324 30388 148376 30394
rect 148324 30330 148376 30336
rect 148888 8634 148916 34054
rect 149440 30462 149468 34054
rect 149428 30456 149480 30462
rect 149428 30398 149480 30404
rect 149992 30394 150020 34054
rect 150176 34054 150236 34082
rect 150788 34054 151124 34082
rect 151340 34054 151676 34082
rect 151892 34054 152228 34082
rect 152444 34054 152780 34082
rect 148968 30388 149020 30394
rect 148968 30330 149020 30336
rect 149980 30388 150032 30394
rect 149980 30330 150032 30336
rect 148876 8628 148928 8634
rect 148876 8570 148928 8576
rect 148980 6633 149008 30330
rect 150176 8770 150204 34054
rect 150348 30456 150400 30462
rect 150348 30398 150400 30404
rect 150256 30388 150308 30394
rect 150256 30330 150308 30336
rect 150164 8764 150216 8770
rect 150164 8706 150216 8712
rect 148966 6624 149022 6633
rect 148966 6559 149022 6568
rect 150268 6497 150296 30330
rect 150254 6488 150310 6497
rect 150254 6423 150310 6432
rect 147128 5160 147180 5166
rect 147128 5102 147180 5108
rect 147588 5160 147640 5166
rect 147588 5102 147640 5108
rect 145932 2984 145984 2990
rect 145932 2926 145984 2932
rect 145944 480 145972 2926
rect 147140 480 147168 5102
rect 150360 5098 150388 30398
rect 151096 30394 151124 34054
rect 151084 30388 151136 30394
rect 151084 30330 151136 30336
rect 151648 6322 151676 34054
rect 152200 30394 152228 34054
rect 152752 30462 152780 34054
rect 152982 33810 153010 34068
rect 153548 34054 153884 34082
rect 154100 34054 154528 34082
rect 154652 34054 154988 34082
rect 155296 34054 155724 34082
rect 152982 33782 153056 33810
rect 152740 30456 152792 30462
rect 152740 30398 152792 30404
rect 151728 30388 151780 30394
rect 151728 30330 151780 30336
rect 152188 30388 152240 30394
rect 152188 30330 152240 30336
rect 152924 30388 152976 30394
rect 152924 30330 152976 30336
rect 150624 6316 150676 6322
rect 150624 6258 150676 6264
rect 151636 6316 151688 6322
rect 151636 6258 151688 6264
rect 148324 5092 148376 5098
rect 148324 5034 148376 5040
rect 150348 5092 150400 5098
rect 150348 5034 150400 5040
rect 148336 480 148364 5034
rect 149520 3052 149572 3058
rect 149520 2994 149572 3000
rect 149532 480 149560 2994
rect 150636 480 150664 6258
rect 151740 5001 151768 30330
rect 152936 8702 152964 30330
rect 152924 8696 152976 8702
rect 152924 8638 152976 8644
rect 153028 6361 153056 33782
rect 153108 30456 153160 30462
rect 153108 30398 153160 30404
rect 153014 6352 153070 6361
rect 153014 6287 153070 6296
rect 153120 5030 153148 30398
rect 153856 30394 153884 34054
rect 153844 30388 153896 30394
rect 153844 30330 153896 30336
rect 154396 30388 154448 30394
rect 154396 30330 154448 30336
rect 154408 8838 154436 30330
rect 154396 8832 154448 8838
rect 154396 8774 154448 8780
rect 154212 6248 154264 6254
rect 154212 6190 154264 6196
rect 151820 5024 151872 5030
rect 151726 4992 151782 5001
rect 151820 4966 151872 4972
rect 153108 5024 153160 5030
rect 153108 4966 153160 4972
rect 151726 4927 151782 4936
rect 151832 480 151860 4966
rect 153016 3120 153068 3126
rect 153016 3062 153068 3068
rect 153028 480 153056 3062
rect 154224 480 154252 6190
rect 154500 4865 154528 34054
rect 154960 30394 154988 34054
rect 155224 31612 155276 31618
rect 155224 31554 155276 31560
rect 154948 30388 155000 30394
rect 154948 30330 155000 30336
rect 154486 4856 154542 4865
rect 154486 4791 154542 4800
rect 155236 3126 155264 31554
rect 155696 8906 155724 34054
rect 155834 33810 155862 34068
rect 156400 34054 156736 34082
rect 156952 34054 157196 34082
rect 157504 34054 157840 34082
rect 158056 34054 158392 34082
rect 155834 33782 155908 33810
rect 155776 30388 155828 30394
rect 155776 30330 155828 30336
rect 155684 8900 155736 8906
rect 155684 8842 155736 8848
rect 155788 6254 155816 30330
rect 155776 6248 155828 6254
rect 155776 6190 155828 6196
rect 155880 4962 155908 33782
rect 156604 31680 156656 31686
rect 156604 31622 156656 31628
rect 155408 4956 155460 4962
rect 155408 4898 155460 4904
rect 155868 4956 155920 4962
rect 155868 4898 155920 4904
rect 155224 3120 155276 3126
rect 155224 3062 155276 3068
rect 155420 480 155448 4898
rect 156616 3058 156644 31622
rect 156708 30394 156736 34054
rect 156696 30388 156748 30394
rect 156696 30330 156748 30336
rect 157168 9654 157196 34054
rect 157812 30394 157840 34054
rect 157984 31544 158036 31550
rect 157984 31486 158036 31492
rect 157248 30388 157300 30394
rect 157248 30330 157300 30336
rect 157800 30388 157852 30394
rect 157800 30330 157852 30336
rect 157156 9648 157208 9654
rect 157156 9590 157208 9596
rect 157260 6225 157288 30330
rect 157246 6216 157302 6225
rect 157246 6151 157302 6160
rect 157800 5568 157852 5574
rect 157800 5510 157852 5516
rect 156604 3052 156656 3058
rect 156604 2994 156656 3000
rect 156604 2916 156656 2922
rect 156604 2858 156656 2864
rect 156616 480 156644 2858
rect 157812 480 157840 5510
rect 157996 2922 158024 31486
rect 158364 30462 158392 34054
rect 158548 34054 158608 34082
rect 159160 34054 159496 34082
rect 159712 34054 160048 34082
rect 160264 34054 160600 34082
rect 160816 34054 161152 34082
rect 158352 30456 158404 30462
rect 158352 30398 158404 30404
rect 158444 30388 158496 30394
rect 158444 30330 158496 30336
rect 158456 13462 158484 30330
rect 158444 13456 158496 13462
rect 158444 13398 158496 13404
rect 158548 9586 158576 34054
rect 159364 31476 159416 31482
rect 159364 31418 159416 31424
rect 158628 30456 158680 30462
rect 158628 30398 158680 30404
rect 158536 9580 158588 9586
rect 158536 9522 158588 9528
rect 158640 7002 158668 30398
rect 158628 6996 158680 7002
rect 158628 6938 158680 6944
rect 158904 4888 158956 4894
rect 158904 4830 158956 4836
rect 157984 2916 158036 2922
rect 157984 2858 158036 2864
rect 158916 480 158944 4830
rect 159376 2854 159404 31418
rect 159468 30394 159496 34054
rect 159456 30388 159508 30394
rect 159456 30330 159508 30336
rect 159916 30388 159968 30394
rect 159916 30330 159968 30336
rect 159928 13394 159956 30330
rect 159916 13388 159968 13394
rect 159916 13330 159968 13336
rect 160020 9518 160048 34054
rect 160572 30394 160600 34054
rect 160744 31748 160796 31754
rect 160744 31690 160796 31696
rect 160560 30388 160612 30394
rect 160560 30330 160612 30336
rect 160008 9512 160060 9518
rect 160008 9454 160060 9460
rect 160756 3194 160784 31690
rect 161124 30462 161152 34054
rect 161308 34054 161368 34082
rect 161920 34054 162256 34082
rect 162472 34054 162808 34082
rect 163024 34054 163360 34082
rect 163576 34054 163912 34082
rect 161112 30456 161164 30462
rect 161112 30398 161164 30404
rect 161204 30388 161256 30394
rect 161204 30330 161256 30336
rect 161216 9450 161244 30330
rect 161204 9444 161256 9450
rect 161204 9386 161256 9392
rect 161308 9314 161336 34054
rect 162228 31550 162256 34054
rect 162216 31544 162268 31550
rect 162216 31486 162268 31492
rect 161388 30456 161440 30462
rect 161388 30398 161440 30404
rect 161296 9308 161348 9314
rect 161296 9250 161348 9256
rect 161400 4894 161428 30398
rect 162780 13326 162808 34054
rect 163332 30462 163360 34054
rect 163320 30456 163372 30462
rect 163320 30398 163372 30404
rect 163884 30394 163912 34054
rect 163976 34054 164128 34082
rect 164680 34054 165016 34082
rect 165232 34054 165568 34082
rect 165876 34054 166212 34082
rect 166428 34054 166856 34082
rect 163872 30388 163924 30394
rect 163872 30330 163924 30336
rect 162768 13320 162820 13326
rect 162768 13262 162820 13268
rect 163976 13258 164004 34054
rect 164148 30456 164200 30462
rect 164148 30398 164200 30404
rect 164056 30388 164108 30394
rect 164056 30330 164108 30336
rect 163964 13252 164016 13258
rect 163964 13194 164016 13200
rect 164068 11150 164096 30330
rect 164056 11144 164108 11150
rect 164056 11086 164108 11092
rect 164160 9382 164188 30398
rect 164988 30394 165016 34054
rect 165540 31618 165568 34054
rect 165528 31612 165580 31618
rect 165528 31554 165580 31560
rect 166184 30394 166212 34054
rect 166264 31136 166316 31142
rect 166264 31078 166316 31084
rect 164976 30388 165028 30394
rect 164976 30330 165028 30336
rect 165528 30388 165580 30394
rect 165528 30330 165580 30336
rect 166172 30388 166224 30394
rect 166172 30330 166224 30336
rect 164148 9376 164200 9382
rect 164148 9318 164200 9324
rect 165540 9246 165568 30330
rect 165528 9240 165580 9246
rect 165528 9182 165580 9188
rect 166080 5704 166132 5710
rect 166080 5646 166132 5652
rect 162492 5636 162544 5642
rect 162492 5578 162544 5584
rect 161388 4888 161440 4894
rect 161388 4830 161440 4836
rect 160100 3188 160152 3194
rect 160100 3130 160152 3136
rect 160744 3188 160796 3194
rect 160744 3130 160796 3136
rect 159364 2848 159416 2854
rect 159364 2790 159416 2796
rect 160112 480 160140 3130
rect 161296 3120 161348 3126
rect 161296 3062 161348 3068
rect 161308 480 161336 3062
rect 162504 480 162532 5578
rect 163688 4820 163740 4826
rect 163688 4762 163740 4768
rect 163700 480 163728 4762
rect 164884 3052 164936 3058
rect 164884 2994 164936 3000
rect 164896 480 164924 2994
rect 166092 480 166120 5646
rect 166276 2990 166304 31078
rect 166828 9178 166856 34054
rect 166920 34054 166980 34082
rect 167532 34054 167960 34082
rect 168084 34054 168328 34082
rect 168636 34054 168972 34082
rect 169188 34054 169616 34082
rect 166920 31482 166948 34054
rect 166908 31476 166960 31482
rect 166908 31418 166960 31424
rect 167644 31204 167696 31210
rect 167644 31146 167696 31152
rect 166908 30388 166960 30394
rect 166908 30330 166960 30336
rect 166816 9172 166868 9178
rect 166816 9114 166868 9120
rect 166920 4826 166948 30330
rect 166908 4820 166960 4826
rect 166908 4762 166960 4768
rect 167184 3256 167236 3262
rect 167184 3198 167236 3204
rect 166264 2984 166316 2990
rect 166264 2926 166316 2932
rect 167196 480 167224 3198
rect 167656 3058 167684 31146
rect 167932 26234 167960 34054
rect 167932 26206 168236 26234
rect 168208 12510 168236 26206
rect 168196 12504 168248 12510
rect 168196 12446 168248 12452
rect 168300 9042 168328 34054
rect 168944 31142 168972 34054
rect 169024 31340 169076 31346
rect 169024 31282 169076 31288
rect 168932 31136 168984 31142
rect 168932 31078 168984 31084
rect 168288 9036 168340 9042
rect 168288 8978 168340 8984
rect 167644 3052 167696 3058
rect 167644 2994 167696 3000
rect 169036 2922 169064 31282
rect 169588 13190 169616 34054
rect 169680 34054 169740 34082
rect 170292 34054 170628 34082
rect 170844 34054 171088 34082
rect 171396 34054 171732 34082
rect 171948 34054 172284 34082
rect 169576 13184 169628 13190
rect 169576 13126 169628 13132
rect 169680 8974 169708 34054
rect 170404 31408 170456 31414
rect 170404 31350 170456 31356
rect 169668 8968 169720 8974
rect 169668 8910 169720 8916
rect 169576 5772 169628 5778
rect 169576 5714 169628 5720
rect 168380 2916 168432 2922
rect 168380 2858 168432 2864
rect 169024 2916 169076 2922
rect 169024 2858 169076 2864
rect 168392 480 168420 2858
rect 169588 480 169616 5714
rect 170416 3194 170444 31350
rect 170600 30462 170628 34054
rect 170588 30456 170640 30462
rect 170588 30398 170640 30404
rect 171060 13122 171088 34054
rect 171704 30394 171732 34054
rect 172256 30530 172284 34054
rect 172348 34054 172500 34082
rect 173052 34054 173388 34082
rect 173604 34054 173756 34082
rect 174156 34054 174492 34082
rect 174708 34054 175136 34082
rect 172244 30524 172296 30530
rect 172244 30466 172296 30472
rect 171692 30388 171744 30394
rect 171692 30330 171744 30336
rect 171048 13116 171100 13122
rect 171048 13058 171100 13064
rect 172348 12646 172376 34054
rect 173164 30796 173216 30802
rect 173164 30738 173216 30744
rect 172428 30388 172480 30394
rect 172428 30330 172480 30336
rect 172336 12640 172388 12646
rect 172336 12582 172388 12588
rect 172440 8362 172468 30330
rect 173176 16574 173204 30738
rect 173360 30394 173388 34054
rect 173348 30388 173400 30394
rect 173348 30330 173400 30336
rect 173176 16546 173296 16574
rect 172428 8356 172480 8362
rect 172428 8298 172480 8304
rect 173164 5908 173216 5914
rect 173164 5850 173216 5856
rect 170772 5840 170824 5846
rect 170772 5782 170824 5788
rect 170404 3188 170456 3194
rect 170404 3130 170456 3136
rect 170784 480 170812 5782
rect 171968 2848 172020 2854
rect 171968 2790 172020 2796
rect 171980 480 172008 2790
rect 173176 480 173204 5850
rect 173268 2854 173296 16546
rect 173728 13870 173756 34054
rect 174464 30394 174492 34054
rect 173808 30388 173860 30394
rect 173808 30330 173860 30336
rect 174452 30388 174504 30394
rect 174452 30330 174504 30336
rect 175004 30388 175056 30394
rect 175004 30330 175056 30336
rect 173716 13864 173768 13870
rect 173716 13806 173768 13812
rect 173820 9110 173848 30330
rect 175016 26234 175044 30330
rect 175108 30138 175136 34054
rect 175200 34054 175260 34082
rect 175812 34054 176148 34082
rect 176456 34054 176608 34082
rect 177008 34054 177344 34082
rect 177560 34054 177988 34082
rect 178112 34054 178448 34082
rect 178664 34054 179000 34082
rect 179216 34054 179368 34082
rect 179768 34054 180104 34082
rect 180320 34054 180564 34082
rect 180872 34054 181208 34082
rect 181424 34054 181760 34082
rect 175200 30734 175228 34054
rect 175924 31068 175976 31074
rect 175924 31010 175976 31016
rect 175188 30728 175240 30734
rect 175188 30670 175240 30676
rect 175108 30110 175228 30138
rect 175016 26206 175136 26234
rect 175108 12578 175136 26206
rect 175096 12572 175148 12578
rect 175096 12514 175148 12520
rect 173808 9104 173860 9110
rect 173808 9046 173860 9052
rect 175200 8430 175228 30110
rect 175188 8424 175240 8430
rect 175188 8366 175240 8372
rect 174268 3324 174320 3330
rect 174268 3266 174320 3272
rect 173256 2848 173308 2854
rect 173256 2790 173308 2796
rect 174280 480 174308 3266
rect 175936 3262 175964 31010
rect 176120 26234 176148 34054
rect 176120 26206 176516 26234
rect 176488 12714 176516 26206
rect 176476 12708 176528 12714
rect 176476 12650 176528 12656
rect 176580 9353 176608 34054
rect 177212 30660 177264 30666
rect 177212 30602 177264 30608
rect 177224 26234 177252 30602
rect 177316 30394 177344 34054
rect 177396 31000 177448 31006
rect 177396 30942 177448 30948
rect 177304 30388 177356 30394
rect 177304 30330 177356 30336
rect 177224 26206 177344 26234
rect 176566 9344 176622 9353
rect 176566 9279 176622 9288
rect 176660 6180 176712 6186
rect 176660 6122 176712 6128
rect 175924 3256 175976 3262
rect 175924 3198 175976 3204
rect 175464 3120 175516 3126
rect 175464 3062 175516 3068
rect 175476 480 175504 3062
rect 176672 480 176700 6122
rect 177316 3126 177344 26206
rect 177408 3330 177436 30942
rect 177856 30388 177908 30394
rect 177856 30330 177908 30336
rect 177868 13938 177896 30330
rect 177856 13932 177908 13938
rect 177856 13874 177908 13880
rect 177960 12782 177988 34054
rect 178420 30394 178448 34054
rect 178972 30666 179000 34054
rect 178960 30660 179012 30666
rect 178960 30602 179012 30608
rect 178408 30388 178460 30394
rect 178408 30330 178460 30336
rect 179236 30388 179288 30394
rect 179236 30330 179288 30336
rect 177948 12776 178000 12782
rect 177948 12718 178000 12724
rect 179248 9217 179276 30330
rect 179234 9208 179290 9217
rect 179234 9143 179290 9152
rect 179340 6186 179368 34054
rect 179972 30932 180024 30938
rect 179972 30874 180024 30880
rect 179984 26234 180012 30874
rect 180076 30394 180104 34054
rect 180536 31074 180564 34054
rect 180524 31068 180576 31074
rect 180524 31010 180576 31016
rect 181180 30598 181208 34054
rect 181444 30864 181496 30870
rect 181444 30806 181496 30812
rect 181168 30592 181220 30598
rect 181168 30534 181220 30540
rect 180064 30388 180116 30394
rect 180064 30330 180116 30336
rect 180708 30388 180760 30394
rect 180708 30330 180760 30336
rect 179984 26206 180104 26234
rect 179328 6180 179380 6186
rect 179328 6122 179380 6128
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 177396 3324 177448 3330
rect 177396 3266 177448 3272
rect 177304 3120 177356 3126
rect 177304 3062 177356 3068
rect 177868 480 177896 3334
rect 180076 2990 180104 26206
rect 180720 9081 180748 30330
rect 181456 16574 181484 30806
rect 181732 30394 181760 34054
rect 181916 34054 181976 34082
rect 182528 34054 182864 34082
rect 183080 34054 183416 34082
rect 183632 34054 183968 34082
rect 184184 34054 184520 34082
rect 181720 30388 181772 30394
rect 181720 30330 181772 30336
rect 181456 16546 181576 16574
rect 180706 9072 180762 9081
rect 180706 9007 180762 9016
rect 180248 6044 180300 6050
rect 180248 5986 180300 5992
rect 179052 2984 179104 2990
rect 179052 2926 179104 2932
rect 180064 2984 180116 2990
rect 180064 2926 180116 2932
rect 179064 480 179092 2926
rect 180260 480 180288 5986
rect 181444 5976 181496 5982
rect 181444 5918 181496 5924
rect 181456 480 181484 5918
rect 181548 3126 181576 16546
rect 181916 14074 181944 34054
rect 182088 30592 182140 30598
rect 182088 30534 182140 30540
rect 181996 30388 182048 30394
rect 181996 30330 182048 30336
rect 181904 14068 181956 14074
rect 181904 14010 181956 14016
rect 182008 14006 182036 30330
rect 181996 14000 182048 14006
rect 181996 13942 182048 13948
rect 182100 5574 182128 30534
rect 182836 30394 182864 34054
rect 182824 30388 182876 30394
rect 182824 30330 182876 30336
rect 183388 14142 183416 34054
rect 183940 30598 183968 34054
rect 183928 30592 183980 30598
rect 183928 30534 183980 30540
rect 184492 30394 184520 34054
rect 184676 34054 184736 34082
rect 185288 34054 185624 34082
rect 185840 34054 186268 34082
rect 186392 34054 186728 34082
rect 187036 34054 187372 34082
rect 183468 30388 183520 30394
rect 183468 30330 183520 30336
rect 184480 30388 184532 30394
rect 184480 30330 184532 30336
rect 183376 14136 183428 14142
rect 183376 14078 183428 14084
rect 183480 5642 183508 30330
rect 184676 14278 184704 34054
rect 185492 31068 185544 31074
rect 185492 31010 185544 31016
rect 184848 30592 184900 30598
rect 184848 30534 184900 30540
rect 184756 30388 184808 30394
rect 184756 30330 184808 30336
rect 184664 14272 184716 14278
rect 184664 14214 184716 14220
rect 183744 6112 183796 6118
rect 183744 6054 183796 6060
rect 183468 5636 183520 5642
rect 183468 5578 183520 5584
rect 182088 5568 182140 5574
rect 182088 5510 182140 5516
rect 181536 3120 181588 3126
rect 181536 3062 181588 3068
rect 182548 3052 182600 3058
rect 182548 2994 182600 3000
rect 182560 480 182588 2994
rect 183756 480 183784 6054
rect 184768 5710 184796 30330
rect 184756 5704 184808 5710
rect 184756 5646 184808 5652
rect 184860 3058 184888 30534
rect 185504 26234 185532 31010
rect 185596 30802 185624 34054
rect 185584 30796 185636 30802
rect 185584 30738 185636 30744
rect 185504 26206 185624 26234
rect 185596 4146 185624 26206
rect 186240 5778 186268 34054
rect 186700 30394 186728 34054
rect 187344 30598 187372 34054
rect 187528 34054 187588 34082
rect 188140 34054 188476 34082
rect 188692 34054 189028 34082
rect 189244 34054 189580 34082
rect 189796 34054 190224 34082
rect 187332 30592 187384 30598
rect 187332 30534 187384 30540
rect 186688 30388 186740 30394
rect 186688 30330 186740 30336
rect 187424 30388 187476 30394
rect 187424 30330 187476 30336
rect 187436 14210 187464 30330
rect 187424 14204 187476 14210
rect 187424 14146 187476 14152
rect 187332 6792 187384 6798
rect 187332 6734 187384 6740
rect 186228 5772 186280 5778
rect 186228 5714 186280 5720
rect 184940 4140 184992 4146
rect 184940 4082 184992 4088
rect 185584 4140 185636 4146
rect 185584 4082 185636 4088
rect 184848 3052 184900 3058
rect 184848 2994 184900 3000
rect 184952 480 184980 4082
rect 186136 2916 186188 2922
rect 186136 2858 186188 2864
rect 186148 480 186176 2858
rect 187344 480 187372 6734
rect 187528 5846 187556 34054
rect 188448 30870 188476 34054
rect 189000 31754 189028 34054
rect 188988 31748 189040 31754
rect 188988 31690 189040 31696
rect 188436 30864 188488 30870
rect 188436 30806 188488 30812
rect 188988 30864 189040 30870
rect 188988 30806 189040 30812
rect 187608 30592 187660 30598
rect 187608 30534 187660 30540
rect 187516 5840 187568 5846
rect 187516 5782 187568 5788
rect 187620 3058 187648 30534
rect 189000 9790 189028 30806
rect 189552 30394 189580 34054
rect 189540 30388 189592 30394
rect 189540 30330 189592 30336
rect 190196 9858 190224 34054
rect 190334 33810 190362 34068
rect 190900 34054 191236 34082
rect 191452 34054 191696 34082
rect 192004 34054 192340 34082
rect 192556 34054 192892 34082
rect 190334 33782 190408 33810
rect 190276 30388 190328 30394
rect 190276 30330 190328 30336
rect 190184 9852 190236 9858
rect 190184 9794 190236 9800
rect 188988 9784 189040 9790
rect 188988 9726 189040 9732
rect 190288 5914 190316 30330
rect 190276 5908 190328 5914
rect 190276 5850 190328 5856
rect 188528 4072 188580 4078
rect 188528 4014 188580 4020
rect 187608 3052 187660 3058
rect 187608 2994 187660 3000
rect 188540 480 188568 4014
rect 190380 3194 190408 33782
rect 191208 30394 191236 34054
rect 191196 30388 191248 30394
rect 191196 30330 191248 30336
rect 191668 9926 191696 34054
rect 192312 31006 192340 34054
rect 192300 31000 192352 31006
rect 192300 30942 192352 30948
rect 192864 30394 192892 34054
rect 193048 34054 193108 34082
rect 193660 34054 193996 34082
rect 194212 34054 194456 34082
rect 194764 34054 195100 34082
rect 195316 34054 195652 34082
rect 191748 30388 191800 30394
rect 191748 30330 191800 30336
rect 192852 30388 192904 30394
rect 192852 30330 192904 30336
rect 191656 9920 191708 9926
rect 191656 9862 191708 9868
rect 190828 6724 190880 6730
rect 190828 6666 190880 6672
rect 189724 3188 189776 3194
rect 189724 3130 189776 3136
rect 190368 3188 190420 3194
rect 190368 3130 190420 3136
rect 189736 480 189764 3130
rect 190840 480 190868 6666
rect 191760 5982 191788 30330
rect 193048 9994 193076 34054
rect 193968 30394 193996 34054
rect 193128 30388 193180 30394
rect 193128 30330 193180 30336
rect 193956 30388 194008 30394
rect 193956 30330 194008 30336
rect 193036 9988 193088 9994
rect 193036 9930 193088 9936
rect 193140 6050 193168 30330
rect 194324 6656 194376 6662
rect 194324 6598 194376 6604
rect 193128 6044 193180 6050
rect 193128 5986 193180 5992
rect 191748 5976 191800 5982
rect 191748 5918 191800 5924
rect 192024 3936 192076 3942
rect 192024 3878 192076 3884
rect 192036 480 192064 3878
rect 194336 3346 194364 6598
rect 194428 6118 194456 34054
rect 195072 30870 195100 34054
rect 195624 30938 195652 34054
rect 195854 33810 195882 34068
rect 196420 34054 196756 34082
rect 196972 34054 197308 34082
rect 197616 34054 197952 34082
rect 198168 34054 198596 34082
rect 195854 33782 195928 33810
rect 195612 30932 195664 30938
rect 195612 30874 195664 30880
rect 195060 30864 195112 30870
rect 195060 30806 195112 30812
rect 195796 30864 195848 30870
rect 195796 30806 195848 30812
rect 194508 30388 194560 30394
rect 194508 30330 194560 30336
rect 194416 6112 194468 6118
rect 194416 6054 194468 6060
rect 194520 3942 194548 30330
rect 195808 10062 195836 30806
rect 195796 10056 195848 10062
rect 195796 9998 195848 10004
rect 195900 5273 195928 33782
rect 196728 30394 196756 34054
rect 196716 30388 196768 30394
rect 196716 30330 196768 30336
rect 197176 30388 197228 30394
rect 197176 30330 197228 30336
rect 197188 10130 197216 30330
rect 197176 10124 197228 10130
rect 197176 10066 197228 10072
rect 195886 5264 195942 5273
rect 195886 5199 195942 5208
rect 195612 4004 195664 4010
rect 195612 3946 195664 3952
rect 194508 3936 194560 3942
rect 194508 3878 194560 3884
rect 193220 3324 193272 3330
rect 194336 3318 194456 3346
rect 193220 3266 193272 3272
rect 193232 480 193260 3266
rect 194428 480 194456 3318
rect 195624 480 195652 3946
rect 197280 3330 197308 34054
rect 197924 30394 197952 34054
rect 197912 30388 197964 30394
rect 197912 30330 197964 30336
rect 198568 10198 198596 34054
rect 198660 34054 198720 34082
rect 199272 34054 199608 34082
rect 199824 34054 199976 34082
rect 200376 34054 200712 34082
rect 200928 34054 201356 34082
rect 198660 31346 198688 34054
rect 198648 31340 198700 31346
rect 198648 31282 198700 31288
rect 199580 30394 199608 34054
rect 198648 30388 198700 30394
rect 198648 30330 198700 30336
rect 199568 30388 199620 30394
rect 199568 30330 199620 30336
rect 198556 10192 198608 10198
rect 198556 10134 198608 10140
rect 198660 6798 198688 30330
rect 199948 10266 199976 34054
rect 200684 30394 200712 34054
rect 200764 31680 200816 31686
rect 200764 31622 200816 31628
rect 200028 30388 200080 30394
rect 200028 30330 200080 30336
rect 200672 30388 200724 30394
rect 200672 30330 200724 30336
rect 199936 10260 199988 10266
rect 199936 10202 199988 10208
rect 198648 6792 198700 6798
rect 198648 6734 198700 6740
rect 200040 6730 200068 30330
rect 200028 6724 200080 6730
rect 200028 6666 200080 6672
rect 197912 6588 197964 6594
rect 197912 6530 197964 6536
rect 197268 3324 197320 3330
rect 197268 3266 197320 3272
rect 196808 2916 196860 2922
rect 196808 2858 196860 2864
rect 196820 480 196848 2858
rect 197924 480 197952 6530
rect 200776 4214 200804 31622
rect 201224 30388 201276 30394
rect 201224 30330 201276 30336
rect 201236 11014 201264 30330
rect 201224 11008 201276 11014
rect 201224 10950 201276 10956
rect 201328 6662 201356 34054
rect 201420 34054 201480 34082
rect 202032 34054 202368 34082
rect 202584 34054 202828 34082
rect 203136 34054 203472 34082
rect 203688 34054 203932 34082
rect 201420 30394 201448 34054
rect 202340 31006 202368 34054
rect 202328 31000 202380 31006
rect 202328 30942 202380 30948
rect 201408 30388 201460 30394
rect 201408 30330 201460 30336
rect 201408 30252 201460 30258
rect 201408 30194 201460 30200
rect 201316 6656 201368 6662
rect 201316 6598 201368 6604
rect 200304 4208 200356 4214
rect 200304 4150 200356 4156
rect 200764 4208 200816 4214
rect 200764 4150 200816 4156
rect 199108 3868 199160 3874
rect 199108 3810 199160 3816
rect 199120 480 199148 3810
rect 200316 480 200344 4150
rect 201420 4146 201448 30194
rect 202800 12850 202828 34054
rect 203444 30598 203472 34054
rect 203432 30592 203484 30598
rect 203432 30534 203484 30540
rect 203904 30394 203932 34054
rect 203996 34054 204240 34082
rect 204792 34054 205128 34082
rect 205344 34054 205588 34082
rect 205896 34054 206232 34082
rect 206448 34054 206876 34082
rect 203892 30388 203944 30394
rect 203892 30330 203944 30336
rect 203996 12918 204024 34054
rect 204904 31612 204956 31618
rect 204904 31554 204956 31560
rect 204076 30592 204128 30598
rect 204076 30534 204128 30540
rect 203984 12912 204036 12918
rect 203984 12854 204036 12860
rect 202788 12844 202840 12850
rect 202788 12786 202840 12792
rect 204088 10946 204116 30534
rect 204168 30388 204220 30394
rect 204168 30330 204220 30336
rect 204076 10940 204128 10946
rect 204076 10882 204128 10888
rect 201500 8220 201552 8226
rect 201500 8162 201552 8168
rect 201408 4140 201460 4146
rect 201408 4082 201460 4088
rect 201512 480 201540 8162
rect 203892 4480 203944 4486
rect 203892 4422 203944 4428
rect 202696 3868 202748 3874
rect 202696 3810 202748 3816
rect 202708 480 202736 3810
rect 203904 480 203932 4422
rect 204180 4078 204208 30330
rect 204916 4486 204944 31554
rect 205100 30394 205128 34054
rect 205560 31550 205588 34054
rect 205548 31544 205600 31550
rect 205548 31486 205600 31492
rect 206204 30394 206232 34054
rect 205088 30388 205140 30394
rect 205088 30330 205140 30336
rect 205548 30388 205600 30394
rect 205548 30330 205600 30336
rect 206192 30388 206244 30394
rect 206192 30330 206244 30336
rect 206744 30388 206796 30394
rect 206744 30330 206796 30336
rect 205560 10878 205588 30330
rect 206756 14346 206784 30330
rect 206744 14340 206796 14346
rect 206744 14282 206796 14288
rect 205548 10872 205600 10878
rect 205548 10814 205600 10820
rect 206848 10810 206876 34054
rect 206940 34054 207000 34082
rect 207552 34054 208072 34082
rect 208196 34054 208348 34082
rect 208748 34054 209084 34082
rect 209300 34054 209728 34082
rect 209852 34054 210188 34082
rect 210404 34054 210740 34082
rect 206836 10804 206888 10810
rect 206836 10746 206888 10752
rect 205088 8152 205140 8158
rect 205088 8094 205140 8100
rect 204904 4480 204956 4486
rect 204904 4422 204956 4428
rect 204168 4072 204220 4078
rect 204168 4014 204220 4020
rect 205100 480 205128 8094
rect 206940 4010 206968 34054
rect 208044 26234 208072 34054
rect 208044 26206 208256 26234
rect 208228 14414 208256 26206
rect 208216 14408 208268 14414
rect 208216 14350 208268 14356
rect 208320 10742 208348 34054
rect 209056 31618 209084 34054
rect 209044 31612 209096 31618
rect 209044 31554 209096 31560
rect 209044 31476 209096 31482
rect 209044 31418 209096 31424
rect 208308 10736 208360 10742
rect 208308 10678 208360 10684
rect 208584 8084 208636 8090
rect 208584 8026 208636 8032
rect 207388 4344 207440 4350
rect 207388 4286 207440 4292
rect 206192 4004 206244 4010
rect 206192 3946 206244 3952
rect 206928 4004 206980 4010
rect 206928 3946 206980 3952
rect 206204 480 206232 3946
rect 207400 480 207428 4286
rect 208596 480 208624 8026
rect 209056 4350 209084 31418
rect 209700 7070 209728 34054
rect 210160 30394 210188 34054
rect 210712 30598 210740 34054
rect 210942 33810 210970 34068
rect 211508 34054 211844 34082
rect 212060 34054 212396 34082
rect 212612 34054 212948 34082
rect 213164 34054 213592 34082
rect 213716 34054 213868 34082
rect 214268 34054 214604 34082
rect 214820 34054 215156 34082
rect 215372 34054 215708 34082
rect 215924 34054 216260 34082
rect 210942 33782 211016 33810
rect 210700 30592 210752 30598
rect 210700 30534 210752 30540
rect 210148 30388 210200 30394
rect 210148 30330 210200 30336
rect 210884 30388 210936 30394
rect 210884 30330 210936 30336
rect 210896 10674 210924 30330
rect 210884 10668 210936 10674
rect 210884 10610 210936 10616
rect 210988 7138 211016 33782
rect 211068 30592 211120 30598
rect 211068 30534 211120 30540
rect 210976 7132 211028 7138
rect 210976 7074 211028 7080
rect 209688 7064 209740 7070
rect 209688 7006 209740 7012
rect 210976 4412 211028 4418
rect 210976 4354 211028 4360
rect 209044 4344 209096 4350
rect 209044 4286 209096 4292
rect 209780 3800 209832 3806
rect 209780 3742 209832 3748
rect 209792 480 209820 3742
rect 210988 480 211016 4354
rect 211080 3942 211108 30534
rect 211816 30394 211844 34054
rect 212368 31210 212396 34054
rect 212356 31204 212408 31210
rect 212356 31146 212408 31152
rect 212920 30394 212948 34054
rect 213184 31136 213236 31142
rect 213184 31078 213236 31084
rect 211804 30388 211856 30394
rect 211804 30330 211856 30336
rect 212448 30388 212500 30394
rect 212448 30330 212500 30336
rect 212908 30388 212960 30394
rect 212908 30330 212960 30336
rect 212460 10606 212488 30330
rect 212448 10600 212500 10606
rect 212448 10542 212500 10548
rect 213196 4418 213224 31078
rect 213564 26234 213592 34054
rect 213736 30388 213788 30394
rect 213736 30330 213788 30336
rect 213564 26206 213684 26234
rect 213656 10538 213684 26206
rect 213644 10532 213696 10538
rect 213644 10474 213696 10480
rect 213748 7206 213776 30330
rect 213736 7200 213788 7206
rect 213736 7142 213788 7148
rect 213184 4412 213236 4418
rect 213184 4354 213236 4360
rect 211068 3936 211120 3942
rect 211068 3878 211120 3884
rect 213840 3874 213868 34054
rect 214576 30394 214604 34054
rect 214564 30388 214616 30394
rect 214564 30330 214616 30336
rect 215128 10470 215156 34054
rect 215680 31686 215708 34054
rect 215668 31680 215720 31686
rect 215668 31622 215720 31628
rect 216232 30394 216260 34054
rect 216462 33810 216490 34068
rect 217028 34054 217364 34082
rect 217580 34054 217916 34082
rect 218132 34054 218468 34082
rect 218776 34054 219112 34082
rect 216462 33782 216536 33810
rect 215208 30388 215260 30394
rect 215208 30330 215260 30336
rect 216220 30388 216272 30394
rect 216220 30330 216272 30336
rect 215116 10464 215168 10470
rect 215116 10406 215168 10412
rect 215220 7274 215248 30330
rect 216508 10402 216536 33782
rect 217336 30394 217364 34054
rect 216588 30388 216640 30394
rect 216588 30330 216640 30336
rect 217324 30388 217376 30394
rect 217324 30330 217376 30336
rect 216496 10396 216548 10402
rect 216496 10338 216548 10344
rect 215668 7948 215720 7954
rect 215668 7890 215720 7896
rect 215208 7268 215260 7274
rect 215208 7210 215260 7216
rect 214472 4276 214524 4282
rect 214472 4218 214524 4224
rect 213828 3868 213880 3874
rect 213828 3810 213880 3816
rect 212172 3664 212224 3670
rect 212172 3606 212224 3612
rect 212184 480 212212 3606
rect 213368 3596 213420 3602
rect 213368 3538 213420 3544
rect 213380 480 213408 3538
rect 214484 480 214512 4218
rect 215680 480 215708 7890
rect 216600 7342 216628 30330
rect 217888 7410 217916 34054
rect 218440 30394 218468 34054
rect 219084 31414 219112 34054
rect 219314 33810 219342 34068
rect 219880 34054 220216 34082
rect 220432 34054 220768 34082
rect 220984 34054 221320 34082
rect 221536 34054 221964 34082
rect 219314 33782 219388 33810
rect 219072 31408 219124 31414
rect 219072 31350 219124 31356
rect 217968 30388 218020 30394
rect 217968 30330 218020 30336
rect 218428 30388 218480 30394
rect 218428 30330 218480 30336
rect 219256 30388 219308 30394
rect 219256 30330 219308 30336
rect 217876 7404 217928 7410
rect 217876 7346 217928 7352
rect 216588 7336 216640 7342
rect 216588 7278 216640 7284
rect 217980 3806 218008 30330
rect 219268 10334 219296 30330
rect 219256 10328 219308 10334
rect 219256 10270 219308 10276
rect 219256 8016 219308 8022
rect 219256 7958 219308 7964
rect 218060 4548 218112 4554
rect 218060 4490 218112 4496
rect 217968 3800 218020 3806
rect 216862 3768 216918 3777
rect 217968 3742 218020 3748
rect 216862 3703 216918 3712
rect 216876 480 216904 3703
rect 218072 480 218100 4490
rect 219268 480 219296 7958
rect 219360 7478 219388 33782
rect 220188 30394 220216 34054
rect 220176 30388 220228 30394
rect 220176 30330 220228 30336
rect 220636 30388 220688 30394
rect 220636 30330 220688 30336
rect 220648 10713 220676 30330
rect 220634 10704 220690 10713
rect 220634 10639 220690 10648
rect 219348 7472 219400 7478
rect 219348 7414 219400 7420
rect 220740 3738 220768 34054
rect 221292 30394 221320 34054
rect 221280 30388 221332 30394
rect 221280 30330 221332 30336
rect 221936 26234 221964 34054
rect 222028 34054 222088 34082
rect 222640 34054 222976 34082
rect 223192 34054 223436 34082
rect 223744 34054 224080 34082
rect 224296 34054 224632 34082
rect 222028 31142 222056 34054
rect 222016 31136 222068 31142
rect 222016 31078 222068 31084
rect 222948 30394 222976 34054
rect 222108 30388 222160 30394
rect 222108 30330 222160 30336
rect 222936 30388 222988 30394
rect 222936 30330 222988 30336
rect 221936 26206 222056 26234
rect 222028 10577 222056 26206
rect 222014 10568 222070 10577
rect 222014 10503 222070 10512
rect 222120 7546 222148 30330
rect 223408 10441 223436 34054
rect 224052 30598 224080 34054
rect 224040 30592 224092 30598
rect 224040 30534 224092 30540
rect 224604 30394 224632 34054
rect 224696 34054 224848 34082
rect 225400 34054 225736 34082
rect 225952 34054 226288 34082
rect 226504 34054 226840 34082
rect 227056 34054 227392 34082
rect 223488 30388 223540 30394
rect 223488 30330 223540 30336
rect 224592 30388 224644 30394
rect 224592 30330 224644 30336
rect 223394 10432 223450 10441
rect 223394 10367 223450 10376
rect 223500 8294 223528 30330
rect 224696 10305 224724 34054
rect 225708 31278 225736 34054
rect 225696 31272 225748 31278
rect 225696 31214 225748 31220
rect 224868 30592 224920 30598
rect 224868 30534 224920 30540
rect 224776 30388 224828 30394
rect 224776 30330 224828 30336
rect 224682 10296 224738 10305
rect 224682 10231 224738 10240
rect 223488 8288 223540 8294
rect 223488 8230 223540 8236
rect 224788 8226 224816 30330
rect 224776 8220 224828 8226
rect 224776 8162 224828 8168
rect 222752 7880 222804 7886
rect 222752 7822 222804 7828
rect 222108 7540 222160 7546
rect 222108 7482 222160 7488
rect 221556 4616 221608 4622
rect 221556 4558 221608 4564
rect 220728 3732 220780 3738
rect 220728 3674 220780 3680
rect 220452 3528 220504 3534
rect 220452 3470 220504 3476
rect 220464 480 220492 3470
rect 221568 480 221596 4558
rect 222764 480 222792 7822
rect 224880 3670 224908 30534
rect 226260 8158 226288 34054
rect 226812 30394 226840 34054
rect 227364 30598 227392 34054
rect 227548 34054 227608 34082
rect 228160 34054 228496 34082
rect 228712 34054 228956 34082
rect 229356 34054 229692 34082
rect 229908 34054 230244 34082
rect 227352 30592 227404 30598
rect 227352 30534 227404 30540
rect 226800 30388 226852 30394
rect 226800 30330 226852 30336
rect 227444 30388 227496 30394
rect 227444 30330 227496 30336
rect 227456 15162 227484 30330
rect 227444 15156 227496 15162
rect 227444 15098 227496 15104
rect 226248 8152 226300 8158
rect 226248 8094 226300 8100
rect 227548 8022 227576 34054
rect 227628 30592 227680 30598
rect 227628 30534 227680 30540
rect 227536 8016 227588 8022
rect 227536 7958 227588 7964
rect 226340 7812 226392 7818
rect 226340 7754 226392 7760
rect 225144 4684 225196 4690
rect 225144 4626 225196 4632
rect 224868 3664 224920 3670
rect 223946 3632 224002 3641
rect 224868 3606 224920 3612
rect 223946 3567 224002 3576
rect 223960 480 223988 3567
rect 225156 480 225184 4626
rect 226352 480 226380 7754
rect 227640 3602 227668 30534
rect 228468 30394 228496 34054
rect 228928 31074 228956 34054
rect 228916 31068 228968 31074
rect 228916 31010 228968 31016
rect 229664 30394 229692 34054
rect 228456 30388 228508 30394
rect 228456 30330 228508 30336
rect 229008 30388 229060 30394
rect 229008 30330 229060 30336
rect 229652 30388 229704 30394
rect 229652 30330 229704 30336
rect 229020 15094 229048 30330
rect 229008 15088 229060 15094
rect 229008 15030 229060 15036
rect 230216 15026 230244 34054
rect 230400 34054 230460 34082
rect 231012 34054 231348 34082
rect 231564 34054 231716 34082
rect 232116 34054 232452 34082
rect 232668 34054 233004 34082
rect 230296 30388 230348 30394
rect 230296 30330 230348 30336
rect 230204 15020 230256 15026
rect 230204 14962 230256 14968
rect 230308 8090 230336 30330
rect 230296 8084 230348 8090
rect 230296 8026 230348 8032
rect 228732 4752 228784 4758
rect 228732 4694 228784 4700
rect 227628 3596 227680 3602
rect 227628 3538 227680 3544
rect 227534 3496 227590 3505
rect 227534 3431 227590 3440
rect 227548 480 227576 3431
rect 228744 480 228772 4694
rect 230400 3534 230428 34054
rect 231320 30394 231348 34054
rect 231308 30388 231360 30394
rect 231308 30330 231360 30336
rect 231688 14958 231716 34054
rect 232424 30598 232452 34054
rect 232412 30592 232464 30598
rect 232412 30534 232464 30540
rect 232976 30394 233004 34054
rect 233068 34054 233220 34082
rect 233772 34054 234200 34082
rect 234324 34054 234568 34082
rect 234876 34054 235212 34082
rect 235428 34054 235764 34082
rect 231768 30388 231820 30394
rect 231768 30330 231820 30336
rect 232964 30388 233016 30394
rect 232964 30330 233016 30336
rect 231676 14952 231728 14958
rect 231676 14894 231728 14900
rect 231780 7954 231808 30330
rect 233068 14890 233096 34054
rect 233148 30388 233200 30394
rect 233148 30330 233200 30336
rect 233056 14884 233108 14890
rect 233056 14826 233108 14832
rect 231768 7948 231820 7954
rect 231768 7890 231820 7896
rect 233160 7886 233188 30330
rect 234172 26234 234200 34054
rect 234172 26206 234476 26234
rect 234448 16114 234476 26206
rect 234436 16108 234488 16114
rect 234436 16050 234488 16056
rect 233148 7880 233200 7886
rect 233148 7822 233200 7828
rect 234540 7818 234568 34054
rect 235184 30394 235212 34054
rect 235172 30388 235224 30394
rect 235172 30330 235224 30336
rect 235736 30326 235764 34054
rect 235920 34054 235980 34082
rect 236532 34054 236960 34082
rect 237084 34054 237328 34082
rect 237636 34054 237972 34082
rect 238188 34054 238616 34082
rect 235816 30388 235868 30394
rect 235816 30330 235868 30336
rect 235724 30320 235776 30326
rect 235724 30262 235776 30268
rect 235828 11218 235856 30330
rect 235816 11212 235868 11218
rect 235816 11154 235868 11160
rect 234528 7812 234580 7818
rect 234528 7754 234580 7760
rect 235920 7750 235948 34054
rect 236932 26234 236960 34054
rect 236932 26206 237236 26234
rect 234620 7744 234672 7750
rect 234620 7686 234672 7692
rect 235908 7744 235960 7750
rect 235908 7686 235960 7692
rect 232228 5500 232280 5506
rect 232228 5442 232280 5448
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 231032 3460 231084 3466
rect 231032 3402 231084 3408
rect 229836 2848 229888 2854
rect 229836 2790 229888 2796
rect 229848 480 229876 2790
rect 231044 480 231072 3402
rect 232240 480 232268 5442
rect 233424 2984 233476 2990
rect 233424 2926 233476 2932
rect 233436 480 233464 2926
rect 234632 480 234660 7686
rect 237208 6594 237236 26206
rect 237196 6588 237248 6594
rect 237196 6530 237248 6536
rect 235814 5128 235870 5137
rect 235814 5063 235870 5072
rect 235828 480 235856 5063
rect 237300 3466 237328 34054
rect 237944 31482 237972 34054
rect 237932 31476 237984 31482
rect 237932 31418 237984 31424
rect 238588 11286 238616 34054
rect 238680 34054 238740 34082
rect 239292 34054 239628 34082
rect 238680 31634 238708 34054
rect 238680 31606 238800 31634
rect 238668 31476 238720 31482
rect 238668 31418 238720 31424
rect 238576 11280 238628 11286
rect 238576 11222 238628 11228
rect 238680 7993 238708 31418
rect 238772 30977 238800 31606
rect 238758 30968 238814 30977
rect 238758 30903 238814 30912
rect 239600 30394 239628 34054
rect 239922 33810 239950 34068
rect 240488 34054 240824 34082
rect 241040 34054 241468 34082
rect 241592 34054 241928 34082
rect 242144 34054 242480 34082
rect 242696 34054 242848 34082
rect 243248 34054 243584 34082
rect 243800 34054 244136 34082
rect 244352 34054 244688 34082
rect 244904 34054 245332 34082
rect 239922 33782 239996 33810
rect 239588 30388 239640 30394
rect 239588 30330 239640 30336
rect 239968 11354 239996 33782
rect 240796 30394 240824 34054
rect 240048 30388 240100 30394
rect 240048 30330 240100 30336
rect 240784 30388 240836 30394
rect 240784 30330 240836 30336
rect 241336 30388 241388 30394
rect 241336 30330 241388 30336
rect 239956 11348 240008 11354
rect 239956 11290 240008 11296
rect 238666 7984 238722 7993
rect 238666 7919 238722 7928
rect 240060 7857 240088 30330
rect 241348 16046 241376 30330
rect 241336 16040 241388 16046
rect 241336 15982 241388 15988
rect 240046 7848 240102 7857
rect 240046 7783 240102 7792
rect 241440 7721 241468 34054
rect 241900 30394 241928 34054
rect 242452 30462 242480 34054
rect 242164 30456 242216 30462
rect 242164 30398 242216 30404
rect 242440 30456 242492 30462
rect 242440 30398 242492 30404
rect 241888 30388 241940 30394
rect 241888 30330 241940 30336
rect 241426 7712 241482 7721
rect 241426 7647 241482 7656
rect 241704 7676 241756 7682
rect 241704 7618 241756 7624
rect 240508 6860 240560 6866
rect 240508 6802 240560 6808
rect 239312 5432 239364 5438
rect 239312 5374 239364 5380
rect 237288 3460 237340 3466
rect 237288 3402 237340 3408
rect 238114 3360 238170 3369
rect 238114 3295 238170 3304
rect 237012 3120 237064 3126
rect 237012 3062 237064 3068
rect 237024 480 237052 3062
rect 238128 480 238156 3295
rect 239324 480 239352 5374
rect 240520 480 240548 6802
rect 241716 480 241744 7618
rect 242176 6866 242204 30398
rect 242716 30388 242768 30394
rect 242716 30330 242768 30336
rect 242728 11422 242756 30330
rect 242716 11416 242768 11422
rect 242716 11358 242768 11364
rect 242820 7682 242848 34054
rect 243556 30394 243584 34054
rect 243544 30388 243596 30394
rect 243544 30330 243596 30336
rect 244108 15978 244136 34054
rect 244660 30394 244688 34054
rect 244924 30524 244976 30530
rect 244924 30466 244976 30472
rect 244188 30388 244240 30394
rect 244188 30330 244240 30336
rect 244648 30388 244700 30394
rect 244648 30330 244700 30336
rect 244096 15972 244148 15978
rect 244096 15914 244148 15920
rect 244200 11490 244228 30330
rect 244188 11484 244240 11490
rect 244188 11426 244240 11432
rect 244936 9722 244964 30466
rect 245304 26234 245332 34054
rect 245442 33810 245470 34068
rect 246008 34054 246344 34082
rect 246560 34054 246896 34082
rect 247112 34054 247448 34082
rect 247664 34054 248092 34082
rect 248216 34054 248368 34082
rect 248768 34054 249104 34082
rect 249320 34054 249748 34082
rect 249872 34054 250208 34082
rect 250516 34054 250852 34082
rect 245442 33782 245516 33810
rect 245488 30462 245516 33782
rect 245476 30456 245528 30462
rect 245476 30398 245528 30404
rect 246316 30394 246344 34054
rect 245568 30388 245620 30394
rect 245568 30330 245620 30336
rect 246304 30388 246356 30394
rect 246304 30330 246356 30336
rect 245304 26206 245516 26234
rect 245488 11558 245516 26206
rect 245476 11552 245528 11558
rect 245476 11494 245528 11500
rect 244924 9716 244976 9722
rect 244924 9658 244976 9664
rect 242808 7676 242860 7682
rect 242808 7618 242860 7624
rect 245580 7614 245608 30330
rect 246868 11626 246896 34054
rect 247420 30394 247448 34054
rect 248064 30546 248092 34054
rect 248064 30518 248276 30546
rect 246948 30388 247000 30394
rect 246948 30330 247000 30336
rect 247408 30388 247460 30394
rect 247408 30330 247460 30336
rect 248144 30388 248196 30394
rect 248144 30330 248196 30336
rect 246856 11620 246908 11626
rect 246856 11562 246908 11568
rect 245200 7608 245252 7614
rect 245200 7550 245252 7556
rect 245568 7608 245620 7614
rect 246960 7585 246988 30330
rect 248156 15910 248184 30330
rect 248144 15904 248196 15910
rect 248144 15846 248196 15852
rect 248248 14822 248276 30518
rect 248236 14816 248288 14822
rect 248236 14758 248288 14764
rect 248340 11694 248368 34054
rect 249076 31249 249104 34054
rect 249062 31240 249118 31249
rect 249062 31175 249118 31184
rect 249720 14754 249748 34054
rect 250180 30530 250208 34054
rect 250824 31822 250852 34054
rect 251008 34054 251068 34082
rect 251620 34054 251956 34082
rect 252172 34054 252508 34082
rect 252724 34054 253060 34082
rect 253276 34054 253704 34082
rect 250812 31816 250864 31822
rect 250812 31758 250864 31764
rect 251008 30818 251036 34054
rect 251088 31816 251140 31822
rect 251088 31758 251140 31764
rect 250916 30790 251036 30818
rect 250168 30524 250220 30530
rect 250168 30466 250220 30472
rect 249708 14748 249760 14754
rect 249708 14690 249760 14696
rect 250916 14618 250944 30790
rect 250996 30524 251048 30530
rect 250996 30466 251048 30472
rect 250904 14612 250956 14618
rect 250904 14554 250956 14560
rect 251008 12442 251036 30466
rect 250996 12436 251048 12442
rect 250996 12378 251048 12384
rect 248328 11688 248380 11694
rect 248328 11630 248380 11636
rect 248788 8492 248840 8498
rect 248788 8434 248840 8440
rect 245568 7550 245620 7556
rect 246946 7576 247002 7585
rect 242164 6860 242216 6866
rect 242164 6802 242216 6808
rect 244096 6520 244148 6526
rect 244096 6462 244148 6468
rect 242900 5364 242952 5370
rect 242900 5306 242952 5312
rect 242912 480 242940 5306
rect 244108 480 244136 6462
rect 245212 480 245240 7550
rect 246946 7511 247002 7520
rect 247592 6452 247644 6458
rect 247592 6394 247644 6400
rect 246396 5296 246448 5302
rect 246396 5238 246448 5244
rect 246408 480 246436 5238
rect 247604 480 247632 6394
rect 248800 480 248828 8434
rect 249984 5228 250036 5234
rect 249984 5170 250036 5176
rect 249996 480 250024 5170
rect 251100 3505 251128 31758
rect 251928 30530 251956 34054
rect 252480 31113 252508 34054
rect 252466 31104 252522 31113
rect 252466 31039 252522 31048
rect 253032 30530 253060 34054
rect 251916 30524 251968 30530
rect 251916 30466 251968 30472
rect 252468 30524 252520 30530
rect 252468 30466 252520 30472
rect 253020 30524 253072 30530
rect 253020 30466 253072 30472
rect 253572 30524 253624 30530
rect 253572 30466 253624 30472
rect 252480 12374 252508 30466
rect 253584 26234 253612 30466
rect 253676 30138 253704 34054
rect 253814 33810 253842 34068
rect 254380 34054 254716 34082
rect 254932 34054 255268 34082
rect 255484 34054 255820 34082
rect 256036 34054 256464 34082
rect 253814 33782 253888 33810
rect 253676 30110 253796 30138
rect 253584 26206 253704 26234
rect 253676 14686 253704 26206
rect 253664 14680 253716 14686
rect 253664 14622 253716 14628
rect 252468 12368 252520 12374
rect 252468 12310 252520 12316
rect 253768 12306 253796 30110
rect 253756 12300 253808 12306
rect 253756 12242 253808 12248
rect 252376 8560 252428 8566
rect 252376 8502 252428 8508
rect 251180 6384 251232 6390
rect 251180 6326 251232 6332
rect 251086 3496 251142 3505
rect 251086 3431 251142 3440
rect 251192 480 251220 6326
rect 252388 480 252416 8502
rect 253480 5160 253532 5166
rect 253480 5102 253532 5108
rect 253492 480 253520 5102
rect 253860 3369 253888 33782
rect 254688 30530 254716 34054
rect 254676 30524 254728 30530
rect 254676 30466 254728 30472
rect 255136 30524 255188 30530
rect 255136 30466 255188 30472
rect 255148 12986 255176 30466
rect 255136 12980 255188 12986
rect 255136 12922 255188 12928
rect 255240 8498 255268 34054
rect 255792 30530 255820 34054
rect 255780 30524 255832 30530
rect 255780 30466 255832 30472
rect 256436 13054 256464 34054
rect 256574 33810 256602 34068
rect 257140 34054 257476 34082
rect 257692 34054 257936 34082
rect 258244 34054 258580 34082
rect 258796 34054 259132 34082
rect 256574 33782 256648 33810
rect 256516 30524 256568 30530
rect 256516 30466 256568 30472
rect 256424 13048 256476 13054
rect 256424 12990 256476 12996
rect 256528 12238 256556 30466
rect 256516 12232 256568 12238
rect 256516 12174 256568 12180
rect 255872 8628 255924 8634
rect 255872 8570 255924 8576
rect 255228 8492 255280 8498
rect 255228 8434 255280 8440
rect 254674 6624 254730 6633
rect 254674 6559 254730 6568
rect 253846 3360 253902 3369
rect 253846 3295 253902 3304
rect 254688 480 254716 6559
rect 255884 480 255912 8570
rect 256620 8566 256648 33782
rect 257448 30530 257476 34054
rect 257436 30524 257488 30530
rect 257436 30466 257488 30472
rect 257908 13802 257936 34054
rect 257988 30524 258040 30530
rect 257988 30466 258040 30472
rect 257896 13796 257948 13802
rect 257896 13738 257948 13744
rect 258000 12170 258028 30466
rect 258552 27334 258580 34054
rect 259104 30530 259132 34054
rect 259196 34054 259348 34082
rect 259900 34054 260236 34082
rect 260452 34054 260696 34082
rect 261096 34054 261432 34082
rect 261648 34054 261984 34082
rect 259092 30524 259144 30530
rect 259092 30466 259144 30472
rect 258540 27328 258592 27334
rect 258540 27270 258592 27276
rect 259196 13734 259224 34054
rect 260208 30530 260236 34054
rect 259276 30524 259328 30530
rect 259276 30466 259328 30472
rect 260196 30524 260248 30530
rect 260196 30466 260248 30472
rect 259184 13728 259236 13734
rect 259184 13670 259236 13676
rect 257988 12164 258040 12170
rect 257988 12106 258040 12112
rect 259288 12102 259316 30466
rect 259368 27328 259420 27334
rect 259368 27270 259420 27276
rect 259276 12096 259328 12102
rect 259276 12038 259328 12044
rect 259380 8634 259408 27270
rect 260668 12034 260696 34054
rect 261404 30530 261432 34054
rect 261956 31822 261984 34054
rect 262048 34054 262200 34082
rect 262752 34054 263088 34082
rect 263304 34054 263456 34082
rect 263856 34054 264192 34082
rect 264408 34054 264744 34082
rect 261944 31816 261996 31822
rect 261944 31758 261996 31764
rect 260748 30524 260800 30530
rect 260748 30466 260800 30472
rect 261392 30524 261444 30530
rect 261392 30466 261444 30472
rect 261944 30524 261996 30530
rect 261944 30466 261996 30472
rect 260656 12028 260708 12034
rect 260656 11970 260708 11976
rect 259460 8764 259512 8770
rect 259460 8706 259512 8712
rect 259368 8628 259420 8634
rect 259368 8570 259420 8576
rect 256608 8560 256660 8566
rect 256608 8502 256660 8508
rect 258262 6488 258318 6497
rect 258262 6423 258318 6432
rect 257068 5092 257120 5098
rect 257068 5034 257120 5040
rect 257080 480 257108 5034
rect 258276 480 258304 6423
rect 259472 480 259500 8706
rect 260760 6526 260788 30466
rect 261956 13666 261984 30466
rect 261944 13660 261996 13666
rect 261944 13602 261996 13608
rect 262048 11966 262076 34054
rect 262128 31816 262180 31822
rect 262128 31758 262180 31764
rect 262036 11960 262088 11966
rect 262036 11902 262088 11908
rect 262140 8770 262168 31758
rect 263060 30530 263088 34054
rect 263048 30524 263100 30530
rect 263048 30466 263100 30472
rect 263428 8770 263456 34054
rect 264164 30530 264192 34054
rect 264716 31822 264744 34054
rect 264808 34054 264960 34082
rect 265512 34054 265940 34082
rect 266064 34054 266308 34082
rect 266616 34054 266952 34082
rect 267168 34054 267504 34082
rect 264704 31816 264756 31822
rect 264704 31758 264756 31764
rect 263508 30524 263560 30530
rect 263508 30466 263560 30472
rect 264152 30524 264204 30530
rect 264152 30466 264204 30472
rect 264704 30524 264756 30530
rect 264704 30466 264756 30472
rect 262128 8764 262180 8770
rect 262128 8706 262180 8712
rect 263416 8764 263468 8770
rect 263416 8706 263468 8712
rect 262956 8696 263008 8702
rect 262956 8638 263008 8644
rect 260748 6520 260800 6526
rect 260748 6462 260800 6468
rect 261760 6316 261812 6322
rect 261760 6258 261812 6264
rect 260654 4992 260710 5001
rect 260654 4927 260710 4936
rect 260668 480 260696 4927
rect 261772 480 261800 6258
rect 262968 480 262996 8638
rect 263520 4690 263548 30466
rect 264716 11898 264744 30466
rect 264704 11892 264756 11898
rect 264704 11834 264756 11840
rect 264808 6458 264836 34054
rect 264888 31816 264940 31822
rect 264888 31758 264940 31764
rect 264796 6452 264848 6458
rect 264796 6394 264848 6400
rect 264900 5098 264928 31758
rect 265912 26234 265940 34054
rect 265912 26206 266216 26234
rect 266188 11830 266216 26206
rect 266176 11824 266228 11830
rect 266176 11766 266228 11772
rect 265346 6352 265402 6361
rect 265346 6287 265402 6296
rect 264888 5092 264940 5098
rect 264888 5034 264940 5040
rect 264152 5024 264204 5030
rect 264152 4966 264204 4972
rect 263508 4684 263560 4690
rect 263508 4626 263560 4632
rect 264164 480 264192 4966
rect 265360 480 265388 6287
rect 266280 5030 266308 34054
rect 266924 30530 266952 34054
rect 266912 30524 266964 30530
rect 266912 30466 266964 30472
rect 267476 11762 267504 34054
rect 267660 34054 267720 34082
rect 268272 34054 268608 34082
rect 268824 34054 268976 34082
rect 269376 34054 269712 34082
rect 269928 34054 270356 34082
rect 267556 30524 267608 30530
rect 267556 30466 267608 30472
rect 267464 11756 267516 11762
rect 267464 11698 267516 11704
rect 267568 8838 267596 30466
rect 266544 8832 266596 8838
rect 266544 8774 266596 8780
rect 267556 8832 267608 8838
rect 267556 8774 267608 8780
rect 266268 5024 266320 5030
rect 266268 4966 266320 4972
rect 266556 480 266584 8774
rect 267660 4486 267688 34054
rect 268580 30530 268608 34054
rect 268568 30524 268620 30530
rect 268568 30466 268620 30472
rect 268948 12073 268976 34054
rect 269684 30666 269712 34054
rect 269672 30660 269724 30666
rect 269672 30602 269724 30608
rect 269028 30524 269080 30530
rect 269028 30466 269080 30472
rect 270224 30524 270276 30530
rect 270224 30466 270276 30472
rect 268934 12064 268990 12073
rect 268934 11999 268990 12008
rect 269040 6390 269068 30466
rect 270236 11801 270264 30466
rect 270222 11792 270278 11801
rect 270222 11727 270278 11736
rect 270328 8906 270356 34054
rect 270420 34054 270480 34082
rect 271032 34054 271368 34082
rect 270420 30530 270448 34054
rect 270500 30660 270552 30666
rect 270500 30602 270552 30608
rect 270408 30524 270460 30530
rect 270408 30466 270460 30472
rect 270512 30410 270540 30602
rect 271340 30530 271368 34054
rect 271662 33810 271690 34068
rect 272228 34054 272564 34082
rect 272780 34054 273208 34082
rect 273332 34054 273668 34082
rect 273884 34054 274312 34082
rect 274436 34054 274588 34082
rect 274988 34054 275324 34082
rect 275540 34054 275876 34082
rect 276092 34054 276428 34082
rect 276644 34054 276980 34082
rect 271662 33782 271736 33810
rect 271328 30524 271380 30530
rect 271328 30466 271380 30472
rect 270420 30382 270540 30410
rect 270040 8900 270092 8906
rect 270040 8842 270092 8848
rect 270316 8900 270368 8906
rect 270316 8842 270368 8848
rect 269028 6384 269080 6390
rect 269028 6326 269080 6332
rect 268844 6248 268896 6254
rect 268844 6190 268896 6196
rect 267738 4856 267794 4865
rect 267738 4791 267794 4800
rect 267648 4480 267700 4486
rect 267648 4422 267700 4428
rect 267752 480 267780 4791
rect 268856 480 268884 6190
rect 270052 480 270080 8842
rect 270420 4486 270448 30382
rect 271708 6322 271736 33782
rect 272536 30530 272564 34054
rect 271788 30524 271840 30530
rect 271788 30466 271840 30472
rect 272524 30524 272576 30530
rect 272524 30466 272576 30472
rect 273076 30524 273128 30530
rect 273076 30466 273128 30472
rect 271696 6316 271748 6322
rect 271696 6258 271748 6264
rect 271800 5166 271828 30466
rect 273088 11937 273116 30466
rect 273074 11928 273130 11937
rect 273074 11863 273130 11872
rect 272430 6216 272486 6225
rect 272430 6151 272486 6160
rect 271788 5160 271840 5166
rect 271788 5102 271840 5108
rect 271236 4956 271288 4962
rect 271236 4898 271288 4904
rect 270408 4480 270460 4486
rect 270408 4422 270460 4428
rect 271248 480 271276 4898
rect 272444 480 272472 6151
rect 273180 5098 273208 34054
rect 273640 30530 273668 34054
rect 273628 30524 273680 30530
rect 273628 30466 273680 30472
rect 274284 26234 274312 34054
rect 274456 30524 274508 30530
rect 274456 30466 274508 30472
rect 274284 26206 274404 26234
rect 274376 11665 274404 26206
rect 274362 11656 274418 11665
rect 274362 11591 274418 11600
rect 274468 9654 274496 30466
rect 273628 9648 273680 9654
rect 273628 9590 273680 9596
rect 274456 9648 274508 9654
rect 274456 9590 274508 9596
rect 273168 5092 273220 5098
rect 273168 5034 273220 5040
rect 273640 480 273668 9590
rect 274560 5438 274588 34054
rect 275296 30530 275324 34054
rect 275284 30524 275336 30530
rect 275284 30466 275336 30472
rect 275848 13598 275876 34054
rect 276400 30666 276428 34054
rect 276296 30660 276348 30666
rect 276296 30602 276348 30608
rect 276388 30660 276440 30666
rect 276388 30602 276440 30608
rect 275928 30524 275980 30530
rect 275928 30466 275980 30472
rect 275836 13592 275888 13598
rect 275836 13534 275888 13540
rect 274824 13456 274876 13462
rect 274824 13398 274876 13404
rect 274548 5432 274600 5438
rect 274548 5374 274600 5380
rect 274836 480 274864 13398
rect 275940 6254 275968 30466
rect 276308 26234 276336 30602
rect 276952 30530 276980 34054
rect 277136 34054 277196 34082
rect 277748 34054 278084 34082
rect 278300 34054 278636 34082
rect 278852 34054 279188 34082
rect 279404 34054 279740 34082
rect 276940 30524 276992 30530
rect 276940 30466 276992 30472
rect 276308 26206 276704 26234
rect 276676 7002 276704 26206
rect 277136 13530 277164 34054
rect 277308 30660 277360 30666
rect 277308 30602 277360 30608
rect 277216 30524 277268 30530
rect 277216 30466 277268 30472
rect 277124 13524 277176 13530
rect 277124 13466 277176 13472
rect 277228 9586 277256 30466
rect 277124 9580 277176 9586
rect 277124 9522 277176 9528
rect 277216 9580 277268 9586
rect 277216 9522 277268 9528
rect 276020 6996 276072 7002
rect 276020 6938 276072 6944
rect 276664 6996 276716 7002
rect 276664 6938 276716 6944
rect 275928 6248 275980 6254
rect 275928 6190 275980 6196
rect 276032 480 276060 6938
rect 277136 480 277164 9522
rect 277320 5370 277348 30602
rect 278056 30530 278084 34054
rect 278044 30524 278096 30530
rect 278044 30466 278096 30472
rect 278320 13388 278372 13394
rect 278320 13330 278372 13336
rect 277308 5364 277360 5370
rect 277308 5306 277360 5312
rect 278332 480 278360 13330
rect 278608 6633 278636 34054
rect 279160 30530 279188 34054
rect 279712 30666 279740 34054
rect 279942 33810 279970 34068
rect 280508 34054 280844 34082
rect 281060 34054 281488 34082
rect 281612 34054 281948 34082
rect 282256 34054 282684 34082
rect 279942 33782 280016 33810
rect 279700 30660 279752 30666
rect 279700 30602 279752 30608
rect 278688 30524 278740 30530
rect 278688 30466 278740 30472
rect 279148 30524 279200 30530
rect 279148 30466 279200 30472
rect 279884 30524 279936 30530
rect 279884 30466 279936 30472
rect 278594 6624 278650 6633
rect 278594 6559 278650 6568
rect 278700 5506 278728 30466
rect 279896 13462 279924 30466
rect 279884 13456 279936 13462
rect 279884 13398 279936 13404
rect 279516 9512 279568 9518
rect 279516 9454 279568 9460
rect 278688 5500 278740 5506
rect 278688 5442 278740 5448
rect 279528 480 279556 9454
rect 279988 9450 280016 33782
rect 280068 30660 280120 30666
rect 280068 30602 280120 30608
rect 279976 9444 280028 9450
rect 279976 9386 280028 9392
rect 280080 5438 280108 30602
rect 280816 30530 280844 34054
rect 280804 30524 280856 30530
rect 280804 30466 280856 30472
rect 281356 30524 281408 30530
rect 281356 30466 281408 30472
rect 281368 13394 281396 30466
rect 281356 13388 281408 13394
rect 281356 13330 281408 13336
rect 280712 9512 280764 9518
rect 280712 9454 280764 9460
rect 280068 5432 280120 5438
rect 280068 5374 280120 5380
rect 280724 480 280752 9454
rect 281460 5030 281488 34054
rect 281920 30530 281948 34054
rect 281908 30524 281960 30530
rect 281908 30466 281960 30472
rect 282656 13433 282684 34054
rect 282794 33810 282822 34068
rect 283360 34054 283696 34082
rect 283912 34054 284156 34082
rect 284464 34054 284800 34082
rect 285016 34054 285352 34082
rect 282794 33782 282868 33810
rect 282736 30524 282788 30530
rect 282736 30466 282788 30472
rect 282642 13424 282698 13433
rect 282642 13359 282698 13368
rect 282748 9518 282776 30466
rect 282736 9512 282788 9518
rect 282736 9454 282788 9460
rect 282840 5370 282868 33782
rect 283668 30530 283696 34054
rect 283656 30524 283708 30530
rect 283656 30466 283708 30472
rect 284128 13297 284156 34054
rect 284772 30666 284800 34054
rect 284760 30660 284812 30666
rect 284760 30602 284812 30608
rect 285324 30530 285352 34054
rect 285416 34054 285568 34082
rect 286120 34054 286456 34082
rect 286672 34054 286916 34082
rect 287224 34054 287560 34082
rect 287776 34054 288112 34082
rect 284208 30524 284260 30530
rect 284208 30466 284260 30472
rect 285312 30524 285364 30530
rect 285312 30466 285364 30472
rect 284114 13288 284170 13297
rect 284114 13223 284170 13232
rect 284220 9450 284248 30466
rect 285416 13326 285444 34054
rect 285588 30660 285640 30666
rect 285588 30602 285640 30608
rect 285496 30524 285548 30530
rect 285496 30466 285548 30472
rect 284944 13320 284996 13326
rect 284944 13262 284996 13268
rect 285404 13320 285456 13326
rect 285404 13262 285456 13268
rect 284208 9444 284260 9450
rect 284208 9386 284260 9392
rect 283104 9308 283156 9314
rect 283104 9250 283156 9256
rect 282828 5364 282880 5370
rect 282828 5306 282880 5312
rect 281908 5228 281960 5234
rect 281908 5170 281960 5176
rect 281448 5024 281500 5030
rect 281448 4966 281500 4972
rect 281920 480 281948 5170
rect 283116 480 283144 9250
rect 284300 5296 284352 5302
rect 284300 5238 284352 5244
rect 284312 480 284340 5238
rect 284956 490 284984 13262
rect 285508 6497 285536 30466
rect 285494 6488 285550 6497
rect 285494 6423 285550 6432
rect 285600 5302 285628 30602
rect 286428 30530 286456 34054
rect 286416 30524 286468 30530
rect 286416 30466 286468 30472
rect 286600 9376 286652 9382
rect 286600 9318 286652 9324
rect 285588 5296 285640 5302
rect 285588 5238 285640 5244
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 9318
rect 286888 9314 286916 34054
rect 287532 30530 287560 34054
rect 288084 30666 288112 34054
rect 288268 34054 288328 34082
rect 288880 34054 289216 34082
rect 289432 34054 289768 34082
rect 289984 34054 290320 34082
rect 290536 34054 290964 34082
rect 288072 30660 288124 30666
rect 288072 30602 288124 30608
rect 286968 30524 287020 30530
rect 286968 30466 287020 30472
rect 287520 30524 287572 30530
rect 287520 30466 287572 30472
rect 288164 30524 288216 30530
rect 288164 30466 288216 30472
rect 286876 9308 286928 9314
rect 286876 9250 286928 9256
rect 286980 5166 287008 30466
rect 288176 13161 288204 30466
rect 288162 13152 288218 13161
rect 288162 13087 288218 13096
rect 287336 11144 287388 11150
rect 287336 11086 287388 11092
rect 286968 5160 287020 5166
rect 286968 5102 287020 5108
rect 287348 490 287376 11086
rect 288268 8945 288296 34054
rect 288348 30660 288400 30666
rect 288348 30602 288400 30608
rect 288254 8936 288310 8945
rect 288254 8871 288310 8880
rect 288360 5234 288388 30602
rect 289188 30530 289216 34054
rect 289176 30524 289228 30530
rect 289176 30466 289228 30472
rect 289636 30524 289688 30530
rect 289636 30466 289688 30472
rect 289648 13258 289676 30466
rect 288992 13252 289044 13258
rect 288992 13194 289044 13200
rect 289636 13252 289688 13258
rect 289636 13194 289688 13200
rect 288348 5228 288400 5234
rect 288348 5170 288400 5176
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 13194
rect 289740 5137 289768 34054
rect 290292 30530 290320 34054
rect 290280 30524 290332 30530
rect 290280 30466 290332 30472
rect 290936 14550 290964 34054
rect 291074 33810 291102 34068
rect 291640 34054 291976 34082
rect 292192 34054 292528 34082
rect 292836 34054 293172 34082
rect 293388 34054 293816 34082
rect 291074 33782 291148 33810
rect 291016 30524 291068 30530
rect 291016 30466 291068 30472
rect 290924 14544 290976 14550
rect 290924 14486 290976 14492
rect 290188 9240 290240 9246
rect 290188 9182 290240 9188
rect 289726 5128 289782 5137
rect 289726 5063 289782 5072
rect 290200 480 290228 9182
rect 291028 6361 291056 30466
rect 291014 6352 291070 6361
rect 291014 6287 291070 6296
rect 291120 5001 291148 33782
rect 291948 30530 291976 34054
rect 291936 30524 291988 30530
rect 291936 30466 291988 30472
rect 292396 30524 292448 30530
rect 292396 30466 292448 30472
rect 292408 14482 292436 30466
rect 292500 14793 292528 34054
rect 293144 30666 293172 34054
rect 293132 30660 293184 30666
rect 293132 30602 293184 30608
rect 293684 30524 293736 30530
rect 293684 30466 293736 30472
rect 292486 14784 292542 14793
rect 292486 14719 292542 14728
rect 292396 14476 292448 14482
rect 292396 14418 292448 14424
rect 293696 13025 293724 30466
rect 293682 13016 293738 13025
rect 293682 12951 293738 12960
rect 293788 9246 293816 34054
rect 293880 34054 293940 34082
rect 294492 34054 294828 34082
rect 295044 34054 295196 34082
rect 295596 34054 295932 34082
rect 296148 34054 296576 34082
rect 293880 30530 293908 34054
rect 293960 30660 294012 30666
rect 293960 30602 294012 30608
rect 293868 30524 293920 30530
rect 293868 30466 293920 30472
rect 293972 30410 294000 30602
rect 294800 30530 294828 34054
rect 294788 30524 294840 30530
rect 294788 30466 294840 30472
rect 293880 30382 294000 30410
rect 293776 9240 293828 9246
rect 293776 9182 293828 9188
rect 293684 9172 293736 9178
rect 293684 9114 293736 9120
rect 291660 5228 291712 5234
rect 291660 5170 291712 5176
rect 291672 5114 291700 5170
rect 291672 5098 291976 5114
rect 291672 5092 291988 5098
rect 291672 5086 291936 5092
rect 291936 5034 291988 5040
rect 291106 4992 291162 5001
rect 291106 4927 291162 4936
rect 291384 4888 291436 4894
rect 291384 4830 291436 4836
rect 291396 480 291424 4830
rect 292580 4820 292632 4826
rect 292580 4762 292632 4768
rect 292592 480 292620 4762
rect 293696 480 293724 9114
rect 293880 4826 293908 30382
rect 295168 9178 295196 34054
rect 295904 30530 295932 34054
rect 295248 30524 295300 30530
rect 295248 30466 295300 30472
rect 295892 30524 295944 30530
rect 295892 30466 295944 30472
rect 296444 30524 296496 30530
rect 296444 30466 296496 30472
rect 295156 9172 295208 9178
rect 295156 9114 295208 9120
rect 295260 5030 295288 30466
rect 296456 12510 296484 30466
rect 296548 30138 296576 34054
rect 296640 34054 296700 34082
rect 297252 34054 297680 34082
rect 297804 34054 298048 34082
rect 298356 34054 298692 34082
rect 298908 34054 299244 34082
rect 296640 30258 296668 34054
rect 296628 30252 296680 30258
rect 296628 30194 296680 30200
rect 296548 30110 296668 30138
rect 296536 30048 296588 30054
rect 296536 29990 296588 29996
rect 295616 12504 295668 12510
rect 295616 12446 295668 12452
rect 296444 12504 296496 12510
rect 296444 12446 296496 12452
rect 295248 5024 295300 5030
rect 295248 4966 295300 4972
rect 294880 4888 294932 4894
rect 294880 4830 294932 4836
rect 293868 4820 293920 4826
rect 293868 4762 293920 4768
rect 294892 480 294920 4830
rect 295628 490 295656 12446
rect 296548 6225 296576 29990
rect 296534 6216 296590 6225
rect 296534 6151 296590 6160
rect 296640 4894 296668 30110
rect 297652 26234 297680 34054
rect 297652 26206 297956 26234
rect 297928 14657 297956 26206
rect 297914 14648 297970 14657
rect 297914 14583 297970 14592
rect 297272 9036 297324 9042
rect 297272 8978 297324 8984
rect 296628 4888 296680 4894
rect 296628 4830 296680 4836
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 8978
rect 298020 4865 298048 34054
rect 298664 30530 298692 34054
rect 298652 30524 298704 30530
rect 298652 30466 298704 30472
rect 299216 14521 299244 34054
rect 299400 34054 299460 34082
rect 300012 34054 300440 34082
rect 300564 34054 300808 34082
rect 301116 34054 301452 34082
rect 301668 34054 302004 34082
rect 299296 30524 299348 30530
rect 299296 30466 299348 30472
rect 299202 14512 299258 14521
rect 299202 14447 299258 14456
rect 299308 9042 299336 30466
rect 299296 9036 299348 9042
rect 299296 8978 299348 8984
rect 299400 4962 299428 34054
rect 300412 26234 300440 34054
rect 300412 26206 300716 26234
rect 300688 13190 300716 26206
rect 299664 13184 299716 13190
rect 299664 13126 299716 13132
rect 300676 13184 300728 13190
rect 300676 13126 300728 13132
rect 298468 4956 298520 4962
rect 298468 4898 298520 4904
rect 299388 4956 299440 4962
rect 299388 4898 299440 4904
rect 298006 4856 298062 4865
rect 298006 4791 298062 4800
rect 298480 480 298508 4898
rect 299676 480 299704 13126
rect 300780 12730 300808 34054
rect 301424 30666 301452 34054
rect 301504 30728 301556 30734
rect 301504 30670 301556 30676
rect 301412 30660 301464 30666
rect 301412 30602 301464 30608
rect 300688 12702 300808 12730
rect 300688 9042 300716 12702
rect 300676 9036 300728 9042
rect 300676 8978 300728 8984
rect 300768 8968 300820 8974
rect 300768 8910 300820 8916
rect 300780 480 300808 8910
rect 301516 6866 301544 30670
rect 301976 30530 302004 34054
rect 302160 34054 302220 34082
rect 302160 31385 302188 34054
rect 302146 31376 302202 31385
rect 302146 31311 302202 31320
rect 301964 30524 302016 30530
rect 301964 30466 302016 30472
rect 302896 20670 302924 312015
rect 303068 310072 303120 310078
rect 303068 310014 303120 310020
rect 302974 309360 303030 309369
rect 302974 309295 303030 309304
rect 302988 33114 303016 309295
rect 303080 46918 303108 310014
rect 303172 86970 303200 312151
rect 303252 310208 303304 310214
rect 303252 310150 303304 310156
rect 303264 167006 303292 310150
rect 303252 167000 303304 167006
rect 303252 166942 303304 166948
rect 303356 126954 303384 312287
rect 303528 310412 303580 310418
rect 303528 310354 303580 310360
rect 303436 310276 303488 310282
rect 303436 310218 303488 310224
rect 303448 206990 303476 310218
rect 303540 273222 303568 310354
rect 304356 310344 304408 310350
rect 304356 310286 304408 310292
rect 304264 310140 304316 310146
rect 304264 310082 304316 310088
rect 303528 273216 303580 273222
rect 303528 273158 303580 273164
rect 303436 206984 303488 206990
rect 303436 206926 303488 206932
rect 303344 126948 303396 126954
rect 303344 126890 303396 126896
rect 303160 86964 303212 86970
rect 303160 86906 303212 86912
rect 304276 73166 304304 310082
rect 304368 153202 304396 310286
rect 304460 233238 304488 312423
rect 304540 310480 304592 310486
rect 304540 310422 304592 310428
rect 304552 245614 304580 310422
rect 304644 259418 304672 312938
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 304724 310004 304776 310010
rect 304724 309946 304776 309952
rect 304736 299470 304764 309946
rect 580816 309596 580868 309602
rect 580816 309538 580868 309544
rect 580632 309528 580684 309534
rect 580632 309470 580684 309476
rect 580540 309392 580592 309398
rect 580540 309334 580592 309340
rect 580356 309324 580408 309330
rect 580356 309266 580408 309272
rect 315302 309224 315358 309233
rect 315302 309159 315358 309168
rect 580264 309188 580316 309194
rect 304724 299464 304776 299470
rect 304724 299406 304776 299412
rect 304632 259412 304684 259418
rect 304632 259354 304684 259360
rect 304540 245608 304592 245614
rect 304540 245550 304592 245556
rect 304448 233232 304500 233238
rect 304448 233174 304500 233180
rect 304356 153196 304408 153202
rect 304356 153138 304408 153144
rect 304264 73160 304316 73166
rect 304264 73102 304316 73108
rect 303068 46912 303120 46918
rect 303068 46854 303120 46860
rect 302976 33108 303028 33114
rect 302976 33050 303028 33056
rect 308404 30660 308456 30666
rect 308404 30602 308456 30608
rect 304264 30524 304316 30530
rect 304264 30466 304316 30472
rect 302884 20664 302936 20670
rect 302884 20606 302936 20612
rect 304276 13122 304304 30466
rect 307760 13864 307812 13870
rect 307760 13806 307812 13812
rect 303160 13116 303212 13122
rect 303160 13058 303212 13064
rect 304264 13116 304316 13122
rect 304264 13058 304316 13064
rect 301412 6860 301464 6866
rect 301412 6802 301464 6808
rect 301504 6860 301556 6866
rect 301504 6802 301556 6808
rect 301424 490 301452 6802
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301424 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 13058
rect 306380 12640 306432 12646
rect 306380 12582 306432 12588
rect 305552 9716 305604 9722
rect 305552 9658 305604 9664
rect 304356 8356 304408 8362
rect 304356 8298 304408 8304
rect 304368 480 304396 8298
rect 305564 480 305592 9658
rect 306392 490 306420 12582
rect 307772 3126 307800 13806
rect 308416 9110 308444 30602
rect 309784 30592 309836 30598
rect 309784 30534 309836 30540
rect 309692 12572 309744 12578
rect 309692 12514 309744 12520
rect 307944 9104 307996 9110
rect 307944 9046 307996 9052
rect 308404 9104 308456 9110
rect 308404 9046 308456 9052
rect 307760 3120 307812 3126
rect 307760 3062 307812 3068
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 9046
rect 309048 3120 309100 3126
rect 309048 3062 309100 3068
rect 309060 480 309088 3062
rect 309704 490 309732 12514
rect 309796 3126 309824 30534
rect 312544 30388 312596 30394
rect 312544 30330 312596 30336
rect 311440 8424 311492 8430
rect 311440 8366 311492 8372
rect 309784 3120 309836 3126
rect 309784 3062 309836 3068
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309704 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 8366
rect 312556 2854 312584 30330
rect 313832 12708 313884 12714
rect 313832 12650 313884 12656
rect 312636 6860 312688 6866
rect 312636 6802 312688 6808
rect 312544 2848 312596 2854
rect 312544 2790 312596 2796
rect 312648 480 312676 6802
rect 313844 480 313872 12650
rect 315026 9344 315082 9353
rect 315026 9279 315082 9288
rect 315040 480 315068 9279
rect 315316 6866 315344 309159
rect 580264 309130 580316 309136
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 579988 273216 580040 273222
rect 579988 273158 580040 273164
rect 580000 272241 580028 273158
rect 579986 272232 580042 272241
rect 579986 272167 580042 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 579620 206984 579672 206990
rect 579620 206926 579672 206932
rect 579632 205737 579660 206926
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 579620 126948 579672 126954
rect 579620 126890 579672 126896
rect 579632 126041 579660 126890
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580276 59673 580304 309130
rect 580368 99521 580396 309266
rect 580448 309256 580500 309262
rect 580448 309198 580500 309204
rect 580460 112849 580488 309198
rect 580552 139369 580580 309334
rect 580644 179217 580672 309470
rect 580724 309460 580776 309466
rect 580724 309402 580776 309408
rect 580736 192545 580764 309402
rect 580828 219065 580856 309538
rect 580814 219056 580870 219065
rect 580814 218991 580870 219000
rect 580722 192536 580778 192545
rect 580722 192471 580778 192480
rect 580630 179208 580686 179217
rect 580630 179143 580686 179152
rect 580538 139360 580594 139369
rect 580538 139295 580594 139304
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580354 99512 580410 99521
rect 580354 99447 580410 99456
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 330484 31748 330536 31754
rect 330484 31690 330536 31696
rect 322202 31376 322258 31385
rect 322202 31311 322258 31320
rect 315396 30456 315448 30462
rect 315396 30398 315448 30404
rect 315304 6860 315356 6866
rect 315304 6802 315356 6808
rect 315408 2990 315436 30398
rect 316040 13932 316092 13938
rect 316040 13874 316092 13880
rect 316052 3482 316080 13874
rect 317328 12776 317380 12782
rect 317328 12718 317380 12724
rect 316052 3454 316264 3482
rect 315396 2984 315448 2990
rect 315396 2926 315448 2932
rect 316236 480 316264 3454
rect 317340 480 317368 12718
rect 318522 9208 318578 9217
rect 318522 9143 318578 9152
rect 318536 480 318564 9143
rect 322110 9072 322166 9081
rect 322110 9007 322166 9016
rect 319720 6996 319772 7002
rect 319720 6938 319772 6944
rect 319732 480 319760 6938
rect 320916 6180 320968 6186
rect 320916 6122 320968 6128
rect 320928 480 320956 6122
rect 322124 480 322152 9007
rect 322216 6186 322244 31311
rect 323582 31240 323638 31249
rect 323582 31175 323638 31184
rect 322204 6180 322256 6186
rect 322204 6122 322256 6128
rect 323596 3641 323624 31175
rect 323676 30796 323728 30802
rect 323676 30738 323728 30744
rect 323582 3632 323638 3641
rect 323582 3567 323638 3576
rect 323688 2922 323716 30738
rect 328736 14136 328788 14142
rect 328736 14078 328788 14084
rect 326344 14068 326396 14074
rect 326344 14010 326396 14016
rect 324320 14000 324372 14006
rect 324320 13942 324372 13948
rect 323308 2916 323360 2922
rect 323308 2858 323360 2864
rect 323676 2916 323728 2922
rect 323676 2858 323728 2864
rect 323320 480 323348 2858
rect 324332 2786 324360 13942
rect 324412 5568 324464 5574
rect 324412 5510 324464 5516
rect 324320 2780 324372 2786
rect 324320 2722 324372 2728
rect 324424 480 324452 5510
rect 325608 2780 325660 2786
rect 325608 2722 325660 2728
rect 325620 480 325648 2722
rect 326356 490 326384 14010
rect 328000 5636 328052 5642
rect 328000 5578 328052 5584
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 5578
rect 328748 490 328776 14078
rect 330496 3058 330524 31690
rect 358084 31680 358136 31686
rect 358084 31622 358136 31628
rect 351184 31612 351236 31618
rect 351184 31554 351236 31560
rect 348424 31544 348476 31550
rect 348424 31486 348476 31492
rect 341524 31340 341576 31346
rect 341524 31282 341576 31288
rect 337384 30932 337436 30938
rect 337384 30874 337436 30880
rect 333244 30864 333296 30870
rect 333244 30806 333296 30812
rect 332692 14272 332744 14278
rect 332692 14214 332744 14220
rect 331588 5704 331640 5710
rect 331588 5646 331640 5652
rect 330392 3052 330444 3058
rect 330392 2994 330444 3000
rect 330484 3052 330536 3058
rect 330484 2994 330536 3000
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 2994
rect 331600 480 331628 5646
rect 332704 480 332732 14214
rect 333256 3058 333284 30806
rect 337396 16574 337424 30874
rect 337396 16546 337608 16574
rect 336280 14204 336332 14210
rect 336280 14146 336332 14152
rect 335084 5772 335136 5778
rect 335084 5714 335136 5720
rect 333244 3052 333296 3058
rect 333244 2994 333296 3000
rect 333888 2916 333940 2922
rect 333888 2858 333940 2864
rect 333900 480 333928 2858
rect 335096 480 335124 5714
rect 336292 480 336320 14146
rect 337580 3194 337608 16546
rect 339500 9784 339552 9790
rect 339500 9726 339552 9732
rect 338672 5840 338724 5846
rect 338672 5782 338724 5788
rect 337476 3188 337528 3194
rect 337476 3130 337528 3136
rect 337568 3188 337620 3194
rect 337568 3130 337620 3136
rect 337488 480 337516 3130
rect 338684 480 338712 5782
rect 339512 490 339540 9726
rect 341536 2922 341564 31282
rect 344284 31000 344336 31006
rect 344284 30942 344336 30948
rect 342904 9852 342956 9858
rect 342904 9794 342956 9800
rect 342168 5908 342220 5914
rect 342168 5850 342220 5856
rect 340972 2916 341024 2922
rect 340972 2858 341024 2864
rect 341524 2916 341576 2922
rect 341524 2858 341576 2864
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 2858
rect 342180 480 342208 5850
rect 342916 490 342944 9794
rect 344296 3194 344324 30942
rect 346952 9920 347004 9926
rect 346952 9862 347004 9868
rect 345756 5976 345808 5982
rect 345756 5918 345808 5924
rect 344560 3256 344612 3262
rect 344560 3198 344612 3204
rect 344284 3188 344336 3194
rect 344284 3130 344336 3136
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3198
rect 345768 480 345796 5918
rect 346964 480 346992 9862
rect 348436 3233 348464 31486
rect 349160 9988 349212 9994
rect 349160 9930 349212 9936
rect 349172 3330 349200 9930
rect 349252 6044 349304 6050
rect 349252 5986 349304 5992
rect 349160 3324 349212 3330
rect 349160 3266 349212 3272
rect 348422 3224 348478 3233
rect 348422 3159 348478 3168
rect 348056 3052 348108 3058
rect 348056 2994 348108 3000
rect 348068 480 348096 2994
rect 349264 480 349292 5986
rect 351196 3330 351224 31554
rect 355324 31204 355376 31210
rect 355324 31146 355376 31152
rect 353576 10056 353628 10062
rect 353576 9998 353628 10004
rect 352840 6112 352892 6118
rect 352840 6054 352892 6060
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 351184 3324 351236 3330
rect 351184 3266 351236 3272
rect 351828 3324 351880 3330
rect 351828 3266 351880 3272
rect 350460 480 350488 3266
rect 351644 3256 351696 3262
rect 351840 3233 351868 3266
rect 351644 3198 351696 3204
rect 351826 3224 351882 3233
rect 351656 480 351684 3198
rect 351826 3159 351882 3168
rect 352852 480 352880 6054
rect 353588 490 353616 9998
rect 355336 2922 355364 31146
rect 357532 10124 357584 10130
rect 357532 10066 357584 10072
rect 356334 5264 356390 5273
rect 356334 5199 356390 5208
rect 355968 3392 356020 3398
rect 355888 3340 355968 3346
rect 355888 3334 356020 3340
rect 355888 3318 356008 3334
rect 355888 3262 355916 3318
rect 355876 3256 355928 3262
rect 355876 3198 355928 3204
rect 355232 2916 355284 2922
rect 355232 2858 355284 2864
rect 355324 2916 355376 2922
rect 355324 2858 355376 2864
rect 353864 598 354076 626
rect 353864 490 353892 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 462 353892 490
rect 354048 480 354076 598
rect 355244 480 355272 2858
rect 356348 480 356376 5199
rect 357544 480 357572 10066
rect 358096 3398 358124 31622
rect 376024 31476 376076 31482
rect 376024 31418 376076 31424
rect 362224 31408 362276 31414
rect 362224 31350 362276 31356
rect 362236 16574 362264 31350
rect 369124 31272 369176 31278
rect 369124 31214 369176 31220
rect 366364 31136 366416 31142
rect 366364 31078 366416 31084
rect 362236 16546 362448 16574
rect 361120 10192 361172 10198
rect 361120 10134 361172 10140
rect 359924 6792 359976 6798
rect 359924 6734 359976 6740
rect 358084 3392 358136 3398
rect 358084 3334 358136 3340
rect 358728 2916 358780 2922
rect 358728 2858 358780 2864
rect 358740 480 358768 2858
rect 359936 480 359964 6734
rect 361132 480 361160 10134
rect 362420 3058 362448 16546
rect 364616 10260 364668 10266
rect 364616 10202 364668 10208
rect 363512 6724 363564 6730
rect 363512 6666 363564 6672
rect 362316 3052 362368 3058
rect 362316 2994 362368 3000
rect 362408 3052 362460 3058
rect 362408 2994 362460 3000
rect 362328 480 362356 2994
rect 363524 480 363552 6666
rect 364628 480 364656 10202
rect 366376 4146 366404 31078
rect 369136 16574 369164 31214
rect 373264 31068 373316 31074
rect 373264 31010 373316 31016
rect 369136 16546 369532 16574
rect 367744 11008 367796 11014
rect 367744 10950 367796 10956
rect 367008 6656 367060 6662
rect 367008 6598 367060 6604
rect 365812 4140 365864 4146
rect 365812 4082 365864 4088
rect 366364 4140 366416 4146
rect 366364 4082 366416 4088
rect 365824 480 365852 4082
rect 367020 480 367048 6598
rect 367756 490 367784 10950
rect 369504 3398 369532 16546
rect 370136 12844 370188 12850
rect 370136 12786 370188 12792
rect 369492 3392 369544 3398
rect 369492 3334 369544 3340
rect 369400 3256 369452 3262
rect 369400 3198 369452 3204
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 3198
rect 370148 490 370176 12786
rect 371240 10940 371292 10946
rect 371240 10882 371292 10888
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371252 490 371280 10882
rect 372896 4072 372948 4078
rect 372896 4014 372948 4020
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 370566 -960 370678 480
rect 371252 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 4014
rect 373276 3398 373304 31010
rect 376036 16574 376064 31418
rect 382922 31104 382978 31113
rect 382922 31039 382978 31048
rect 380162 30968 380218 30977
rect 380162 30903 380218 30912
rect 376036 16546 376616 16574
rect 374092 12912 374144 12918
rect 374092 12854 374144 12860
rect 373264 3392 373316 3398
rect 373264 3334 373316 3340
rect 374104 480 374132 12854
rect 375288 10872 375340 10878
rect 375288 10814 375340 10820
rect 375300 480 375328 10814
rect 376588 4078 376616 16546
rect 377680 14340 377732 14346
rect 377680 14282 377732 14288
rect 376484 4072 376536 4078
rect 376484 4014 376536 4020
rect 376576 4072 376628 4078
rect 376576 4014 376628 4020
rect 376496 480 376524 4014
rect 377692 480 377720 14282
rect 378416 10804 378468 10810
rect 378416 10746 378468 10752
rect 378428 490 378456 10746
rect 380176 4078 380204 30903
rect 381176 14408 381228 14414
rect 381176 14350 381228 14356
rect 380164 4072 380216 4078
rect 380164 4014 380216 4020
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 3946
rect 381188 480 381216 14350
rect 382372 10736 382424 10742
rect 382372 10678 382424 10684
rect 382384 480 382412 10678
rect 382936 4010 382964 31039
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 436744 16108 436796 16114
rect 436744 16050 436796 16056
rect 420920 15156 420972 15162
rect 420920 15098 420972 15104
rect 418804 12504 418856 12510
rect 418804 12446 418856 12452
rect 407210 10704 407266 10713
rect 385960 10668 386012 10674
rect 407210 10639 407266 10648
rect 385960 10610 386012 10616
rect 384764 7064 384816 7070
rect 384764 7006 384816 7012
rect 383476 4140 383528 4146
rect 383476 4082 383528 4088
rect 382924 4004 382976 4010
rect 382924 3946 382976 3952
rect 383488 3754 383516 4082
rect 383488 3726 383608 3754
rect 383580 3330 383608 3726
rect 383476 3324 383528 3330
rect 383476 3266 383528 3272
rect 383568 3324 383620 3330
rect 383568 3266 383620 3272
rect 383488 1714 383516 3266
rect 383488 1686 383608 1714
rect 383580 480 383608 1686
rect 384776 480 384804 7006
rect 385972 480 386000 10610
rect 389456 10600 389508 10606
rect 389456 10542 389508 10548
rect 388260 7132 388312 7138
rect 388260 7074 388312 7080
rect 387156 3936 387208 3942
rect 387156 3878 387208 3884
rect 387168 480 387196 3878
rect 388272 480 388300 7074
rect 389468 480 389496 10542
rect 392584 10532 392636 10538
rect 392584 10474 392636 10480
rect 391848 7200 391900 7206
rect 391848 7142 391900 7148
rect 390652 2916 390704 2922
rect 390652 2858 390704 2864
rect 390664 480 390692 2858
rect 391860 480 391888 7142
rect 392596 490 392624 10474
rect 396080 10464 396132 10470
rect 396080 10406 396132 10412
rect 395344 7268 395396 7274
rect 395344 7210 395396 7216
rect 394240 3868 394292 3874
rect 394240 3810 394292 3816
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 3810
rect 395356 480 395384 7210
rect 396092 490 396120 10406
rect 398840 10396 398892 10402
rect 398840 10338 398892 10344
rect 398852 3806 398880 10338
rect 403624 10328 403676 10334
rect 403624 10270 403676 10276
rect 402520 7404 402572 7410
rect 402520 7346 402572 7352
rect 398932 7336 398984 7342
rect 398932 7278 398984 7284
rect 398840 3800 398892 3806
rect 398840 3742 398892 3748
rect 397736 3052 397788 3058
rect 397736 2994 397788 3000
rect 396368 598 396580 626
rect 396368 490 396396 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 2994
rect 398944 480 398972 7278
rect 401324 3868 401376 3874
rect 401324 3810 401376 3816
rect 400128 3800 400180 3806
rect 400128 3742 400180 3748
rect 400140 480 400168 3742
rect 401336 480 401364 3810
rect 402532 480 402560 7346
rect 403636 480 403664 10270
rect 406016 7472 406068 7478
rect 406016 7414 406068 7420
rect 404820 3188 404872 3194
rect 404820 3130 404872 3136
rect 404832 480 404860 3130
rect 406028 480 406056 7414
rect 407224 480 407252 10639
rect 410798 10568 410854 10577
rect 410798 10503 410854 10512
rect 409604 7540 409656 7546
rect 409604 7482 409656 7488
rect 408408 3732 408460 3738
rect 408408 3674 408460 3680
rect 408420 480 408448 3674
rect 409616 480 409644 7482
rect 410812 480 410840 10503
rect 414294 10432 414350 10441
rect 414294 10367 414350 10376
rect 413100 8288 413152 8294
rect 413100 8230 413152 8236
rect 411904 3256 411956 3262
rect 411904 3198 411956 3204
rect 411916 480 411944 3198
rect 413112 480 413140 8230
rect 414308 480 414336 10367
rect 417422 10296 417478 10305
rect 417422 10231 417478 10240
rect 416688 8220 416740 8226
rect 416688 8162 416740 8168
rect 415492 3664 415544 3670
rect 415492 3606 415544 3612
rect 415504 480 415532 3606
rect 416700 480 416728 8162
rect 417436 490 417464 10231
rect 418816 3670 418844 12446
rect 420184 8152 420236 8158
rect 420184 8094 420236 8100
rect 418804 3664 418856 3670
rect 418804 3606 418856 3612
rect 418988 3324 419040 3330
rect 418988 3266 419040 3272
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 419000 480 419028 3266
rect 420196 480 420224 8094
rect 420932 490 420960 15098
rect 423680 15088 423732 15094
rect 423680 15030 423732 15036
rect 422576 3596 422628 3602
rect 422576 3538 422628 3544
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 3538
rect 423692 3534 423720 15030
rect 428464 15020 428516 15026
rect 428464 14962 428516 14968
rect 427268 8084 427320 8090
rect 427268 8026 427320 8032
rect 423772 8016 423824 8022
rect 423772 7958 423824 7964
rect 423680 3528 423732 3534
rect 423680 3470 423732 3476
rect 423784 480 423812 7958
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 424980 480 425008 3470
rect 426164 3392 426216 3398
rect 426164 3334 426216 3340
rect 426176 480 426204 3334
rect 427280 480 427308 8026
rect 428476 480 428504 14962
rect 432052 14952 432104 14958
rect 432052 14894 432104 14900
rect 430856 7948 430908 7954
rect 430856 7890 430908 7896
rect 429660 3596 429712 3602
rect 429660 3538 429712 3544
rect 429672 480 429700 3538
rect 430868 480 430896 7890
rect 432064 480 432092 14894
rect 435088 14884 435140 14890
rect 435088 14826 435140 14832
rect 434444 7880 434496 7886
rect 434444 7822 434496 7828
rect 433248 4140 433300 4146
rect 433248 4082 433300 4088
rect 433260 480 433288 4082
rect 434456 480 434484 7822
rect 435100 490 435128 14826
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 16050
rect 450912 16040 450964 16046
rect 450912 15982 450964 15988
rect 448520 11348 448572 11354
rect 448520 11290 448572 11296
rect 445760 11280 445812 11286
rect 445760 11222 445812 11228
rect 439136 11212 439188 11218
rect 439136 11154 439188 11160
rect 437940 7812 437992 7818
rect 437940 7754 437992 7760
rect 437952 480 437980 7754
rect 439148 480 439176 11154
rect 445022 7984 445078 7993
rect 445022 7919 445078 7928
rect 441528 7744 441580 7750
rect 441528 7686 441580 7692
rect 440332 2848 440384 2854
rect 440332 2790 440384 2796
rect 440344 480 440372 2790
rect 441540 480 441568 7686
rect 442632 6588 442684 6594
rect 442632 6530 442684 6536
rect 442644 480 442672 6530
rect 443828 3460 443880 3466
rect 443828 3402 443880 3408
rect 443840 480 443868 3402
rect 445036 480 445064 7919
rect 445772 490 445800 11222
rect 447416 4072 447468 4078
rect 447416 4014 447468 4020
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 4014
rect 448532 3534 448560 11290
rect 448610 7848 448666 7857
rect 448610 7783 448666 7792
rect 448520 3528 448572 3534
rect 448520 3470 448572 3476
rect 448624 480 448652 7783
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 449820 480 449848 3470
rect 450924 480 450952 15982
rect 456800 15972 456852 15978
rect 456800 15914 456852 15920
rect 453304 11416 453356 11422
rect 453304 11358 453356 11364
rect 452106 7712 452162 7721
rect 452106 7647 452162 7656
rect 452120 480 452148 7647
rect 453316 480 453344 11358
rect 455696 7676 455748 7682
rect 455696 7618 455748 7624
rect 454500 2984 454552 2990
rect 454500 2926 454552 2932
rect 454512 480 454540 2926
rect 455708 480 455736 7618
rect 456812 3534 456840 15914
rect 465172 15904 465224 15910
rect 465172 15846 465224 15852
rect 463976 11620 464028 11626
rect 463976 11562 464028 11568
rect 459928 11552 459980 11558
rect 459928 11494 459980 11500
rect 456892 11484 456944 11490
rect 456892 11426 456944 11432
rect 456800 3528 456852 3534
rect 456800 3470 456852 3476
rect 456904 480 456932 11426
rect 459192 7608 459244 7614
rect 459192 7550 459244 7556
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 458100 480 458128 3470
rect 459204 480 459232 7550
rect 459940 490 459968 11494
rect 462778 7576 462834 7585
rect 462778 7511 462834 7520
rect 461584 3120 461636 3126
rect 461584 3062 461636 3068
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3062
rect 462792 480 462820 7511
rect 463988 480 464016 11562
rect 465184 480 465212 15846
rect 465816 14816 465868 14822
rect 465816 14758 465868 14764
rect 560390 14784 560446 14793
rect 465828 490 465856 14758
rect 469864 14748 469916 14754
rect 560390 14719 560446 14728
rect 469864 14690 469916 14696
rect 467472 11688 467524 11694
rect 467472 11630 467524 11636
rect 466104 598 466316 626
rect 466104 490 466132 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 462 466132 490
rect 466288 480 466316 598
rect 467484 480 467512 11630
rect 468666 3632 468722 3641
rect 468666 3567 468722 3576
rect 468680 480 468708 3567
rect 469876 480 469904 14690
rect 476488 14680 476540 14686
rect 476488 14622 476540 14628
rect 473452 14612 473504 14618
rect 473452 14554 473504 14560
rect 470600 12436 470652 12442
rect 470600 12378 470652 12384
rect 470612 490 470640 12378
rect 472254 3496 472310 3505
rect 472254 3431 472310 3440
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 3431
rect 473464 480 473492 14554
rect 474096 12368 474148 12374
rect 474096 12310 474148 12316
rect 474108 490 474136 12310
rect 475752 4004 475804 4010
rect 475752 3946 475804 3952
rect 474384 598 474596 626
rect 474384 490 474412 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 462 474412 490
rect 474568 480 474596 598
rect 475764 480 475792 3946
rect 476500 490 476528 14622
rect 556896 14544 556948 14550
rect 556896 14486 556948 14492
rect 487160 13796 487212 13802
rect 487160 13738 487212 13744
rect 484032 13048 484084 13054
rect 484032 12990 484084 12996
rect 480536 12980 480588 12986
rect 480536 12922 480588 12928
rect 478144 12300 478196 12306
rect 478144 12242 478196 12248
rect 476776 598 476988 626
rect 476776 490 476804 598
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 462 476804 490
rect 476960 480 476988 598
rect 478156 480 478184 12242
rect 479338 3360 479394 3369
rect 479338 3295 479394 3304
rect 479352 480 479380 3295
rect 480548 480 480576 12922
rect 482376 12232 482428 12238
rect 482376 12174 482428 12180
rect 481732 8492 481784 8498
rect 481732 8434 481784 8440
rect 481744 480 481772 8434
rect 482388 490 482416 12174
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 12990
rect 486424 12164 486476 12170
rect 486424 12106 486476 12112
rect 485228 8560 485280 8566
rect 485228 8502 485280 8508
rect 485240 480 485268 8502
rect 486436 480 486464 12106
rect 487172 490 487200 13738
rect 489920 13728 489972 13734
rect 489920 13670 489972 13676
rect 488816 8628 488868 8634
rect 488816 8570 488868 8576
rect 487448 598 487660 626
rect 487448 490 487476 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 462 487476 490
rect 487632 480 487660 598
rect 488828 480 488856 8570
rect 489932 3602 489960 13670
rect 494704 13660 494756 13666
rect 494704 13602 494756 13608
rect 490012 12096 490064 12102
rect 490012 12038 490064 12044
rect 489920 3596 489972 3602
rect 489920 3538 489972 3544
rect 490024 3482 490052 12038
rect 493048 12028 493100 12034
rect 493048 11970 493100 11976
rect 492312 6520 492364 6526
rect 492312 6462 492364 6468
rect 491116 3596 491168 3602
rect 491116 3538 491168 3544
rect 489932 3454 490052 3482
rect 489932 480 489960 3454
rect 491128 480 491156 3538
rect 492324 480 492352 6462
rect 493060 490 493088 11970
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 13602
rect 525432 13592 525484 13598
rect 525432 13534 525484 13540
rect 511262 12064 511318 12073
rect 511262 11999 511318 12008
rect 497096 11960 497148 11966
rect 497096 11902 497148 11908
rect 495900 8696 495952 8702
rect 495900 8638 495952 8644
rect 495912 480 495940 8638
rect 497108 480 497136 11902
rect 500592 11892 500644 11898
rect 500592 11834 500644 11840
rect 499396 8764 499448 8770
rect 499396 8706 499448 8712
rect 498200 4208 498252 4214
rect 498200 4150 498252 4156
rect 498212 480 498240 4150
rect 499408 480 499436 8706
rect 500604 480 500632 11834
rect 503720 11824 503772 11830
rect 503720 11766 503772 11772
rect 502984 6452 503036 6458
rect 502984 6394 503036 6400
rect 501788 4276 501840 4282
rect 501788 4218 501840 4224
rect 501800 480 501828 4218
rect 502996 480 503024 6394
rect 503732 490 503760 11766
rect 507216 11756 507268 11762
rect 507216 11698 507268 11704
rect 506480 8832 506532 8838
rect 506480 8774 506532 8780
rect 505376 4344 505428 4350
rect 505376 4286 505428 4292
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 4286
rect 506492 480 506520 8774
rect 507228 490 507256 11698
rect 510068 6384 510120 6390
rect 510068 6326 510120 6332
rect 508872 4412 508924 4418
rect 508872 4354 508924 4360
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 4354
rect 510080 480 510108 6326
rect 511276 480 511304 11999
rect 517886 11928 517942 11937
rect 517886 11863 517942 11872
rect 514758 11792 514814 11801
rect 514758 11727 514814 11736
rect 513564 8900 513616 8906
rect 513564 8842 513616 8848
rect 512460 4480 512512 4486
rect 512460 4422 512512 4428
rect 512472 480 512500 4422
rect 513576 480 513604 8842
rect 514772 480 514800 11727
rect 517152 6316 517204 6322
rect 517152 6258 517204 6264
rect 515956 4548 516008 4554
rect 515956 4490 516008 4496
rect 515968 480 515996 4490
rect 517164 480 517192 6258
rect 517900 490 517928 11863
rect 521842 11656 521898 11665
rect 521842 11591 521898 11600
rect 520740 9648 520792 9654
rect 520740 9590 520792 9596
rect 519544 4616 519596 4622
rect 519544 4558 519596 4564
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 4558
rect 520752 480 520780 9590
rect 521856 480 521884 11591
rect 524236 6248 524288 6254
rect 524236 6190 524288 6196
rect 523040 4752 523092 4758
rect 523040 4694 523092 4700
rect 523052 480 523080 4694
rect 524248 480 524276 6190
rect 525444 480 525472 13534
rect 528560 13524 528612 13530
rect 528560 13466 528612 13472
rect 527824 9580 527876 9586
rect 527824 9522 527876 9528
rect 526628 4684 526680 4690
rect 526628 4626 526680 4632
rect 526640 480 526668 4626
rect 527836 480 527864 9522
rect 528572 490 528600 13466
rect 532056 13456 532108 13462
rect 532056 13398 532108 13404
rect 539598 13424 539654 13433
rect 531318 6624 531374 6633
rect 531318 6559 531374 6568
rect 530124 5500 530176 5506
rect 530124 5442 530176 5448
rect 528848 598 529060 626
rect 528848 490 528876 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 5442
rect 531332 480 531360 6559
rect 532068 490 532096 13398
rect 536104 13388 536156 13394
rect 539598 13359 539654 13368
rect 536104 13330 536156 13336
rect 534908 9512 534960 9518
rect 534908 9454 534960 9460
rect 533712 5432 533764 5438
rect 533712 5374 533764 5380
rect 532344 598 532556 626
rect 532344 490 532372 598
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 462 532372 490
rect 532528 480 532556 598
rect 533724 480 533752 5374
rect 534920 480 534948 9454
rect 536116 480 536144 13330
rect 538404 9444 538456 9450
rect 538404 9386 538456 9392
rect 537208 5364 537260 5370
rect 537208 5306 537260 5312
rect 537220 480 537248 5306
rect 538416 480 538444 9386
rect 539612 480 539640 13359
rect 546684 13320 546736 13326
rect 542726 13288 542782 13297
rect 546684 13262 546736 13268
rect 542726 13223 542782 13232
rect 541992 9376 542044 9382
rect 541992 9318 542044 9324
rect 540796 5296 540848 5302
rect 540796 5238 540848 5244
rect 540808 480 540836 5238
rect 542004 480 542032 9318
rect 542740 490 542768 13223
rect 545486 6488 545542 6497
rect 545486 6423 545542 6432
rect 544384 5228 544436 5234
rect 544384 5170 544436 5176
rect 543016 598 543228 626
rect 543016 490 543044 598
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 5170
rect 545500 480 545528 6423
rect 546696 480 546724 13262
rect 553768 13252 553820 13258
rect 553768 13194 553820 13200
rect 550270 13152 550326 13161
rect 550270 13087 550326 13096
rect 549076 9308 549128 9314
rect 549076 9250 549128 9256
rect 547880 5160 547932 5166
rect 547880 5102 547932 5108
rect 547892 480 547920 5102
rect 549088 480 549116 9250
rect 550284 480 550312 13087
rect 552662 8936 552718 8945
rect 552662 8871 552718 8880
rect 551468 5092 551520 5098
rect 551468 5034 551520 5040
rect 551480 480 551508 5034
rect 552676 480 552704 8871
rect 553780 480 553808 13194
rect 556158 6352 556214 6361
rect 556158 6287 556214 6296
rect 554962 5128 555018 5137
rect 554962 5063 555018 5072
rect 554976 480 555004 5063
rect 556172 480 556200 6287
rect 556908 490 556936 14486
rect 559288 14476 559340 14482
rect 559288 14418 559340 14424
rect 558550 4992 558606 5001
rect 558550 4927 558606 4936
rect 557184 598 557396 626
rect 557184 490 557212 598
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 462 557212 490
rect 557368 480 557396 598
rect 558564 480 558592 4927
rect 559300 490 559328 14418
rect 559576 598 559788 626
rect 559576 490 559604 598
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 462 559604 490
rect 559760 480 559788 598
rect 560404 490 560432 14719
rect 571522 14648 571578 14657
rect 571522 14583 571578 14592
rect 564438 13016 564494 13025
rect 564438 12951 564494 12960
rect 563244 9240 563296 9246
rect 563244 9182 563296 9188
rect 562048 5024 562100 5030
rect 562048 4966 562100 4972
rect 560680 598 560892 626
rect 560680 490 560708 598
rect 559718 -960 559830 480
rect 560404 462 560708 490
rect 560864 480 560892 598
rect 562060 480 562088 4966
rect 563256 480 563284 9182
rect 564452 480 564480 12951
rect 566832 9172 566884 9178
rect 566832 9114 566884 9120
rect 565636 4956 565688 4962
rect 565636 4898 565688 4904
rect 565648 480 565676 4898
rect 566844 480 566872 9114
rect 570326 6216 570382 6225
rect 570326 6151 570382 6160
rect 569132 4888 569184 4894
rect 569132 4830 569184 4836
rect 568028 3664 568080 3670
rect 568028 3606 568080 3612
rect 568040 480 568068 3606
rect 569144 480 569172 4830
rect 570340 480 570368 6151
rect 571536 480 571564 14583
rect 575110 14512 575166 14521
rect 575110 14447 575166 14456
rect 573916 9036 573968 9042
rect 573916 8978 573968 8984
rect 572718 4856 572774 4865
rect 572718 4791 572774 4800
rect 572732 480 572760 4791
rect 573928 480 573956 8978
rect 575124 480 575152 14447
rect 576952 13184 577004 13190
rect 576952 13126 577004 13132
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 576320 480 576348 4762
rect 576964 490 576992 13126
rect 581736 13116 581788 13122
rect 581736 13058 581788 13064
rect 581000 9104 581052 9110
rect 581000 9046 581052 9052
rect 578608 8968 578660 8974
rect 578608 8910 578660 8916
rect 577240 598 577452 626
rect 577240 490 577268 598
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 462 577268 490
rect 577424 480 577452 598
rect 578620 480 578648 8910
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 9046
rect 581748 490 581776 13058
rect 583392 3120 583444 3126
rect 583392 3062 583444 3068
rect 582024 598 582236 626
rect 582024 490 582052 598
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 462 582052 490
rect 582208 480 582236 598
rect 583404 480 583432 3062
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3146 593000 3202 593056
rect 3330 553832 3386 553888
rect 3330 540776 3386 540832
rect 3330 527856 3386 527912
rect 3330 501744 3386 501800
rect 3146 488688 3202 488744
rect 3054 475632 3110 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 3330 436600 3386 436656
rect 3146 423544 3202 423600
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3330 345344 3386 345400
rect 3698 644272 3754 644328
rect 3514 632032 3570 632088
rect 3790 619112 3846 619168
rect 3698 566888 3754 566944
rect 3606 514800 3662 514856
rect 3882 358400 3938 358456
rect 3606 319232 3662 319288
rect 2962 306212 2964 306232
rect 2964 306212 3016 306232
rect 3016 306212 3018 306232
rect 2962 306176 3018 306212
rect 2778 293120 2834 293176
rect 2778 267180 2780 267200
rect 2780 267180 2832 267200
rect 2832 267180 2834 267200
rect 2778 267144 2834 267180
rect 3514 311888 3570 311944
rect 3330 254088 3386 254144
rect 2778 214956 2780 214976
rect 2780 214956 2832 214976
rect 2832 214956 2834 214976
rect 2778 214920 2834 214956
rect 2778 162832 2834 162888
rect 2778 123664 2834 123720
rect 2778 110608 2834 110664
rect 2778 97552 2834 97608
rect 2778 84632 2834 84688
rect 2778 71612 2780 71632
rect 2780 71612 2832 71632
rect 2832 71612 2834 71632
rect 2778 71576 2834 71612
rect 3146 45500 3148 45520
rect 3148 45500 3200 45520
rect 3200 45500 3202 45520
rect 3146 45464 3202 45500
rect 2778 32408 2834 32464
rect 4066 241032 4122 241088
rect 3974 201864 4030 201920
rect 3882 188808 3938 188864
rect 3790 149776 3846 149832
rect 3698 136720 3754 136776
rect 40130 650120 40186 650176
rect 104714 645360 104770 645416
rect 98642 644292 98698 644328
rect 98642 644272 98644 644292
rect 98644 644272 98696 644292
rect 98696 644272 98698 644292
rect 104254 644292 104310 644328
rect 104254 644272 104256 644292
rect 104256 644272 104308 644292
rect 104308 644272 104310 644292
rect 133878 643592 133934 643648
rect 40130 625640 40186 625696
rect 40038 623464 40094 623520
rect 40038 582120 40094 582176
rect 40222 606736 40278 606792
rect 114466 606056 114522 606112
rect 118606 590688 118662 590744
rect 3606 58520 3662 58576
rect 68006 312432 68062 312488
rect 50986 312296 51042 312352
rect 43994 312160 44050 312216
rect 34334 312024 34390 312080
rect 121366 576816 121422 576872
rect 153106 643864 153162 643920
rect 167458 590688 167514 590744
rect 167458 580216 167514 580272
rect 167458 576816 167514 576872
rect 192390 645360 192446 645416
rect 192758 645360 192814 645416
rect 192206 644272 192262 644328
rect 189722 644000 189778 644056
rect 192758 644000 192814 644056
rect 189722 643728 189778 643784
rect 196898 644272 196954 644328
rect 196530 644000 196586 644056
rect 192206 643592 192262 643648
rect 192758 643592 192814 643648
rect 196622 643612 196678 643648
rect 196622 643592 196624 643612
rect 196624 643592 196676 643612
rect 196676 643592 196678 643612
rect 192206 643320 192262 643376
rect 190918 642932 190974 642968
rect 190918 642912 190920 642932
rect 190920 642912 190972 642932
rect 190972 642912 190974 642932
rect 192206 642132 192208 642152
rect 192208 642132 192260 642152
rect 192260 642132 192262 642152
rect 192206 642096 192262 642132
rect 300766 665216 300822 665272
rect 202694 645396 202696 645416
rect 202696 645396 202748 645416
rect 202748 645396 202750 645416
rect 202694 645360 202750 645396
rect 201774 644816 201830 644872
rect 199014 644272 199070 644328
rect 199290 644272 199346 644328
rect 198094 643592 198150 643648
rect 199290 643592 199346 643648
rect 199658 643592 199714 643648
rect 202510 643728 202566 643784
rect 202786 643728 202842 643784
rect 202234 643592 202290 643648
rect 208398 643592 208454 643648
rect 202234 643184 202290 643240
rect 206558 643184 206614 643240
rect 236182 644292 236238 644328
rect 236182 644272 236184 644292
rect 236184 644272 236236 644292
rect 236236 644272 236238 644292
rect 240690 644292 240746 644328
rect 240690 644272 240692 644292
rect 240692 644272 240744 644292
rect 240744 644272 240746 644292
rect 236182 642268 236184 642288
rect 236184 642268 236236 642288
rect 236236 642268 236238 642288
rect 236182 642232 236238 642268
rect 241610 642268 241612 642288
rect 241612 642268 241664 642288
rect 241664 642268 241666 642288
rect 241610 642232 241666 642268
rect 230478 639920 230534 639976
rect 230478 639648 230534 639704
rect 224866 639548 224868 639568
rect 224868 639548 224920 639568
rect 224920 639548 224922 639568
rect 224866 639512 224922 639548
rect 463330 688644 463332 688664
rect 463332 688644 463384 688664
rect 463384 688644 463386 688664
rect 463330 688608 463386 688644
rect 465538 688608 465594 688664
rect 459558 640464 459614 640520
rect 468666 640464 468722 640520
rect 469034 640464 469090 640520
rect 471794 640464 471850 640520
rect 404266 628088 404322 628144
rect 391846 559408 391902 559464
rect 391386 543496 391442 543552
rect 427818 551520 427874 551576
rect 580262 697176 580318 697232
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 579618 484608 579674 484664
rect 579986 471416 580042 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 579618 418240 579674 418296
rect 580170 404912 580226 404968
rect 579618 378392 579674 378448
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 579986 325216 580042 325272
rect 580538 683848 580594 683904
rect 580354 670656 580410 670712
rect 580446 644000 580502 644056
rect 580538 630808 580594 630864
rect 580630 617480 580686 617536
rect 580722 564304 580778 564360
rect 304446 312432 304502 312488
rect 303342 312296 303398 312352
rect 303158 312160 303214 312216
rect 302882 312024 302938 312080
rect 300950 311888 301006 311944
rect 29550 309984 29606 310040
rect 31758 309984 31814 310040
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 79966 3576 80022 3632
rect 84014 3440 84070 3496
rect 84106 3304 84162 3360
rect 110510 3576 110566 3632
rect 117594 3440 117650 3496
rect 118790 3304 118846 3360
rect 131026 3712 131082 3768
rect 133786 3576 133842 3632
rect 135166 3440 135222 3496
rect 139306 5072 139362 5128
rect 140686 3304 140742 3360
rect 148966 6568 149022 6624
rect 150254 6432 150310 6488
rect 153014 6296 153070 6352
rect 151726 4936 151782 4992
rect 154486 4800 154542 4856
rect 157246 6160 157302 6216
rect 176566 9288 176622 9344
rect 179234 9152 179290 9208
rect 180706 9016 180762 9072
rect 195886 5208 195942 5264
rect 216862 3712 216918 3768
rect 220634 10648 220690 10704
rect 222014 10512 222070 10568
rect 223394 10376 223450 10432
rect 224682 10240 224738 10296
rect 223946 3576 224002 3632
rect 227534 3440 227590 3496
rect 235814 5072 235870 5128
rect 238758 30912 238814 30968
rect 238666 7928 238722 7984
rect 240046 7792 240102 7848
rect 241426 7656 241482 7712
rect 238114 3304 238170 3360
rect 249062 31184 249118 31240
rect 246946 7520 247002 7576
rect 252466 31048 252522 31104
rect 251086 3440 251142 3496
rect 254674 6568 254730 6624
rect 253846 3304 253902 3360
rect 258262 6432 258318 6488
rect 260654 4936 260710 4992
rect 265346 6296 265402 6352
rect 268934 12008 268990 12064
rect 270222 11736 270278 11792
rect 267738 4800 267794 4856
rect 273074 11872 273130 11928
rect 272430 6160 272486 6216
rect 274362 11600 274418 11656
rect 278594 6568 278650 6624
rect 282642 13368 282698 13424
rect 284114 13232 284170 13288
rect 285494 6432 285550 6488
rect 288162 13096 288218 13152
rect 288254 8880 288310 8936
rect 289726 5072 289782 5128
rect 291014 6296 291070 6352
rect 292486 14728 292542 14784
rect 293682 12960 293738 13016
rect 291106 4936 291162 4992
rect 296534 6160 296590 6216
rect 297914 14592 297970 14648
rect 299202 14456 299258 14512
rect 298006 4800 298062 4856
rect 302146 31320 302202 31376
rect 302974 309304 303030 309360
rect 580170 312024 580226 312080
rect 315302 309168 315358 309224
rect 315026 9288 315082 9344
rect 580170 298696 580226 298752
rect 579986 272176 580042 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 579618 205672 579674 205728
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 579618 125976 579674 126032
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580814 219000 580870 219056
rect 580722 192480 580778 192536
rect 580630 179152 580686 179208
rect 580538 139304 580594 139360
rect 580446 112784 580502 112840
rect 580354 99456 580410 99512
rect 580262 59608 580318 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 322202 31320 322258 31376
rect 318522 9152 318578 9208
rect 322110 9016 322166 9072
rect 323582 31184 323638 31240
rect 323582 3576 323638 3632
rect 348422 3168 348478 3224
rect 351826 3168 351882 3224
rect 356334 5208 356390 5264
rect 382922 31048 382978 31104
rect 380162 30912 380218 30968
rect 579986 19760 580042 19816
rect 407210 10648 407266 10704
rect 410798 10512 410854 10568
rect 414294 10376 414350 10432
rect 417422 10240 417478 10296
rect 445022 7928 445078 7984
rect 448610 7792 448666 7848
rect 452106 7656 452162 7712
rect 462778 7520 462834 7576
rect 560390 14728 560446 14784
rect 468666 3576 468722 3632
rect 472254 3440 472310 3496
rect 479338 3304 479394 3360
rect 511262 12008 511318 12064
rect 517886 11872 517942 11928
rect 514758 11736 514814 11792
rect 521842 11600 521898 11656
rect 531318 6568 531374 6624
rect 539598 13368 539654 13424
rect 542726 13232 542782 13288
rect 545486 6432 545542 6488
rect 550270 13096 550326 13152
rect 552662 8880 552718 8936
rect 556158 6296 556214 6352
rect 554962 5072 555018 5128
rect 558550 4936 558606 4992
rect 571522 14592 571578 14648
rect 564438 12960 564494 13016
rect 570326 6160 570382 6216
rect 575110 14456 575166 14512
rect 572718 4800 572774 4856
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect 463325 688666 463391 688669
rect 465533 688666 465599 688669
rect 463325 688664 465599 688666
rect 463325 688608 463330 688664
rect 463386 688608 465538 688664
rect 465594 688608 465599 688664
rect 463325 688606 465599 688608
rect 463325 688603 463391 688606
rect 465533 688603 465599 688606
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580533 683906 580599 683909
rect 583520 683906 584960 683996
rect 580533 683904 584960 683906
rect 580533 683848 580538 683904
rect 580594 683848 584960 683904
rect 580533 683846 584960 683848
rect 580533 683843 580599 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580349 670714 580415 670717
rect 583520 670714 584960 670804
rect 580349 670712 584960 670714
rect 580349 670656 580354 670712
rect 580410 670656 584960 670712
rect 580349 670654 584960 670656
rect 580349 670651 580415 670654
rect 583520 670564 584960 670654
rect 300761 665274 300827 665277
rect 300761 665272 528570 665274
rect 300761 665216 300766 665272
rect 300822 665216 528570 665272
rect 300761 665214 528570 665216
rect 300761 665211 300827 665214
rect 528510 664972 528570 665214
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect 40174 650181 40234 650284
rect 40125 650176 40234 650181
rect 40125 650120 40130 650176
rect 40186 650120 40234 650176
rect 40125 650118 40234 650120
rect 40125 650115 40191 650118
rect 104709 645418 104775 645421
rect 192385 645418 192451 645421
rect 104709 645416 192451 645418
rect 104709 645360 104714 645416
rect 104770 645360 192390 645416
rect 192446 645360 192451 645416
rect 104709 645358 192451 645360
rect 104709 645355 104775 645358
rect 192385 645355 192451 645358
rect 192753 645418 192819 645421
rect 202689 645418 202755 645421
rect 192753 645416 202755 645418
rect 192753 645360 192758 645416
rect 192814 645360 202694 645416
rect 202750 645360 202755 645416
rect 192753 645358 202755 645360
rect 192753 645355 192819 645358
rect -960 644996 480 645236
rect 201726 644877 201786 645358
rect 202689 645355 202755 645358
rect 201726 644872 201835 644877
rect 201726 644816 201774 644872
rect 201830 644816 201835 644872
rect 201726 644814 201835 644816
rect 201769 644811 201835 644814
rect 128310 644542 133890 644602
rect 3693 644330 3759 644333
rect 98637 644330 98703 644333
rect 3693 644328 98703 644330
rect 3693 644272 3698 644328
rect 3754 644272 98642 644328
rect 98698 644272 98703 644328
rect 3693 644270 98703 644272
rect 3693 644267 3759 644270
rect 98637 644267 98703 644270
rect 104249 644330 104315 644333
rect 128310 644330 128370 644542
rect 104249 644328 128370 644330
rect 104249 644272 104254 644328
rect 104310 644272 128370 644328
rect 104249 644270 128370 644272
rect 133830 644330 133890 644542
rect 192201 644330 192267 644333
rect 133830 644328 192267 644330
rect 133830 644272 192206 644328
rect 192262 644272 192267 644328
rect 133830 644270 192267 644272
rect 104249 644267 104315 644270
rect 192201 644267 192267 644270
rect 196893 644330 196959 644333
rect 199009 644330 199075 644333
rect 196893 644328 199075 644330
rect 196893 644272 196898 644328
rect 196954 644272 199014 644328
rect 199070 644272 199075 644328
rect 196893 644270 199075 644272
rect 196893 644267 196959 644270
rect 199009 644267 199075 644270
rect 199285 644330 199351 644333
rect 236177 644330 236243 644333
rect 240685 644330 240751 644333
rect 199285 644328 199762 644330
rect 199285 644272 199290 644328
rect 199346 644272 199762 644328
rect 199285 644270 199762 644272
rect 199285 644267 199351 644270
rect 189717 644058 189783 644061
rect 180750 644056 189783 644058
rect 180750 644000 189722 644056
rect 189778 644000 189783 644056
rect 180750 643998 189783 644000
rect 153101 643922 153167 643925
rect 180750 643922 180810 643998
rect 189717 643995 189783 643998
rect 192753 644058 192819 644061
rect 196525 644058 196591 644061
rect 192753 644056 196591 644058
rect 192753 644000 192758 644056
rect 192814 644000 196530 644056
rect 196586 644000 196591 644056
rect 192753 643998 196591 644000
rect 192753 643995 192819 643998
rect 196525 643995 196591 643998
rect 153101 643920 180810 643922
rect 153101 643864 153106 643920
rect 153162 643864 180810 643920
rect 153101 643862 180810 643864
rect 185534 643862 190470 643922
rect 153101 643859 153167 643862
rect 133873 643650 133939 643653
rect 185534 643650 185594 643862
rect 189717 643786 189783 643789
rect 189717 643784 189826 643786
rect 189717 643728 189722 643784
rect 189778 643728 189826 643784
rect 189717 643723 189826 643728
rect 133873 643648 185594 643650
rect 133873 643592 133878 643648
rect 133934 643592 185594 643648
rect 133873 643590 185594 643592
rect 133873 643587 133939 643590
rect 189766 643242 189826 643723
rect 190410 643650 190470 643862
rect 199702 643786 199762 644270
rect 236177 644328 240751 644330
rect 236177 644272 236182 644328
rect 236238 644272 240690 644328
rect 240746 644272 240751 644328
rect 236177 644270 240751 644272
rect 236177 644267 236243 644270
rect 240685 644267 240751 644270
rect 580441 644058 580507 644061
rect 583520 644058 584960 644148
rect 580441 644056 584960 644058
rect 580441 644000 580446 644056
rect 580502 644000 584960 644056
rect 580441 643998 584960 644000
rect 580441 643995 580507 643998
rect 583520 643908 584960 643998
rect 202505 643786 202571 643789
rect 199702 643784 202571 643786
rect 199702 643728 202510 643784
rect 202566 643728 202571 643784
rect 199702 643726 202571 643728
rect 202505 643723 202571 643726
rect 202781 643786 202847 643789
rect 202781 643784 205650 643786
rect 202781 643728 202786 643784
rect 202842 643728 205650 643784
rect 202781 643726 205650 643728
rect 202781 643723 202847 643726
rect 192201 643650 192267 643653
rect 190410 643648 192267 643650
rect 190410 643592 192206 643648
rect 192262 643592 192267 643648
rect 190410 643590 192267 643592
rect 192201 643587 192267 643590
rect 192753 643650 192819 643653
rect 196617 643650 196683 643653
rect 192753 643648 196683 643650
rect 192753 643592 192758 643648
rect 192814 643592 196622 643648
rect 196678 643592 196683 643648
rect 192753 643590 196683 643592
rect 192753 643587 192819 643590
rect 196617 643587 196683 643590
rect 198089 643650 198155 643653
rect 199285 643650 199351 643653
rect 198089 643648 199351 643650
rect 198089 643592 198094 643648
rect 198150 643592 199290 643648
rect 199346 643592 199351 643648
rect 198089 643590 199351 643592
rect 198089 643587 198155 643590
rect 199285 643587 199351 643590
rect 199653 643650 199719 643653
rect 202229 643650 202295 643653
rect 199653 643648 202295 643650
rect 199653 643592 199658 643648
rect 199714 643592 202234 643648
rect 202290 643592 202295 643648
rect 199653 643590 202295 643592
rect 205590 643650 205650 643726
rect 208393 643650 208459 643653
rect 205590 643648 208459 643650
rect 205590 643592 208398 643648
rect 208454 643592 208459 643648
rect 205590 643590 208459 643592
rect 199653 643587 199719 643590
rect 202229 643587 202295 643590
rect 208393 643587 208459 643590
rect 192201 643378 192267 643381
rect 190410 643376 192267 643378
rect 190410 643320 192206 643376
rect 192262 643320 192267 643376
rect 190410 643318 192267 643320
rect 190410 643242 190470 643318
rect 192201 643315 192267 643318
rect 189766 643212 190470 643242
rect 189796 643182 190470 643212
rect 202229 643242 202295 643245
rect 206553 643242 206619 643245
rect 202229 643240 206619 643242
rect 202229 643184 202234 643240
rect 202290 643184 206558 643240
rect 206614 643184 206619 643240
rect 202229 643182 206619 643184
rect 202229 643179 202295 643182
rect 206553 643179 206619 643182
rect 190913 642970 190979 642973
rect 190913 642968 191452 642970
rect 190913 642912 190918 642968
rect 190974 642940 191452 642968
rect 190974 642912 191482 642940
rect 190913 642910 191482 642912
rect 190913 642907 190979 642910
rect 191422 642154 191482 642910
rect 236177 642290 236243 642293
rect 241605 642290 241671 642293
rect 236177 642288 241671 642290
rect 236177 642232 236182 642288
rect 236238 642232 241610 642288
rect 241666 642232 241671 642288
rect 236177 642230 241671 642232
rect 236177 642227 236243 642230
rect 241605 642227 241671 642230
rect 192201 642154 192267 642157
rect 191422 642152 192267 642154
rect 191422 642124 192206 642152
rect 191452 642096 192206 642124
rect 192262 642096 192267 642152
rect 191452 642094 192267 642096
rect 192201 642091 192267 642094
rect 459553 640522 459619 640525
rect 468661 640522 468727 640525
rect 459553 640520 468727 640522
rect 459553 640464 459558 640520
rect 459614 640464 468666 640520
rect 468722 640464 468727 640520
rect 459553 640462 468727 640464
rect 459553 640459 459619 640462
rect 468661 640459 468727 640462
rect 469029 640522 469095 640525
rect 471789 640522 471855 640525
rect 469029 640520 471855 640522
rect 469029 640464 469034 640520
rect 469090 640464 471794 640520
rect 471850 640464 471855 640520
rect 469029 640462 471855 640464
rect 469029 640459 469095 640462
rect 471789 640459 471855 640462
rect 230473 639978 230539 639981
rect 230430 639976 230539 639978
rect 230430 639920 230478 639976
rect 230534 639920 230539 639976
rect 230430 639915 230539 639920
rect 224910 639573 224970 639812
rect 230430 639709 230490 639915
rect 230430 639704 230539 639709
rect 230430 639648 230478 639704
rect 230534 639648 230539 639704
rect 230430 639646 230539 639648
rect 230473 639643 230539 639646
rect 224861 639568 224970 639573
rect 224861 639512 224866 639568
rect 224922 639512 224970 639568
rect 224861 639510 224970 639512
rect 224861 639507 224927 639510
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580533 630866 580599 630869
rect 583520 630866 584960 630956
rect 580533 630864 584960 630866
rect 580533 630808 580538 630864
rect 580594 630808 584960 630864
rect 580533 630806 584960 630808
rect 580533 630803 580599 630806
rect 583520 630716 584960 630806
rect 404261 628146 404327 628149
rect 404261 628144 406364 628146
rect 404261 628088 404266 628144
rect 404322 628088 406364 628144
rect 404261 628086 406364 628088
rect 404261 628083 404327 628086
rect 40174 625701 40234 626076
rect 40125 625696 40234 625701
rect 40125 625640 40130 625696
rect 40186 625640 40234 625696
rect 40125 625638 40234 625640
rect 40125 625635 40191 625638
rect 40033 623522 40099 623525
rect 40174 623522 40234 623764
rect 40033 623520 40234 623522
rect 40033 623464 40038 623520
rect 40094 623464 40234 623520
rect 40033 623462 40234 623464
rect 40033 623459 40099 623462
rect -960 619170 480 619260
rect 3785 619170 3851 619173
rect -960 619168 3851 619170
rect -960 619112 3790 619168
rect 3846 619112 3851 619168
rect -960 619110 3851 619112
rect -960 619020 480 619110
rect 3785 619107 3851 619110
rect 580625 617538 580691 617541
rect 583520 617538 584960 617628
rect 580625 617536 584960 617538
rect 580625 617480 580630 617536
rect 580686 617480 584960 617536
rect 580625 617478 584960 617480
rect 580625 617475 580691 617478
rect 583520 617388 584960 617478
rect 40217 606794 40283 606797
rect 40174 606792 40283 606794
rect 40174 606736 40222 606792
rect 40278 606736 40283 606792
rect 40174 606731 40283 606736
rect 40174 606628 40234 606731
rect -960 606114 480 606204
rect 114461 606114 114527 606117
rect -960 606112 114527 606114
rect -960 606056 114466 606112
rect 114522 606056 114527 606112
rect -960 606054 114527 606056
rect -960 605964 480 606054
rect 114461 606051 114527 606054
rect 583520 604060 584960 604300
rect -960 593058 480 593148
rect 3141 593058 3207 593061
rect -960 593056 3207 593058
rect -960 593000 3146 593056
rect 3202 593000 3207 593056
rect -960 592998 3207 593000
rect -960 592908 480 592998
rect 3141 592995 3207 592998
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect 118601 590746 118667 590749
rect 167453 590746 167519 590749
rect 118601 590744 167519 590746
rect 118601 590688 118606 590744
rect 118662 590688 167458 590744
rect 167514 590688 167519 590744
rect 118601 590686 167519 590688
rect 118601 590683 118667 590686
rect 167453 590683 167519 590686
rect 40033 582178 40099 582181
rect 40174 582178 40234 582284
rect 40033 582176 40234 582178
rect 40033 582120 40038 582176
rect 40094 582120 40234 582176
rect 40033 582118 40234 582120
rect 40033 582115 40099 582118
rect 167453 580274 167519 580277
rect 6870 580272 167519 580274
rect 6870 580216 167458 580272
rect 167514 580216 167519 580272
rect 6870 580214 167519 580216
rect -960 580002 480 580092
rect 6870 580002 6930 580214
rect 167453 580211 167519 580214
rect -960 579942 6930 580002
rect -960 579852 480 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 121361 576874 121427 576877
rect 167453 576874 167519 576877
rect 121361 576872 167519 576874
rect 121361 576816 121366 576872
rect 121422 576816 167458 576872
rect 167514 576816 167519 576872
rect 121361 576814 167519 576816
rect 121361 576811 121427 576814
rect 167453 576811 167519 576814
rect -960 566946 480 567036
rect 3693 566946 3759 566949
rect -960 566944 3759 566946
rect -960 566888 3698 566944
rect 3754 566888 3759 566944
rect -960 566886 3759 566888
rect -960 566796 480 566886
rect 3693 566883 3759 566886
rect 580717 564362 580783 564365
rect 583520 564362 584960 564452
rect 580717 564360 584960 564362
rect 580717 564304 580722 564360
rect 580778 564304 584960 564360
rect 580717 564302 584960 564304
rect 580717 564299 580783 564302
rect 583520 564212 584960 564302
rect 391841 559466 391907 559469
rect 391841 559464 394036 559466
rect 391841 559408 391846 559464
rect 391902 559408 394036 559464
rect 391841 559406 394036 559408
rect 391841 559403 391907 559406
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 427813 551578 427879 551581
rect 425868 551576 427879 551578
rect 425868 551520 427818 551576
rect 427874 551520 427879 551576
rect 425868 551518 427879 551520
rect 427813 551515 427879 551518
rect 583520 551020 584960 551260
rect 391381 543554 391447 543557
rect 391381 543552 394036 543554
rect 391381 543496 391386 543552
rect 391442 543496 394036 543552
rect 391381 543494 394036 543496
rect 391381 543491 391447 543494
rect -960 540834 480 540924
rect 3325 540834 3391 540837
rect -960 540832 3391 540834
rect -960 540776 3330 540832
rect 3386 540776 3391 540832
rect -960 540774 3391 540776
rect -960 540684 480 540774
rect 3325 540771 3391 540774
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488746 480 488836
rect 3141 488746 3207 488749
rect -960 488744 3207 488746
rect -960 488688 3146 488744
rect 3202 488688 3207 488744
rect -960 488686 3207 488688
rect -960 488596 480 488686
rect 3141 488683 3207 488686
rect 579613 484666 579679 484669
rect 583520 484666 584960 484756
rect 579613 484664 584960 484666
rect 579613 484608 579618 484664
rect 579674 484608 584960 484664
rect 579613 484606 584960 484608
rect 579613 484603 579679 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436658 480 436748
rect 3325 436658 3391 436661
rect -960 436656 3391 436658
rect -960 436600 3330 436656
rect 3386 436600 3391 436656
rect -960 436598 3391 436600
rect -960 436508 480 436598
rect 3325 436595 3391 436598
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 579613 418298 579679 418301
rect 583520 418298 584960 418388
rect 579613 418296 584960 418298
rect 579613 418240 579618 418296
rect 579674 418240 584960 418296
rect 579613 418238 584960 418240
rect 579613 418235 579679 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579613 378450 579679 378453
rect 583520 378450 584960 378540
rect 579613 378448 584960 378450
rect 579613 378392 579618 378448
rect 579674 378392 584960 378448
rect 579613 378390 584960 378392
rect 579613 378387 579679 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3877 358458 3943 358461
rect -960 358456 3943 358458
rect -960 358400 3882 358456
rect 3938 358400 3943 358456
rect -960 358398 3943 358400
rect -960 358308 480 358398
rect 3877 358395 3943 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3601 319290 3667 319293
rect -960 319288 3667 319290
rect -960 319232 3606 319288
rect 3662 319232 3667 319288
rect -960 319230 3667 319232
rect -960 319140 480 319230
rect 3601 319227 3667 319230
rect 68001 312490 68067 312493
rect 304441 312490 304507 312493
rect 68001 312488 304507 312490
rect 68001 312432 68006 312488
rect 68062 312432 304446 312488
rect 304502 312432 304507 312488
rect 68001 312430 304507 312432
rect 68001 312427 68067 312430
rect 304441 312427 304507 312430
rect 50981 312354 51047 312357
rect 303337 312354 303403 312357
rect 50981 312352 303403 312354
rect 50981 312296 50986 312352
rect 51042 312296 303342 312352
rect 303398 312296 303403 312352
rect 50981 312294 303403 312296
rect 50981 312291 51047 312294
rect 303337 312291 303403 312294
rect 43989 312218 44055 312221
rect 303153 312218 303219 312221
rect 43989 312216 303219 312218
rect 43989 312160 43994 312216
rect 44050 312160 303158 312216
rect 303214 312160 303219 312216
rect 43989 312158 303219 312160
rect 43989 312155 44055 312158
rect 303153 312155 303219 312158
rect 34329 312082 34395 312085
rect 302877 312082 302943 312085
rect 34329 312080 302943 312082
rect 34329 312024 34334 312080
rect 34390 312024 302882 312080
rect 302938 312024 302943 312080
rect 34329 312022 302943 312024
rect 34329 312019 34395 312022
rect 302877 312019 302943 312022
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 3509 311946 3575 311949
rect 300945 311946 301011 311949
rect 3509 311944 301011 311946
rect 3509 311888 3514 311944
rect 3570 311888 300950 311944
rect 301006 311888 301011 311944
rect 583520 311932 584960 312022
rect 3509 311886 301011 311888
rect 3509 311883 3575 311886
rect 300945 311883 301011 311886
rect 29545 310042 29611 310045
rect 31753 310042 31819 310045
rect 29545 310040 31586 310042
rect 29545 309984 29550 310040
rect 29606 309984 31586 310040
rect 29545 309982 31586 309984
rect 29545 309979 29611 309982
rect 31526 309226 31586 309982
rect 31753 310040 35910 310042
rect 31753 309984 31758 310040
rect 31814 309984 35910 310040
rect 31753 309982 35910 309984
rect 31753 309979 31819 309982
rect 35850 309362 35910 309982
rect 302969 309362 303035 309365
rect 35850 309360 303035 309362
rect 35850 309304 302974 309360
rect 303030 309304 303035 309360
rect 35850 309302 303035 309304
rect 302969 309299 303035 309302
rect 315297 309226 315363 309229
rect 31526 309224 315363 309226
rect 31526 309168 315302 309224
rect 315358 309168 315363 309224
rect 31526 309166 315363 309168
rect 315297 309163 315363 309166
rect -960 306234 480 306324
rect 2957 306234 3023 306237
rect -960 306232 3023 306234
rect -960 306176 2962 306232
rect 3018 306176 3023 306232
rect -960 306174 3023 306176
rect -960 306084 480 306174
rect 2957 306171 3023 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579981 272234 580047 272237
rect 583520 272234 584960 272324
rect 579981 272232 584960 272234
rect 579981 272176 579986 272232
rect 580042 272176 584960 272232
rect 579981 272174 584960 272176
rect 579981 272171 580047 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2773 267202 2839 267205
rect -960 267200 2839 267202
rect -960 267144 2778 267200
rect 2834 267144 2839 267200
rect -960 267142 2839 267144
rect -960 267052 480 267142
rect 2773 267139 2839 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 4061 241090 4127 241093
rect -960 241088 4127 241090
rect -960 241032 4066 241088
rect 4122 241032 4127 241088
rect -960 241030 4127 241032
rect -960 240940 480 241030
rect 4061 241027 4127 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580809 219058 580875 219061
rect 583520 219058 584960 219148
rect 580809 219056 584960 219058
rect 580809 219000 580814 219056
rect 580870 219000 584960 219056
rect 580809 218998 584960 219000
rect 580809 218995 580875 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3969 201922 4035 201925
rect -960 201920 4035 201922
rect -960 201864 3974 201920
rect 4030 201864 4035 201920
rect -960 201862 4035 201864
rect -960 201772 480 201862
rect 3969 201859 4035 201862
rect 580717 192538 580783 192541
rect 583520 192538 584960 192628
rect 580717 192536 584960 192538
rect 580717 192480 580722 192536
rect 580778 192480 584960 192536
rect 580717 192478 584960 192480
rect 580717 192475 580783 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3877 188866 3943 188869
rect -960 188864 3943 188866
rect -960 188808 3882 188864
rect 3938 188808 3943 188864
rect -960 188806 3943 188808
rect -960 188716 480 188806
rect 3877 188803 3943 188806
rect 580625 179210 580691 179213
rect 583520 179210 584960 179300
rect 580625 179208 584960 179210
rect 580625 179152 580630 179208
rect 580686 179152 584960 179208
rect 580625 179150 584960 179152
rect 580625 179147 580691 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3785 149834 3851 149837
rect -960 149832 3851 149834
rect -960 149776 3790 149832
rect 3846 149776 3851 149832
rect -960 149774 3851 149776
rect -960 149684 480 149774
rect 3785 149771 3851 149774
rect 580533 139362 580599 139365
rect 583520 139362 584960 139452
rect 580533 139360 584960 139362
rect 580533 139304 580538 139360
rect 580594 139304 584960 139360
rect 580533 139302 584960 139304
rect 580533 139299 580599 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3693 136778 3759 136781
rect -960 136776 3759 136778
rect -960 136720 3698 136776
rect 3754 136720 3759 136776
rect -960 136718 3759 136720
rect -960 136628 480 136718
rect 3693 136715 3759 136718
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 2773 123722 2839 123725
rect -960 123720 2839 123722
rect -960 123664 2778 123720
rect 2834 123664 2839 123720
rect -960 123662 2839 123664
rect -960 123572 480 123662
rect 2773 123659 2839 123662
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 2773 110666 2839 110669
rect -960 110664 2839 110666
rect -960 110608 2778 110664
rect 2834 110608 2839 110664
rect -960 110606 2839 110608
rect -960 110516 480 110606
rect 2773 110603 2839 110606
rect 580349 99514 580415 99517
rect 583520 99514 584960 99604
rect 580349 99512 584960 99514
rect 580349 99456 580354 99512
rect 580410 99456 584960 99512
rect 580349 99454 584960 99456
rect 580349 99451 580415 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2773 71634 2839 71637
rect -960 71632 2839 71634
rect -960 71576 2778 71632
rect 2834 71576 2839 71632
rect -960 71574 2839 71576
rect -960 71484 480 71574
rect 2773 71571 2839 71574
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3141 45522 3207 45525
rect -960 45520 3207 45522
rect -960 45464 3146 45520
rect 3202 45464 3207 45520
rect -960 45462 3207 45464
rect -960 45372 480 45462
rect 3141 45459 3207 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 302141 31378 302207 31381
rect 322197 31378 322263 31381
rect 302141 31376 322263 31378
rect 302141 31320 302146 31376
rect 302202 31320 322202 31376
rect 322258 31320 322263 31376
rect 302141 31318 322263 31320
rect 302141 31315 302207 31318
rect 322197 31315 322263 31318
rect 249057 31242 249123 31245
rect 323577 31242 323643 31245
rect 249057 31240 323643 31242
rect 249057 31184 249062 31240
rect 249118 31184 323582 31240
rect 323638 31184 323643 31240
rect 249057 31182 323643 31184
rect 249057 31179 249123 31182
rect 323577 31179 323643 31182
rect 252461 31106 252527 31109
rect 382917 31106 382983 31109
rect 252461 31104 382983 31106
rect 252461 31048 252466 31104
rect 252522 31048 382922 31104
rect 382978 31048 382983 31104
rect 252461 31046 382983 31048
rect 252461 31043 252527 31046
rect 382917 31043 382983 31046
rect 238753 30970 238819 30973
rect 380157 30970 380223 30973
rect 238753 30968 380223 30970
rect 238753 30912 238758 30968
rect 238814 30912 380162 30968
rect 380218 30912 380223 30968
rect 238753 30910 380223 30912
rect 238753 30907 238819 30910
rect 380157 30907 380223 30910
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 292481 14786 292547 14789
rect 560385 14786 560451 14789
rect 292481 14784 560451 14786
rect 292481 14728 292486 14784
rect 292542 14728 560390 14784
rect 560446 14728 560451 14784
rect 292481 14726 560451 14728
rect 292481 14723 292547 14726
rect 560385 14723 560451 14726
rect 297909 14650 297975 14653
rect 571517 14650 571583 14653
rect 297909 14648 571583 14650
rect 297909 14592 297914 14648
rect 297970 14592 571522 14648
rect 571578 14592 571583 14648
rect 297909 14590 571583 14592
rect 297909 14587 297975 14590
rect 571517 14587 571583 14590
rect 299197 14514 299263 14517
rect 575105 14514 575171 14517
rect 299197 14512 575171 14514
rect 299197 14456 299202 14512
rect 299258 14456 575110 14512
rect 575166 14456 575171 14512
rect 299197 14454 575171 14456
rect 299197 14451 299263 14454
rect 575105 14451 575171 14454
rect 282637 13426 282703 13429
rect 539593 13426 539659 13429
rect 282637 13424 539659 13426
rect 282637 13368 282642 13424
rect 282698 13368 539598 13424
rect 539654 13368 539659 13424
rect 282637 13366 539659 13368
rect 282637 13363 282703 13366
rect 539593 13363 539659 13366
rect 284109 13290 284175 13293
rect 542721 13290 542787 13293
rect 284109 13288 542787 13290
rect 284109 13232 284114 13288
rect 284170 13232 542726 13288
rect 542782 13232 542787 13288
rect 284109 13230 542787 13232
rect 284109 13227 284175 13230
rect 542721 13227 542787 13230
rect 288157 13154 288223 13157
rect 550265 13154 550331 13157
rect 288157 13152 550331 13154
rect 288157 13096 288162 13152
rect 288218 13096 550270 13152
rect 550326 13096 550331 13152
rect 288157 13094 550331 13096
rect 288157 13091 288223 13094
rect 550265 13091 550331 13094
rect 293677 13018 293743 13021
rect 564433 13018 564499 13021
rect 293677 13016 564499 13018
rect 293677 12960 293682 13016
rect 293738 12960 564438 13016
rect 564494 12960 564499 13016
rect 293677 12958 564499 12960
rect 293677 12955 293743 12958
rect 564433 12955 564499 12958
rect 268929 12066 268995 12069
rect 511257 12066 511323 12069
rect 268929 12064 511323 12066
rect 268929 12008 268934 12064
rect 268990 12008 511262 12064
rect 511318 12008 511323 12064
rect 268929 12006 511323 12008
rect 268929 12003 268995 12006
rect 511257 12003 511323 12006
rect 273069 11930 273135 11933
rect 517881 11930 517947 11933
rect 273069 11928 517947 11930
rect 273069 11872 273074 11928
rect 273130 11872 517886 11928
rect 517942 11872 517947 11928
rect 273069 11870 517947 11872
rect 273069 11867 273135 11870
rect 517881 11867 517947 11870
rect 270217 11794 270283 11797
rect 514753 11794 514819 11797
rect 270217 11792 514819 11794
rect 270217 11736 270222 11792
rect 270278 11736 514758 11792
rect 514814 11736 514819 11792
rect 270217 11734 514819 11736
rect 270217 11731 270283 11734
rect 514753 11731 514819 11734
rect 274357 11658 274423 11661
rect 521837 11658 521903 11661
rect 274357 11656 521903 11658
rect 274357 11600 274362 11656
rect 274418 11600 521842 11656
rect 521898 11600 521903 11656
rect 274357 11598 521903 11600
rect 274357 11595 274423 11598
rect 521837 11595 521903 11598
rect 220629 10706 220695 10709
rect 407205 10706 407271 10709
rect 220629 10704 407271 10706
rect 220629 10648 220634 10704
rect 220690 10648 407210 10704
rect 407266 10648 407271 10704
rect 220629 10646 407271 10648
rect 220629 10643 220695 10646
rect 407205 10643 407271 10646
rect 222009 10570 222075 10573
rect 410793 10570 410859 10573
rect 222009 10568 410859 10570
rect 222009 10512 222014 10568
rect 222070 10512 410798 10568
rect 410854 10512 410859 10568
rect 222009 10510 410859 10512
rect 222009 10507 222075 10510
rect 410793 10507 410859 10510
rect 223389 10434 223455 10437
rect 414289 10434 414355 10437
rect 223389 10432 414355 10434
rect 223389 10376 223394 10432
rect 223450 10376 414294 10432
rect 414350 10376 414355 10432
rect 223389 10374 414355 10376
rect 223389 10371 223455 10374
rect 414289 10371 414355 10374
rect 224677 10298 224743 10301
rect 417417 10298 417483 10301
rect 224677 10296 417483 10298
rect 224677 10240 224682 10296
rect 224738 10240 417422 10296
rect 417478 10240 417483 10296
rect 224677 10238 417483 10240
rect 224677 10235 224743 10238
rect 417417 10235 417483 10238
rect 176561 9346 176627 9349
rect 315021 9346 315087 9349
rect 176561 9344 315087 9346
rect 176561 9288 176566 9344
rect 176622 9288 315026 9344
rect 315082 9288 315087 9344
rect 176561 9286 315087 9288
rect 176561 9283 176627 9286
rect 315021 9283 315087 9286
rect 179229 9210 179295 9213
rect 318517 9210 318583 9213
rect 179229 9208 318583 9210
rect 179229 9152 179234 9208
rect 179290 9152 318522 9208
rect 318578 9152 318583 9208
rect 179229 9150 318583 9152
rect 179229 9147 179295 9150
rect 318517 9147 318583 9150
rect 180701 9074 180767 9077
rect 322105 9074 322171 9077
rect 180701 9072 322171 9074
rect 180701 9016 180706 9072
rect 180762 9016 322110 9072
rect 322166 9016 322171 9072
rect 180701 9014 322171 9016
rect 180701 9011 180767 9014
rect 322105 9011 322171 9014
rect 288249 8938 288315 8941
rect 552657 8938 552723 8941
rect 288249 8936 552723 8938
rect 288249 8880 288254 8936
rect 288310 8880 552662 8936
rect 552718 8880 552723 8936
rect 288249 8878 552723 8880
rect 288249 8875 288315 8878
rect 552657 8875 552723 8878
rect 238661 7986 238727 7989
rect 445017 7986 445083 7989
rect 238661 7984 445083 7986
rect 238661 7928 238666 7984
rect 238722 7928 445022 7984
rect 445078 7928 445083 7984
rect 238661 7926 445083 7928
rect 238661 7923 238727 7926
rect 445017 7923 445083 7926
rect 240041 7850 240107 7853
rect 448605 7850 448671 7853
rect 240041 7848 448671 7850
rect 240041 7792 240046 7848
rect 240102 7792 448610 7848
rect 448666 7792 448671 7848
rect 240041 7790 448671 7792
rect 240041 7787 240107 7790
rect 448605 7787 448671 7790
rect 241421 7714 241487 7717
rect 452101 7714 452167 7717
rect 241421 7712 452167 7714
rect 241421 7656 241426 7712
rect 241482 7656 452106 7712
rect 452162 7656 452167 7712
rect 241421 7654 452167 7656
rect 241421 7651 241487 7654
rect 452101 7651 452167 7654
rect 246941 7578 247007 7581
rect 462773 7578 462839 7581
rect 246941 7576 462839 7578
rect 246941 7520 246946 7576
rect 247002 7520 462778 7576
rect 462834 7520 462839 7576
rect 246941 7518 462839 7520
rect 246941 7515 247007 7518
rect 462773 7515 462839 7518
rect 148961 6626 149027 6629
rect 254669 6626 254735 6629
rect 148961 6624 254735 6626
rect -960 6490 480 6580
rect 148961 6568 148966 6624
rect 149022 6568 254674 6624
rect 254730 6568 254735 6624
rect 148961 6566 254735 6568
rect 148961 6563 149027 6566
rect 254669 6563 254735 6566
rect 278589 6626 278655 6629
rect 531313 6626 531379 6629
rect 278589 6624 531379 6626
rect 278589 6568 278594 6624
rect 278650 6568 531318 6624
rect 531374 6568 531379 6624
rect 278589 6566 531379 6568
rect 278589 6563 278655 6566
rect 531313 6563 531379 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 150249 6490 150315 6493
rect 258257 6490 258323 6493
rect 150249 6488 258323 6490
rect 150249 6432 150254 6488
rect 150310 6432 258262 6488
rect 258318 6432 258323 6488
rect 150249 6430 258323 6432
rect 150249 6427 150315 6430
rect 258257 6427 258323 6430
rect 285489 6490 285555 6493
rect 545481 6490 545547 6493
rect 285489 6488 545547 6490
rect 285489 6432 285494 6488
rect 285550 6432 545486 6488
rect 545542 6432 545547 6488
rect 583520 6476 584960 6566
rect 285489 6430 545547 6432
rect 285489 6427 285555 6430
rect 545481 6427 545547 6430
rect 153009 6354 153075 6357
rect 265341 6354 265407 6357
rect 153009 6352 265407 6354
rect 153009 6296 153014 6352
rect 153070 6296 265346 6352
rect 265402 6296 265407 6352
rect 153009 6294 265407 6296
rect 153009 6291 153075 6294
rect 265341 6291 265407 6294
rect 291009 6354 291075 6357
rect 556153 6354 556219 6357
rect 291009 6352 556219 6354
rect 291009 6296 291014 6352
rect 291070 6296 556158 6352
rect 556214 6296 556219 6352
rect 291009 6294 556219 6296
rect 291009 6291 291075 6294
rect 556153 6291 556219 6294
rect 157241 6218 157307 6221
rect 272425 6218 272491 6221
rect 157241 6216 272491 6218
rect 157241 6160 157246 6216
rect 157302 6160 272430 6216
rect 272486 6160 272491 6216
rect 157241 6158 272491 6160
rect 157241 6155 157307 6158
rect 272425 6155 272491 6158
rect 296529 6218 296595 6221
rect 570321 6218 570387 6221
rect 296529 6216 570387 6218
rect 296529 6160 296534 6216
rect 296590 6160 570326 6216
rect 570382 6160 570387 6216
rect 296529 6158 570387 6160
rect 296529 6155 296595 6158
rect 570321 6155 570387 6158
rect 195881 5266 195947 5269
rect 356329 5266 356395 5269
rect 195881 5264 356395 5266
rect 195881 5208 195886 5264
rect 195942 5208 356334 5264
rect 356390 5208 356395 5264
rect 195881 5206 356395 5208
rect 195881 5203 195947 5206
rect 356329 5203 356395 5206
rect 139301 5130 139367 5133
rect 235809 5130 235875 5133
rect 139301 5128 235875 5130
rect 139301 5072 139306 5128
rect 139362 5072 235814 5128
rect 235870 5072 235875 5128
rect 139301 5070 235875 5072
rect 139301 5067 139367 5070
rect 235809 5067 235875 5070
rect 289721 5130 289787 5133
rect 554957 5130 555023 5133
rect 289721 5128 555023 5130
rect 289721 5072 289726 5128
rect 289782 5072 554962 5128
rect 555018 5072 555023 5128
rect 289721 5070 555023 5072
rect 289721 5067 289787 5070
rect 554957 5067 555023 5070
rect 151721 4994 151787 4997
rect 260649 4994 260715 4997
rect 151721 4992 260715 4994
rect 151721 4936 151726 4992
rect 151782 4936 260654 4992
rect 260710 4936 260715 4992
rect 151721 4934 260715 4936
rect 151721 4931 151787 4934
rect 260649 4931 260715 4934
rect 291101 4994 291167 4997
rect 558545 4994 558611 4997
rect 291101 4992 558611 4994
rect 291101 4936 291106 4992
rect 291162 4936 558550 4992
rect 558606 4936 558611 4992
rect 291101 4934 558611 4936
rect 291101 4931 291167 4934
rect 558545 4931 558611 4934
rect 154481 4858 154547 4861
rect 267733 4858 267799 4861
rect 154481 4856 267799 4858
rect 154481 4800 154486 4856
rect 154542 4800 267738 4856
rect 267794 4800 267799 4856
rect 154481 4798 267799 4800
rect 154481 4795 154547 4798
rect 267733 4795 267799 4798
rect 298001 4858 298067 4861
rect 572713 4858 572779 4861
rect 298001 4856 572779 4858
rect 298001 4800 298006 4856
rect 298062 4800 572718 4856
rect 572774 4800 572779 4856
rect 298001 4798 572779 4800
rect 298001 4795 298067 4798
rect 572713 4795 572779 4798
rect 131021 3770 131087 3773
rect 216857 3770 216923 3773
rect 131021 3768 216923 3770
rect 131021 3712 131026 3768
rect 131082 3712 216862 3768
rect 216918 3712 216923 3768
rect 131021 3710 216923 3712
rect 131021 3707 131087 3710
rect 216857 3707 216923 3710
rect 79961 3634 80027 3637
rect 110505 3634 110571 3637
rect 79961 3632 110571 3634
rect 79961 3576 79966 3632
rect 80022 3576 110510 3632
rect 110566 3576 110571 3632
rect 79961 3574 110571 3576
rect 79961 3571 80027 3574
rect 110505 3571 110571 3574
rect 133781 3634 133847 3637
rect 223941 3634 224007 3637
rect 133781 3632 224007 3634
rect 133781 3576 133786 3632
rect 133842 3576 223946 3632
rect 224002 3576 224007 3632
rect 133781 3574 224007 3576
rect 133781 3571 133847 3574
rect 223941 3571 224007 3574
rect 323577 3634 323643 3637
rect 468661 3634 468727 3637
rect 323577 3632 468727 3634
rect 323577 3576 323582 3632
rect 323638 3576 468666 3632
rect 468722 3576 468727 3632
rect 323577 3574 468727 3576
rect 323577 3571 323643 3574
rect 468661 3571 468727 3574
rect 84009 3498 84075 3501
rect 117589 3498 117655 3501
rect 84009 3496 117655 3498
rect 84009 3440 84014 3496
rect 84070 3440 117594 3496
rect 117650 3440 117655 3496
rect 84009 3438 117655 3440
rect 84009 3435 84075 3438
rect 117589 3435 117655 3438
rect 135161 3498 135227 3501
rect 227529 3498 227595 3501
rect 135161 3496 227595 3498
rect 135161 3440 135166 3496
rect 135222 3440 227534 3496
rect 227590 3440 227595 3496
rect 135161 3438 227595 3440
rect 135161 3435 135227 3438
rect 227529 3435 227595 3438
rect 251081 3498 251147 3501
rect 472249 3498 472315 3501
rect 251081 3496 472315 3498
rect 251081 3440 251086 3496
rect 251142 3440 472254 3496
rect 472310 3440 472315 3496
rect 251081 3438 472315 3440
rect 251081 3435 251147 3438
rect 472249 3435 472315 3438
rect 84101 3362 84167 3365
rect 118785 3362 118851 3365
rect 84101 3360 118851 3362
rect 84101 3304 84106 3360
rect 84162 3304 118790 3360
rect 118846 3304 118851 3360
rect 84101 3302 118851 3304
rect 84101 3299 84167 3302
rect 118785 3299 118851 3302
rect 140681 3362 140747 3365
rect 238109 3362 238175 3365
rect 140681 3360 238175 3362
rect 140681 3304 140686 3360
rect 140742 3304 238114 3360
rect 238170 3304 238175 3360
rect 140681 3302 238175 3304
rect 140681 3299 140747 3302
rect 238109 3299 238175 3302
rect 253841 3362 253907 3365
rect 479333 3362 479399 3365
rect 253841 3360 479399 3362
rect 253841 3304 253846 3360
rect 253902 3304 479338 3360
rect 479394 3304 479399 3360
rect 253841 3302 479399 3304
rect 253841 3299 253907 3302
rect 479333 3299 479399 3302
rect 348417 3226 348483 3229
rect 351821 3226 351887 3229
rect 348417 3224 351887 3226
rect 348417 3168 348422 3224
rect 348478 3168 351826 3224
rect 351882 3168 351887 3224
rect 348417 3166 351887 3168
rect 348417 3163 348483 3166
rect 351821 3163 351887 3166
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 312712 27854 316338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 679364 38414 686898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 679364 42134 690618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 679364 45854 694338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 679364 49574 698058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 679364 56414 705242
rect 59514 679364 60134 707162
rect 63234 679364 63854 709082
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 679364 67574 680058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 679364 74414 686898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 679364 78134 690618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 679364 81854 694338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 679364 85574 698058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 679364 92414 705242
rect 95514 679364 96134 707162
rect 99234 679364 99854 709082
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 679364 103574 680058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 679364 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 679364 114134 690618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 679364 117854 694338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 679364 121574 698058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 679364 128414 705242
rect 131514 679364 132134 707162
rect 135234 679364 135854 709082
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 679364 139574 680058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 679364 146414 686898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 679364 150134 690618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 679364 153854 694338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 679364 157574 698058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 679364 164414 705242
rect 167514 679364 168134 707162
rect 171234 679364 171854 709082
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 679364 175574 680058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 679364 182414 686898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 679364 186134 690618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 679364 189854 694338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 679364 193574 698058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 679364 200414 705242
rect 203514 679364 204134 707162
rect 207234 679364 207854 709082
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 679364 211574 680058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 679364 218414 686898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 679364 222134 690618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 679364 225854 694338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 679364 229574 698058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 679364 236414 705242
rect 239514 679364 240134 707162
rect 243234 679364 243854 709082
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 679364 247574 680058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 679364 254414 686898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 679364 258134 690618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 679364 261854 694338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 679364 265574 698058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 679364 272414 705242
rect 275514 679364 276134 707162
rect 279234 679364 279854 709082
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 679364 283574 680058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 679364 290414 686898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 679364 294134 690618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 679364 297854 694338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 679364 301574 698058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 55300 651454 61316 651486
rect 55300 651218 55470 651454
rect 55706 651218 55790 651454
rect 56026 651218 56110 651454
rect 56346 651218 56430 651454
rect 56666 651218 56750 651454
rect 56986 651218 57070 651454
rect 57306 651218 57390 651454
rect 57626 651218 57710 651454
rect 57946 651218 58030 651454
rect 58266 651218 58350 651454
rect 58586 651218 58670 651454
rect 58906 651218 58990 651454
rect 59226 651218 59310 651454
rect 59546 651218 59630 651454
rect 59866 651218 59950 651454
rect 60186 651218 60270 651454
rect 60506 651218 60590 651454
rect 60826 651218 60910 651454
rect 61146 651218 61316 651454
rect 55300 651134 61316 651218
rect 55300 650898 55470 651134
rect 55706 650898 55790 651134
rect 56026 650898 56110 651134
rect 56346 650898 56430 651134
rect 56666 650898 56750 651134
rect 56986 650898 57070 651134
rect 57306 650898 57390 651134
rect 57626 650898 57710 651134
rect 57946 650898 58030 651134
rect 58266 650898 58350 651134
rect 58586 650898 58670 651134
rect 58906 650898 58990 651134
rect 59226 650898 59310 651134
rect 59546 650898 59630 651134
rect 59866 650898 59950 651134
rect 60186 650898 60270 651134
rect 60506 650898 60590 651134
rect 60826 650898 60910 651134
rect 61146 650898 61316 651134
rect 55300 650866 61316 650898
rect 286900 651454 291674 651486
rect 286900 651218 286929 651454
rect 287165 651218 287249 651454
rect 287485 651218 287569 651454
rect 287805 651218 287889 651454
rect 288125 651218 288209 651454
rect 288445 651218 288529 651454
rect 288765 651218 288849 651454
rect 289085 651218 289169 651454
rect 289405 651218 289489 651454
rect 289725 651218 289809 651454
rect 290045 651218 290129 651454
rect 290365 651218 290449 651454
rect 290685 651218 290769 651454
rect 291005 651218 291089 651454
rect 291325 651218 291409 651454
rect 291645 651218 291674 651454
rect 286900 651134 291674 651218
rect 286900 650898 286929 651134
rect 287165 650898 287249 651134
rect 287485 650898 287569 651134
rect 287805 650898 287889 651134
rect 288125 650898 288209 651134
rect 288445 650898 288529 651134
rect 288765 650898 288849 651134
rect 289085 650898 289169 651134
rect 289405 650898 289489 651134
rect 289725 650898 289809 651134
rect 290045 650898 290129 651134
rect 290365 650898 290449 651134
rect 290685 650898 290769 651134
rect 291005 650898 291089 651134
rect 291325 650898 291409 651134
rect 291645 650898 291674 651134
rect 286900 650866 291674 650898
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 44912 633454 52282 633486
rect 44912 633218 44959 633454
rect 45195 633218 45279 633454
rect 45515 633218 45599 633454
rect 45835 633218 45919 633454
rect 46155 633218 46239 633454
rect 46475 633218 46559 633454
rect 46795 633218 46879 633454
rect 47115 633218 47199 633454
rect 47435 633218 47519 633454
rect 47755 633218 47839 633454
rect 48075 633218 48159 633454
rect 48395 633218 48479 633454
rect 48715 633218 48799 633454
rect 49035 633218 49119 633454
rect 49355 633218 49439 633454
rect 49675 633218 49759 633454
rect 49995 633218 50079 633454
rect 50315 633218 50399 633454
rect 50635 633218 50719 633454
rect 50955 633218 51039 633454
rect 51275 633218 51359 633454
rect 51595 633218 51679 633454
rect 51915 633218 51999 633454
rect 52235 633218 52282 633454
rect 44912 633134 52282 633218
rect 44912 632898 44959 633134
rect 45195 632898 45279 633134
rect 45515 632898 45599 633134
rect 45835 632898 45919 633134
rect 46155 632898 46239 633134
rect 46475 632898 46559 633134
rect 46795 632898 46879 633134
rect 47115 632898 47199 633134
rect 47435 632898 47519 633134
rect 47755 632898 47839 633134
rect 48075 632898 48159 633134
rect 48395 632898 48479 633134
rect 48715 632898 48799 633134
rect 49035 632898 49119 633134
rect 49355 632898 49439 633134
rect 49675 632898 49759 633134
rect 49995 632898 50079 633134
rect 50315 632898 50399 633134
rect 50635 632898 50719 633134
rect 50955 632898 51039 633134
rect 51275 632898 51359 633134
rect 51595 632898 51679 633134
rect 51915 632898 51999 633134
rect 52235 632898 52282 633134
rect 44912 632866 52282 632898
rect 295102 633454 300536 633486
rect 295102 633218 295141 633454
rect 295377 633218 295461 633454
rect 295697 633218 295781 633454
rect 296017 633218 296101 633454
rect 296337 633218 296421 633454
rect 296657 633218 296741 633454
rect 296977 633218 297061 633454
rect 297297 633218 297381 633454
rect 297617 633218 297701 633454
rect 297937 633218 298021 633454
rect 298257 633218 298341 633454
rect 298577 633218 298661 633454
rect 298897 633218 298981 633454
rect 299217 633218 299301 633454
rect 299537 633218 299621 633454
rect 299857 633218 299941 633454
rect 300177 633218 300261 633454
rect 300497 633218 300536 633454
rect 295102 633134 300536 633218
rect 295102 632898 295141 633134
rect 295377 632898 295461 633134
rect 295697 632898 295781 633134
rect 296017 632898 296101 633134
rect 296337 632898 296421 633134
rect 296657 632898 296741 633134
rect 296977 632898 297061 633134
rect 297297 632898 297381 633134
rect 297617 632898 297701 633134
rect 297937 632898 298021 633134
rect 298257 632898 298341 633134
rect 298577 632898 298661 633134
rect 298897 632898 298981 633134
rect 299217 632898 299301 633134
rect 299537 632898 299621 633134
rect 299857 632898 299941 633134
rect 300177 632898 300261 633134
rect 300497 632898 300536 633134
rect 295102 632866 300536 632898
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 55300 615454 61316 615486
rect 55300 615218 55470 615454
rect 55706 615218 55790 615454
rect 56026 615218 56110 615454
rect 56346 615218 56430 615454
rect 56666 615218 56750 615454
rect 56986 615218 57070 615454
rect 57306 615218 57390 615454
rect 57626 615218 57710 615454
rect 57946 615218 58030 615454
rect 58266 615218 58350 615454
rect 58586 615218 58670 615454
rect 58906 615218 58990 615454
rect 59226 615218 59310 615454
rect 59546 615218 59630 615454
rect 59866 615218 59950 615454
rect 60186 615218 60270 615454
rect 60506 615218 60590 615454
rect 60826 615218 60910 615454
rect 61146 615218 61316 615454
rect 55300 615134 61316 615218
rect 55300 614898 55470 615134
rect 55706 614898 55790 615134
rect 56026 614898 56110 615134
rect 56346 614898 56430 615134
rect 56666 614898 56750 615134
rect 56986 614898 57070 615134
rect 57306 614898 57390 615134
rect 57626 614898 57710 615134
rect 57946 614898 58030 615134
rect 58266 614898 58350 615134
rect 58586 614898 58670 615134
rect 58906 614898 58990 615134
rect 59226 614898 59310 615134
rect 59546 614898 59630 615134
rect 59866 614898 59950 615134
rect 60186 614898 60270 615134
rect 60506 614898 60590 615134
rect 60826 614898 60910 615134
rect 61146 614898 61316 615134
rect 55300 614866 61316 614898
rect 286900 615454 291674 615486
rect 286900 615218 286929 615454
rect 287165 615218 287249 615454
rect 287485 615218 287569 615454
rect 287805 615218 287889 615454
rect 288125 615218 288209 615454
rect 288445 615218 288529 615454
rect 288765 615218 288849 615454
rect 289085 615218 289169 615454
rect 289405 615218 289489 615454
rect 289725 615218 289809 615454
rect 290045 615218 290129 615454
rect 290365 615218 290449 615454
rect 290685 615218 290769 615454
rect 291005 615218 291089 615454
rect 291325 615218 291409 615454
rect 291645 615218 291674 615454
rect 286900 615134 291674 615218
rect 286900 614898 286929 615134
rect 287165 614898 287249 615134
rect 287485 614898 287569 615134
rect 287805 614898 287889 615134
rect 288125 614898 288209 615134
rect 288445 614898 288529 615134
rect 288765 614898 288849 615134
rect 289085 614898 289169 615134
rect 289405 614898 289489 615134
rect 289725 614898 289809 615134
rect 290045 614898 290129 615134
rect 290365 614898 290449 615134
rect 290685 614898 290769 615134
rect 291005 614898 291089 615134
rect 291325 614898 291409 615134
rect 291645 614898 291674 615134
rect 286900 614866 291674 614898
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 44912 597454 52282 597486
rect 44912 597218 44959 597454
rect 45195 597218 45279 597454
rect 45515 597218 45599 597454
rect 45835 597218 45919 597454
rect 46155 597218 46239 597454
rect 46475 597218 46559 597454
rect 46795 597218 46879 597454
rect 47115 597218 47199 597454
rect 47435 597218 47519 597454
rect 47755 597218 47839 597454
rect 48075 597218 48159 597454
rect 48395 597218 48479 597454
rect 48715 597218 48799 597454
rect 49035 597218 49119 597454
rect 49355 597218 49439 597454
rect 49675 597218 49759 597454
rect 49995 597218 50079 597454
rect 50315 597218 50399 597454
rect 50635 597218 50719 597454
rect 50955 597218 51039 597454
rect 51275 597218 51359 597454
rect 51595 597218 51679 597454
rect 51915 597218 51999 597454
rect 52235 597218 52282 597454
rect 44912 597134 52282 597218
rect 44912 596898 44959 597134
rect 45195 596898 45279 597134
rect 45515 596898 45599 597134
rect 45835 596898 45919 597134
rect 46155 596898 46239 597134
rect 46475 596898 46559 597134
rect 46795 596898 46879 597134
rect 47115 596898 47199 597134
rect 47435 596898 47519 597134
rect 47755 596898 47839 597134
rect 48075 596898 48159 597134
rect 48395 596898 48479 597134
rect 48715 596898 48799 597134
rect 49035 596898 49119 597134
rect 49355 596898 49439 597134
rect 49675 596898 49759 597134
rect 49995 596898 50079 597134
rect 50315 596898 50399 597134
rect 50635 596898 50719 597134
rect 50955 596898 51039 597134
rect 51275 596898 51359 597134
rect 51595 596898 51679 597134
rect 51915 596898 51999 597134
rect 52235 596898 52282 597134
rect 44912 596866 52282 596898
rect 295102 597454 300536 597486
rect 295102 597218 295141 597454
rect 295377 597218 295461 597454
rect 295697 597218 295781 597454
rect 296017 597218 296101 597454
rect 296337 597218 296421 597454
rect 296657 597218 296741 597454
rect 296977 597218 297061 597454
rect 297297 597218 297381 597454
rect 297617 597218 297701 597454
rect 297937 597218 298021 597454
rect 298257 597218 298341 597454
rect 298577 597218 298661 597454
rect 298897 597218 298981 597454
rect 299217 597218 299301 597454
rect 299537 597218 299621 597454
rect 299857 597218 299941 597454
rect 300177 597218 300261 597454
rect 300497 597218 300536 597454
rect 295102 597134 300536 597218
rect 295102 596898 295141 597134
rect 295377 596898 295461 597134
rect 295697 596898 295781 597134
rect 296017 596898 296101 597134
rect 296337 596898 296421 597134
rect 296657 596898 296741 597134
rect 296977 596898 297061 597134
rect 297297 596898 297381 597134
rect 297617 596898 297701 597134
rect 297937 596898 298021 597134
rect 298257 596898 298341 597134
rect 298577 596898 298661 597134
rect 298897 596898 298981 597134
rect 299217 596898 299301 597134
rect 299537 596898 299621 597134
rect 299857 596898 299941 597134
rect 300177 596898 300261 597134
rect 300497 596898 300536 597134
rect 295102 596866 300536 596898
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 286900 579454 291674 579486
rect 286900 579218 286929 579454
rect 287165 579218 287249 579454
rect 287485 579218 287569 579454
rect 287805 579218 287889 579454
rect 288125 579218 288209 579454
rect 288445 579218 288529 579454
rect 288765 579218 288849 579454
rect 289085 579218 289169 579454
rect 289405 579218 289489 579454
rect 289725 579218 289809 579454
rect 290045 579218 290129 579454
rect 290365 579218 290449 579454
rect 290685 579218 290769 579454
rect 291005 579218 291089 579454
rect 291325 579218 291409 579454
rect 291645 579218 291674 579454
rect 286900 579134 291674 579218
rect 286900 578898 286929 579134
rect 287165 578898 287249 579134
rect 287485 578898 287569 579134
rect 287805 578898 287889 579134
rect 288125 578898 288209 579134
rect 288445 578898 288529 579134
rect 288765 578898 288849 579134
rect 289085 578898 289169 579134
rect 289405 578898 289489 579134
rect 289725 578898 289809 579134
rect 290045 578898 290129 579134
rect 290365 578898 290449 579134
rect 290685 578898 290769 579134
rect 291005 578898 291089 579134
rect 291325 578898 291409 579134
rect 291645 578898 291674 579134
rect 286900 578866 291674 578898
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 312712 31574 320058
rect 37794 543454 38414 556000
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 312712 38414 326898
rect 41514 547174 42134 556000
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 312712 42134 330618
rect 45234 550894 45854 556000
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 312712 45854 334338
rect 48954 554614 49574 556000
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 312712 49574 338058
rect 55794 525454 56414 556000
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 312712 56414 344898
rect 59514 529174 60134 556000
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 312712 60134 348618
rect 63234 532894 63854 556000
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 312712 63854 316338
rect 66954 536614 67574 556000
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 312712 67574 320058
rect 73794 543454 74414 556000
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 312712 74414 326898
rect 77514 547174 78134 556000
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 312712 78134 330618
rect 81234 550894 81854 556000
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 312712 81854 334338
rect 84954 554614 85574 556000
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 312712 85574 338058
rect 91794 525454 92414 556000
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 312712 92414 344898
rect 95514 529174 96134 556000
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 312712 96134 348618
rect 99234 532894 99854 556000
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 312712 99854 316338
rect 102954 536614 103574 556000
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 312712 103574 320058
rect 109794 543454 110414 556000
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 312712 110414 326898
rect 113514 547174 114134 556000
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 312712 114134 330618
rect 117234 550894 117854 556000
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 312712 117854 334338
rect 120954 554614 121574 556000
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 312712 121574 338058
rect 127794 525454 128414 556000
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 312712 128414 344898
rect 131514 529174 132134 556000
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 312712 132134 348618
rect 135234 532894 135854 556000
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 312712 135854 316338
rect 138954 536614 139574 556000
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 312712 139574 320058
rect 145794 543454 146414 556000
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 312712 146414 326898
rect 149514 547174 150134 556000
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 312712 150134 330618
rect 153234 550894 153854 556000
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 312712 153854 334338
rect 156954 554614 157574 556000
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 312712 157574 338058
rect 163794 525454 164414 556000
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 312712 164414 344898
rect 167514 529174 168134 556000
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 312712 168134 348618
rect 171234 532894 171854 556000
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 312712 171854 316338
rect 174954 536614 175574 556000
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 312712 175574 320058
rect 181794 543454 182414 556000
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 312712 182414 326898
rect 185514 547174 186134 556000
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 312712 186134 330618
rect 189234 550894 189854 556000
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 312712 189854 334338
rect 192954 554614 193574 556000
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 312712 193574 338058
rect 199794 525454 200414 556000
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 312712 200414 344898
rect 203514 529174 204134 556000
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 312712 204134 348618
rect 207234 532894 207854 556000
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 312712 207854 316338
rect 210954 536614 211574 556000
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 312712 211574 320058
rect 217794 543454 218414 556000
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 312712 218414 326898
rect 221514 547174 222134 556000
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 312712 222134 330618
rect 225234 550894 225854 556000
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 312712 225854 334338
rect 228954 554614 229574 556000
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 312712 229574 338058
rect 235794 525454 236414 556000
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 312712 236414 344898
rect 239514 529174 240134 556000
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 312712 240134 348618
rect 243234 532894 243854 556000
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 312712 243854 316338
rect 246954 536614 247574 556000
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 312712 247574 320058
rect 253794 543454 254414 556000
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 312712 254414 326898
rect 257514 547174 258134 556000
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 312712 258134 330618
rect 261234 550894 261854 556000
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 312712 261854 334338
rect 264954 554614 265574 556000
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 312712 265574 338058
rect 271794 525454 272414 556000
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 312712 272414 344898
rect 275514 529174 276134 556000
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 312712 276134 348618
rect 279234 532894 279854 556000
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 312712 279854 316338
rect 282954 536614 283574 556000
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 312712 283574 320058
rect 289794 543454 290414 556000
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 312712 290414 326898
rect 293514 547174 294134 556000
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 312712 294134 330618
rect 297234 550894 297854 556000
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 312712 297854 334338
rect 300954 554614 301574 556000
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 312712 301574 338058
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 23514 277174 24134 312618
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 32208 291454 32528 291486
rect 32208 291218 32250 291454
rect 32486 291218 32528 291454
rect 32208 291134 32528 291218
rect 32208 290898 32250 291134
rect 32486 290898 32528 291134
rect 32208 290866 32528 290898
rect 62928 291454 63248 291486
rect 62928 291218 62970 291454
rect 63206 291218 63248 291454
rect 62928 291134 63248 291218
rect 62928 290898 62970 291134
rect 63206 290898 63248 291134
rect 62928 290866 63248 290898
rect 93648 291454 93968 291486
rect 93648 291218 93690 291454
rect 93926 291218 93968 291454
rect 93648 291134 93968 291218
rect 93648 290898 93690 291134
rect 93926 290898 93968 291134
rect 93648 290866 93968 290898
rect 124368 291454 124688 291486
rect 124368 291218 124410 291454
rect 124646 291218 124688 291454
rect 124368 291134 124688 291218
rect 124368 290898 124410 291134
rect 124646 290898 124688 291134
rect 124368 290866 124688 290898
rect 155088 291454 155408 291486
rect 155088 291218 155130 291454
rect 155366 291218 155408 291454
rect 155088 291134 155408 291218
rect 155088 290898 155130 291134
rect 155366 290898 155408 291134
rect 155088 290866 155408 290898
rect 185808 291454 186128 291486
rect 185808 291218 185850 291454
rect 186086 291218 186128 291454
rect 185808 291134 186128 291218
rect 185808 290898 185850 291134
rect 186086 290898 186128 291134
rect 185808 290866 186128 290898
rect 216528 291454 216848 291486
rect 216528 291218 216570 291454
rect 216806 291218 216848 291454
rect 216528 291134 216848 291218
rect 216528 290898 216570 291134
rect 216806 290898 216848 291134
rect 216528 290866 216848 290898
rect 247248 291454 247568 291486
rect 247248 291218 247290 291454
rect 247526 291218 247568 291454
rect 247248 291134 247568 291218
rect 247248 290898 247290 291134
rect 247526 290898 247568 291134
rect 247248 290866 247568 290898
rect 277968 291454 278288 291486
rect 277968 291218 278010 291454
rect 278246 291218 278288 291454
rect 277968 291134 278288 291218
rect 277968 290898 278010 291134
rect 278246 290898 278288 291134
rect 277968 290866 278288 290898
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 47568 273454 47888 273486
rect 47568 273218 47610 273454
rect 47846 273218 47888 273454
rect 47568 273134 47888 273218
rect 47568 272898 47610 273134
rect 47846 272898 47888 273134
rect 47568 272866 47888 272898
rect 78288 273454 78608 273486
rect 78288 273218 78330 273454
rect 78566 273218 78608 273454
rect 78288 273134 78608 273218
rect 78288 272898 78330 273134
rect 78566 272898 78608 273134
rect 78288 272866 78608 272898
rect 109008 273454 109328 273486
rect 109008 273218 109050 273454
rect 109286 273218 109328 273454
rect 109008 273134 109328 273218
rect 109008 272898 109050 273134
rect 109286 272898 109328 273134
rect 109008 272866 109328 272898
rect 139728 273454 140048 273486
rect 139728 273218 139770 273454
rect 140006 273218 140048 273454
rect 139728 273134 140048 273218
rect 139728 272898 139770 273134
rect 140006 272898 140048 273134
rect 139728 272866 140048 272898
rect 170448 273454 170768 273486
rect 170448 273218 170490 273454
rect 170726 273218 170768 273454
rect 170448 273134 170768 273218
rect 170448 272898 170490 273134
rect 170726 272898 170768 273134
rect 170448 272866 170768 272898
rect 201168 273454 201488 273486
rect 201168 273218 201210 273454
rect 201446 273218 201488 273454
rect 201168 273134 201488 273218
rect 201168 272898 201210 273134
rect 201446 272898 201488 273134
rect 201168 272866 201488 272898
rect 231888 273454 232208 273486
rect 231888 273218 231930 273454
rect 232166 273218 232208 273454
rect 231888 273134 232208 273218
rect 231888 272898 231930 273134
rect 232166 272898 232208 273134
rect 231888 272866 232208 272898
rect 262608 273454 262928 273486
rect 262608 273218 262650 273454
rect 262886 273218 262928 273454
rect 262608 273134 262928 273218
rect 262608 272898 262650 273134
rect 262886 272898 262928 273134
rect 262608 272866 262928 272898
rect 293328 273454 293648 273486
rect 293328 273218 293370 273454
rect 293606 273218 293648 273454
rect 293328 273134 293648 273218
rect 293328 272898 293370 273134
rect 293606 272898 293648 273134
rect 293328 272866 293648 272898
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 32208 255454 32528 255486
rect 32208 255218 32250 255454
rect 32486 255218 32528 255454
rect 32208 255134 32528 255218
rect 32208 254898 32250 255134
rect 32486 254898 32528 255134
rect 32208 254866 32528 254898
rect 62928 255454 63248 255486
rect 62928 255218 62970 255454
rect 63206 255218 63248 255454
rect 62928 255134 63248 255218
rect 62928 254898 62970 255134
rect 63206 254898 63248 255134
rect 62928 254866 63248 254898
rect 93648 255454 93968 255486
rect 93648 255218 93690 255454
rect 93926 255218 93968 255454
rect 93648 255134 93968 255218
rect 93648 254898 93690 255134
rect 93926 254898 93968 255134
rect 93648 254866 93968 254898
rect 124368 255454 124688 255486
rect 124368 255218 124410 255454
rect 124646 255218 124688 255454
rect 124368 255134 124688 255218
rect 124368 254898 124410 255134
rect 124646 254898 124688 255134
rect 124368 254866 124688 254898
rect 155088 255454 155408 255486
rect 155088 255218 155130 255454
rect 155366 255218 155408 255454
rect 155088 255134 155408 255218
rect 155088 254898 155130 255134
rect 155366 254898 155408 255134
rect 155088 254866 155408 254898
rect 185808 255454 186128 255486
rect 185808 255218 185850 255454
rect 186086 255218 186128 255454
rect 185808 255134 186128 255218
rect 185808 254898 185850 255134
rect 186086 254898 186128 255134
rect 185808 254866 186128 254898
rect 216528 255454 216848 255486
rect 216528 255218 216570 255454
rect 216806 255218 216848 255454
rect 216528 255134 216848 255218
rect 216528 254898 216570 255134
rect 216806 254898 216848 255134
rect 216528 254866 216848 254898
rect 247248 255454 247568 255486
rect 247248 255218 247290 255454
rect 247526 255218 247568 255454
rect 247248 255134 247568 255218
rect 247248 254898 247290 255134
rect 247526 254898 247568 255134
rect 247248 254866 247568 254898
rect 277968 255454 278288 255486
rect 277968 255218 278010 255454
rect 278246 255218 278288 255454
rect 277968 255134 278288 255218
rect 277968 254898 278010 255134
rect 278246 254898 278288 255134
rect 277968 254866 278288 254898
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 47568 237454 47888 237486
rect 47568 237218 47610 237454
rect 47846 237218 47888 237454
rect 47568 237134 47888 237218
rect 47568 236898 47610 237134
rect 47846 236898 47888 237134
rect 47568 236866 47888 236898
rect 78288 237454 78608 237486
rect 78288 237218 78330 237454
rect 78566 237218 78608 237454
rect 78288 237134 78608 237218
rect 78288 236898 78330 237134
rect 78566 236898 78608 237134
rect 78288 236866 78608 236898
rect 109008 237454 109328 237486
rect 109008 237218 109050 237454
rect 109286 237218 109328 237454
rect 109008 237134 109328 237218
rect 109008 236898 109050 237134
rect 109286 236898 109328 237134
rect 109008 236866 109328 236898
rect 139728 237454 140048 237486
rect 139728 237218 139770 237454
rect 140006 237218 140048 237454
rect 139728 237134 140048 237218
rect 139728 236898 139770 237134
rect 140006 236898 140048 237134
rect 139728 236866 140048 236898
rect 170448 237454 170768 237486
rect 170448 237218 170490 237454
rect 170726 237218 170768 237454
rect 170448 237134 170768 237218
rect 170448 236898 170490 237134
rect 170726 236898 170768 237134
rect 170448 236866 170768 236898
rect 201168 237454 201488 237486
rect 201168 237218 201210 237454
rect 201446 237218 201488 237454
rect 201168 237134 201488 237218
rect 201168 236898 201210 237134
rect 201446 236898 201488 237134
rect 201168 236866 201488 236898
rect 231888 237454 232208 237486
rect 231888 237218 231930 237454
rect 232166 237218 232208 237454
rect 231888 237134 232208 237218
rect 231888 236898 231930 237134
rect 232166 236898 232208 237134
rect 231888 236866 232208 236898
rect 262608 237454 262928 237486
rect 262608 237218 262650 237454
rect 262886 237218 262928 237454
rect 262608 237134 262928 237218
rect 262608 236898 262650 237134
rect 262886 236898 262928 237134
rect 262608 236866 262928 236898
rect 293328 237454 293648 237486
rect 293328 237218 293370 237454
rect 293606 237218 293648 237454
rect 293328 237134 293648 237218
rect 293328 236898 293370 237134
rect 293606 236898 293648 237134
rect 293328 236866 293648 236898
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 32208 219454 32528 219486
rect 32208 219218 32250 219454
rect 32486 219218 32528 219454
rect 32208 219134 32528 219218
rect 32208 218898 32250 219134
rect 32486 218898 32528 219134
rect 32208 218866 32528 218898
rect 62928 219454 63248 219486
rect 62928 219218 62970 219454
rect 63206 219218 63248 219454
rect 62928 219134 63248 219218
rect 62928 218898 62970 219134
rect 63206 218898 63248 219134
rect 62928 218866 63248 218898
rect 93648 219454 93968 219486
rect 93648 219218 93690 219454
rect 93926 219218 93968 219454
rect 93648 219134 93968 219218
rect 93648 218898 93690 219134
rect 93926 218898 93968 219134
rect 93648 218866 93968 218898
rect 124368 219454 124688 219486
rect 124368 219218 124410 219454
rect 124646 219218 124688 219454
rect 124368 219134 124688 219218
rect 124368 218898 124410 219134
rect 124646 218898 124688 219134
rect 124368 218866 124688 218898
rect 155088 219454 155408 219486
rect 155088 219218 155130 219454
rect 155366 219218 155408 219454
rect 155088 219134 155408 219218
rect 155088 218898 155130 219134
rect 155366 218898 155408 219134
rect 155088 218866 155408 218898
rect 185808 219454 186128 219486
rect 185808 219218 185850 219454
rect 186086 219218 186128 219454
rect 185808 219134 186128 219218
rect 185808 218898 185850 219134
rect 186086 218898 186128 219134
rect 185808 218866 186128 218898
rect 216528 219454 216848 219486
rect 216528 219218 216570 219454
rect 216806 219218 216848 219454
rect 216528 219134 216848 219218
rect 216528 218898 216570 219134
rect 216806 218898 216848 219134
rect 216528 218866 216848 218898
rect 247248 219454 247568 219486
rect 247248 219218 247290 219454
rect 247526 219218 247568 219454
rect 247248 219134 247568 219218
rect 247248 218898 247290 219134
rect 247526 218898 247568 219134
rect 247248 218866 247568 218898
rect 277968 219454 278288 219486
rect 277968 219218 278010 219454
rect 278246 219218 278288 219454
rect 277968 219134 278288 219218
rect 277968 218898 278010 219134
rect 278246 218898 278288 219134
rect 277968 218866 278288 218898
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 47568 201454 47888 201486
rect 47568 201218 47610 201454
rect 47846 201218 47888 201454
rect 47568 201134 47888 201218
rect 47568 200898 47610 201134
rect 47846 200898 47888 201134
rect 47568 200866 47888 200898
rect 78288 201454 78608 201486
rect 78288 201218 78330 201454
rect 78566 201218 78608 201454
rect 78288 201134 78608 201218
rect 78288 200898 78330 201134
rect 78566 200898 78608 201134
rect 78288 200866 78608 200898
rect 109008 201454 109328 201486
rect 109008 201218 109050 201454
rect 109286 201218 109328 201454
rect 109008 201134 109328 201218
rect 109008 200898 109050 201134
rect 109286 200898 109328 201134
rect 109008 200866 109328 200898
rect 139728 201454 140048 201486
rect 139728 201218 139770 201454
rect 140006 201218 140048 201454
rect 139728 201134 140048 201218
rect 139728 200898 139770 201134
rect 140006 200898 140048 201134
rect 139728 200866 140048 200898
rect 170448 201454 170768 201486
rect 170448 201218 170490 201454
rect 170726 201218 170768 201454
rect 170448 201134 170768 201218
rect 170448 200898 170490 201134
rect 170726 200898 170768 201134
rect 170448 200866 170768 200898
rect 201168 201454 201488 201486
rect 201168 201218 201210 201454
rect 201446 201218 201488 201454
rect 201168 201134 201488 201218
rect 201168 200898 201210 201134
rect 201446 200898 201488 201134
rect 201168 200866 201488 200898
rect 231888 201454 232208 201486
rect 231888 201218 231930 201454
rect 232166 201218 232208 201454
rect 231888 201134 232208 201218
rect 231888 200898 231930 201134
rect 232166 200898 232208 201134
rect 231888 200866 232208 200898
rect 262608 201454 262928 201486
rect 262608 201218 262650 201454
rect 262886 201218 262928 201454
rect 262608 201134 262928 201218
rect 262608 200898 262650 201134
rect 262886 200898 262928 201134
rect 262608 200866 262928 200898
rect 293328 201454 293648 201486
rect 293328 201218 293370 201454
rect 293606 201218 293648 201454
rect 293328 201134 293648 201218
rect 293328 200898 293370 201134
rect 293606 200898 293648 201134
rect 293328 200866 293648 200898
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 32208 183454 32528 183486
rect 32208 183218 32250 183454
rect 32486 183218 32528 183454
rect 32208 183134 32528 183218
rect 32208 182898 32250 183134
rect 32486 182898 32528 183134
rect 32208 182866 32528 182898
rect 62928 183454 63248 183486
rect 62928 183218 62970 183454
rect 63206 183218 63248 183454
rect 62928 183134 63248 183218
rect 62928 182898 62970 183134
rect 63206 182898 63248 183134
rect 62928 182866 63248 182898
rect 93648 183454 93968 183486
rect 93648 183218 93690 183454
rect 93926 183218 93968 183454
rect 93648 183134 93968 183218
rect 93648 182898 93690 183134
rect 93926 182898 93968 183134
rect 93648 182866 93968 182898
rect 124368 183454 124688 183486
rect 124368 183218 124410 183454
rect 124646 183218 124688 183454
rect 124368 183134 124688 183218
rect 124368 182898 124410 183134
rect 124646 182898 124688 183134
rect 124368 182866 124688 182898
rect 155088 183454 155408 183486
rect 155088 183218 155130 183454
rect 155366 183218 155408 183454
rect 155088 183134 155408 183218
rect 155088 182898 155130 183134
rect 155366 182898 155408 183134
rect 155088 182866 155408 182898
rect 185808 183454 186128 183486
rect 185808 183218 185850 183454
rect 186086 183218 186128 183454
rect 185808 183134 186128 183218
rect 185808 182898 185850 183134
rect 186086 182898 186128 183134
rect 185808 182866 186128 182898
rect 216528 183454 216848 183486
rect 216528 183218 216570 183454
rect 216806 183218 216848 183454
rect 216528 183134 216848 183218
rect 216528 182898 216570 183134
rect 216806 182898 216848 183134
rect 216528 182866 216848 182898
rect 247248 183454 247568 183486
rect 247248 183218 247290 183454
rect 247526 183218 247568 183454
rect 247248 183134 247568 183218
rect 247248 182898 247290 183134
rect 247526 182898 247568 183134
rect 247248 182866 247568 182898
rect 277968 183454 278288 183486
rect 277968 183218 278010 183454
rect 278246 183218 278288 183454
rect 277968 183134 278288 183218
rect 277968 182898 278010 183134
rect 278246 182898 278288 183134
rect 277968 182866 278288 182898
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 47568 165454 47888 165486
rect 47568 165218 47610 165454
rect 47846 165218 47888 165454
rect 47568 165134 47888 165218
rect 47568 164898 47610 165134
rect 47846 164898 47888 165134
rect 47568 164866 47888 164898
rect 78288 165454 78608 165486
rect 78288 165218 78330 165454
rect 78566 165218 78608 165454
rect 78288 165134 78608 165218
rect 78288 164898 78330 165134
rect 78566 164898 78608 165134
rect 78288 164866 78608 164898
rect 109008 165454 109328 165486
rect 109008 165218 109050 165454
rect 109286 165218 109328 165454
rect 109008 165134 109328 165218
rect 109008 164898 109050 165134
rect 109286 164898 109328 165134
rect 109008 164866 109328 164898
rect 139728 165454 140048 165486
rect 139728 165218 139770 165454
rect 140006 165218 140048 165454
rect 139728 165134 140048 165218
rect 139728 164898 139770 165134
rect 140006 164898 140048 165134
rect 139728 164866 140048 164898
rect 170448 165454 170768 165486
rect 170448 165218 170490 165454
rect 170726 165218 170768 165454
rect 170448 165134 170768 165218
rect 170448 164898 170490 165134
rect 170726 164898 170768 165134
rect 170448 164866 170768 164898
rect 201168 165454 201488 165486
rect 201168 165218 201210 165454
rect 201446 165218 201488 165454
rect 201168 165134 201488 165218
rect 201168 164898 201210 165134
rect 201446 164898 201488 165134
rect 201168 164866 201488 164898
rect 231888 165454 232208 165486
rect 231888 165218 231930 165454
rect 232166 165218 232208 165454
rect 231888 165134 232208 165218
rect 231888 164898 231930 165134
rect 232166 164898 232208 165134
rect 231888 164866 232208 164898
rect 262608 165454 262928 165486
rect 262608 165218 262650 165454
rect 262886 165218 262928 165454
rect 262608 165134 262928 165218
rect 262608 164898 262650 165134
rect 262886 164898 262928 165134
rect 262608 164866 262928 164898
rect 293328 165454 293648 165486
rect 293328 165218 293370 165454
rect 293606 165218 293648 165454
rect 293328 165134 293648 165218
rect 293328 164898 293370 165134
rect 293606 164898 293648 165134
rect 293328 164866 293648 164898
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 32208 147454 32528 147486
rect 32208 147218 32250 147454
rect 32486 147218 32528 147454
rect 32208 147134 32528 147218
rect 32208 146898 32250 147134
rect 32486 146898 32528 147134
rect 32208 146866 32528 146898
rect 62928 147454 63248 147486
rect 62928 147218 62970 147454
rect 63206 147218 63248 147454
rect 62928 147134 63248 147218
rect 62928 146898 62970 147134
rect 63206 146898 63248 147134
rect 62928 146866 63248 146898
rect 93648 147454 93968 147486
rect 93648 147218 93690 147454
rect 93926 147218 93968 147454
rect 93648 147134 93968 147218
rect 93648 146898 93690 147134
rect 93926 146898 93968 147134
rect 93648 146866 93968 146898
rect 124368 147454 124688 147486
rect 124368 147218 124410 147454
rect 124646 147218 124688 147454
rect 124368 147134 124688 147218
rect 124368 146898 124410 147134
rect 124646 146898 124688 147134
rect 124368 146866 124688 146898
rect 155088 147454 155408 147486
rect 155088 147218 155130 147454
rect 155366 147218 155408 147454
rect 155088 147134 155408 147218
rect 155088 146898 155130 147134
rect 155366 146898 155408 147134
rect 155088 146866 155408 146898
rect 185808 147454 186128 147486
rect 185808 147218 185850 147454
rect 186086 147218 186128 147454
rect 185808 147134 186128 147218
rect 185808 146898 185850 147134
rect 186086 146898 186128 147134
rect 185808 146866 186128 146898
rect 216528 147454 216848 147486
rect 216528 147218 216570 147454
rect 216806 147218 216848 147454
rect 216528 147134 216848 147218
rect 216528 146898 216570 147134
rect 216806 146898 216848 147134
rect 216528 146866 216848 146898
rect 247248 147454 247568 147486
rect 247248 147218 247290 147454
rect 247526 147218 247568 147454
rect 247248 147134 247568 147218
rect 247248 146898 247290 147134
rect 247526 146898 247568 147134
rect 247248 146866 247568 146898
rect 277968 147454 278288 147486
rect 277968 147218 278010 147454
rect 278246 147218 278288 147454
rect 277968 147134 278288 147218
rect 277968 146898 278010 147134
rect 278246 146898 278288 147134
rect 277968 146866 278288 146898
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 47568 129454 47888 129486
rect 47568 129218 47610 129454
rect 47846 129218 47888 129454
rect 47568 129134 47888 129218
rect 47568 128898 47610 129134
rect 47846 128898 47888 129134
rect 47568 128866 47888 128898
rect 78288 129454 78608 129486
rect 78288 129218 78330 129454
rect 78566 129218 78608 129454
rect 78288 129134 78608 129218
rect 78288 128898 78330 129134
rect 78566 128898 78608 129134
rect 78288 128866 78608 128898
rect 109008 129454 109328 129486
rect 109008 129218 109050 129454
rect 109286 129218 109328 129454
rect 109008 129134 109328 129218
rect 109008 128898 109050 129134
rect 109286 128898 109328 129134
rect 109008 128866 109328 128898
rect 139728 129454 140048 129486
rect 139728 129218 139770 129454
rect 140006 129218 140048 129454
rect 139728 129134 140048 129218
rect 139728 128898 139770 129134
rect 140006 128898 140048 129134
rect 139728 128866 140048 128898
rect 170448 129454 170768 129486
rect 170448 129218 170490 129454
rect 170726 129218 170768 129454
rect 170448 129134 170768 129218
rect 170448 128898 170490 129134
rect 170726 128898 170768 129134
rect 170448 128866 170768 128898
rect 201168 129454 201488 129486
rect 201168 129218 201210 129454
rect 201446 129218 201488 129454
rect 201168 129134 201488 129218
rect 201168 128898 201210 129134
rect 201446 128898 201488 129134
rect 201168 128866 201488 128898
rect 231888 129454 232208 129486
rect 231888 129218 231930 129454
rect 232166 129218 232208 129454
rect 231888 129134 232208 129218
rect 231888 128898 231930 129134
rect 232166 128898 232208 129134
rect 231888 128866 232208 128898
rect 262608 129454 262928 129486
rect 262608 129218 262650 129454
rect 262886 129218 262928 129454
rect 262608 129134 262928 129218
rect 262608 128898 262650 129134
rect 262886 128898 262928 129134
rect 262608 128866 262928 128898
rect 293328 129454 293648 129486
rect 293328 129218 293370 129454
rect 293606 129218 293648 129454
rect 293328 129134 293648 129218
rect 293328 128898 293370 129134
rect 293606 128898 293648 129134
rect 293328 128866 293648 128898
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 32208 111454 32528 111486
rect 32208 111218 32250 111454
rect 32486 111218 32528 111454
rect 32208 111134 32528 111218
rect 32208 110898 32250 111134
rect 32486 110898 32528 111134
rect 32208 110866 32528 110898
rect 62928 111454 63248 111486
rect 62928 111218 62970 111454
rect 63206 111218 63248 111454
rect 62928 111134 63248 111218
rect 62928 110898 62970 111134
rect 63206 110898 63248 111134
rect 62928 110866 63248 110898
rect 93648 111454 93968 111486
rect 93648 111218 93690 111454
rect 93926 111218 93968 111454
rect 93648 111134 93968 111218
rect 93648 110898 93690 111134
rect 93926 110898 93968 111134
rect 93648 110866 93968 110898
rect 124368 111454 124688 111486
rect 124368 111218 124410 111454
rect 124646 111218 124688 111454
rect 124368 111134 124688 111218
rect 124368 110898 124410 111134
rect 124646 110898 124688 111134
rect 124368 110866 124688 110898
rect 155088 111454 155408 111486
rect 155088 111218 155130 111454
rect 155366 111218 155408 111454
rect 155088 111134 155408 111218
rect 155088 110898 155130 111134
rect 155366 110898 155408 111134
rect 155088 110866 155408 110898
rect 185808 111454 186128 111486
rect 185808 111218 185850 111454
rect 186086 111218 186128 111454
rect 185808 111134 186128 111218
rect 185808 110898 185850 111134
rect 186086 110898 186128 111134
rect 185808 110866 186128 110898
rect 216528 111454 216848 111486
rect 216528 111218 216570 111454
rect 216806 111218 216848 111454
rect 216528 111134 216848 111218
rect 216528 110898 216570 111134
rect 216806 110898 216848 111134
rect 216528 110866 216848 110898
rect 247248 111454 247568 111486
rect 247248 111218 247290 111454
rect 247526 111218 247568 111454
rect 247248 111134 247568 111218
rect 247248 110898 247290 111134
rect 247526 110898 247568 111134
rect 247248 110866 247568 110898
rect 277968 111454 278288 111486
rect 277968 111218 278010 111454
rect 278246 111218 278288 111454
rect 277968 111134 278288 111218
rect 277968 110898 278010 111134
rect 278246 110898 278288 111134
rect 277968 110866 278288 110898
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 47568 93454 47888 93486
rect 47568 93218 47610 93454
rect 47846 93218 47888 93454
rect 47568 93134 47888 93218
rect 47568 92898 47610 93134
rect 47846 92898 47888 93134
rect 47568 92866 47888 92898
rect 78288 93454 78608 93486
rect 78288 93218 78330 93454
rect 78566 93218 78608 93454
rect 78288 93134 78608 93218
rect 78288 92898 78330 93134
rect 78566 92898 78608 93134
rect 78288 92866 78608 92898
rect 109008 93454 109328 93486
rect 109008 93218 109050 93454
rect 109286 93218 109328 93454
rect 109008 93134 109328 93218
rect 109008 92898 109050 93134
rect 109286 92898 109328 93134
rect 109008 92866 109328 92898
rect 139728 93454 140048 93486
rect 139728 93218 139770 93454
rect 140006 93218 140048 93454
rect 139728 93134 140048 93218
rect 139728 92898 139770 93134
rect 140006 92898 140048 93134
rect 139728 92866 140048 92898
rect 170448 93454 170768 93486
rect 170448 93218 170490 93454
rect 170726 93218 170768 93454
rect 170448 93134 170768 93218
rect 170448 92898 170490 93134
rect 170726 92898 170768 93134
rect 170448 92866 170768 92898
rect 201168 93454 201488 93486
rect 201168 93218 201210 93454
rect 201446 93218 201488 93454
rect 201168 93134 201488 93218
rect 201168 92898 201210 93134
rect 201446 92898 201488 93134
rect 201168 92866 201488 92898
rect 231888 93454 232208 93486
rect 231888 93218 231930 93454
rect 232166 93218 232208 93454
rect 231888 93134 232208 93218
rect 231888 92898 231930 93134
rect 232166 92898 232208 93134
rect 231888 92866 232208 92898
rect 262608 93454 262928 93486
rect 262608 93218 262650 93454
rect 262886 93218 262928 93454
rect 262608 93134 262928 93218
rect 262608 92898 262650 93134
rect 262886 92898 262928 93134
rect 262608 92866 262928 92898
rect 293328 93454 293648 93486
rect 293328 93218 293370 93454
rect 293606 93218 293648 93454
rect 293328 93134 293648 93218
rect 293328 92898 293370 93134
rect 293606 92898 293648 93134
rect 293328 92866 293648 92898
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 32208 75454 32528 75486
rect 32208 75218 32250 75454
rect 32486 75218 32528 75454
rect 32208 75134 32528 75218
rect 32208 74898 32250 75134
rect 32486 74898 32528 75134
rect 32208 74866 32528 74898
rect 62928 75454 63248 75486
rect 62928 75218 62970 75454
rect 63206 75218 63248 75454
rect 62928 75134 63248 75218
rect 62928 74898 62970 75134
rect 63206 74898 63248 75134
rect 62928 74866 63248 74898
rect 93648 75454 93968 75486
rect 93648 75218 93690 75454
rect 93926 75218 93968 75454
rect 93648 75134 93968 75218
rect 93648 74898 93690 75134
rect 93926 74898 93968 75134
rect 93648 74866 93968 74898
rect 124368 75454 124688 75486
rect 124368 75218 124410 75454
rect 124646 75218 124688 75454
rect 124368 75134 124688 75218
rect 124368 74898 124410 75134
rect 124646 74898 124688 75134
rect 124368 74866 124688 74898
rect 155088 75454 155408 75486
rect 155088 75218 155130 75454
rect 155366 75218 155408 75454
rect 155088 75134 155408 75218
rect 155088 74898 155130 75134
rect 155366 74898 155408 75134
rect 155088 74866 155408 74898
rect 185808 75454 186128 75486
rect 185808 75218 185850 75454
rect 186086 75218 186128 75454
rect 185808 75134 186128 75218
rect 185808 74898 185850 75134
rect 186086 74898 186128 75134
rect 185808 74866 186128 74898
rect 216528 75454 216848 75486
rect 216528 75218 216570 75454
rect 216806 75218 216848 75454
rect 216528 75134 216848 75218
rect 216528 74898 216570 75134
rect 216806 74898 216848 75134
rect 216528 74866 216848 74898
rect 247248 75454 247568 75486
rect 247248 75218 247290 75454
rect 247526 75218 247568 75454
rect 247248 75134 247568 75218
rect 247248 74898 247290 75134
rect 247526 74898 247568 75134
rect 247248 74866 247568 74898
rect 277968 75454 278288 75486
rect 277968 75218 278010 75454
rect 278246 75218 278288 75454
rect 277968 75134 278288 75218
rect 277968 74898 278010 75134
rect 278246 74898 278288 75134
rect 277968 74866 278288 74898
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 47568 57454 47888 57486
rect 47568 57218 47610 57454
rect 47846 57218 47888 57454
rect 47568 57134 47888 57218
rect 47568 56898 47610 57134
rect 47846 56898 47888 57134
rect 47568 56866 47888 56898
rect 78288 57454 78608 57486
rect 78288 57218 78330 57454
rect 78566 57218 78608 57454
rect 78288 57134 78608 57218
rect 78288 56898 78330 57134
rect 78566 56898 78608 57134
rect 78288 56866 78608 56898
rect 109008 57454 109328 57486
rect 109008 57218 109050 57454
rect 109286 57218 109328 57454
rect 109008 57134 109328 57218
rect 109008 56898 109050 57134
rect 109286 56898 109328 57134
rect 109008 56866 109328 56898
rect 139728 57454 140048 57486
rect 139728 57218 139770 57454
rect 140006 57218 140048 57454
rect 139728 57134 140048 57218
rect 139728 56898 139770 57134
rect 140006 56898 140048 57134
rect 139728 56866 140048 56898
rect 170448 57454 170768 57486
rect 170448 57218 170490 57454
rect 170726 57218 170768 57454
rect 170448 57134 170768 57218
rect 170448 56898 170490 57134
rect 170726 56898 170768 57134
rect 170448 56866 170768 56898
rect 201168 57454 201488 57486
rect 201168 57218 201210 57454
rect 201446 57218 201488 57454
rect 201168 57134 201488 57218
rect 201168 56898 201210 57134
rect 201446 56898 201488 57134
rect 201168 56866 201488 56898
rect 231888 57454 232208 57486
rect 231888 57218 231930 57454
rect 232166 57218 232208 57454
rect 231888 57134 232208 57218
rect 231888 56898 231930 57134
rect 232166 56898 232208 57134
rect 231888 56866 232208 56898
rect 262608 57454 262928 57486
rect 262608 57218 262650 57454
rect 262886 57218 262928 57454
rect 262608 57134 262928 57218
rect 262608 56898 262650 57134
rect 262886 56898 262928 57134
rect 262608 56866 262928 56898
rect 293328 57454 293648 57486
rect 293328 57218 293370 57454
rect 293606 57218 293648 57454
rect 293328 57134 293648 57218
rect 293328 56898 293370 57134
rect 293606 56898 293648 57134
rect 293328 56866 293648 56898
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 32208 39454 32528 39486
rect 32208 39218 32250 39454
rect 32486 39218 32528 39454
rect 32208 39134 32528 39218
rect 32208 38898 32250 39134
rect 32486 38898 32528 39134
rect 32208 38866 32528 38898
rect 62928 39454 63248 39486
rect 62928 39218 62970 39454
rect 63206 39218 63248 39454
rect 62928 39134 63248 39218
rect 62928 38898 62970 39134
rect 63206 38898 63248 39134
rect 62928 38866 63248 38898
rect 93648 39454 93968 39486
rect 93648 39218 93690 39454
rect 93926 39218 93968 39454
rect 93648 39134 93968 39218
rect 93648 38898 93690 39134
rect 93926 38898 93968 39134
rect 93648 38866 93968 38898
rect 124368 39454 124688 39486
rect 124368 39218 124410 39454
rect 124646 39218 124688 39454
rect 124368 39134 124688 39218
rect 124368 38898 124410 39134
rect 124646 38898 124688 39134
rect 124368 38866 124688 38898
rect 155088 39454 155408 39486
rect 155088 39218 155130 39454
rect 155366 39218 155408 39454
rect 155088 39134 155408 39218
rect 155088 38898 155130 39134
rect 155366 38898 155408 39134
rect 155088 38866 155408 38898
rect 185808 39454 186128 39486
rect 185808 39218 185850 39454
rect 186086 39218 186128 39454
rect 185808 39134 186128 39218
rect 185808 38898 185850 39134
rect 186086 38898 186128 39134
rect 185808 38866 186128 38898
rect 216528 39454 216848 39486
rect 216528 39218 216570 39454
rect 216806 39218 216848 39454
rect 216528 39134 216848 39218
rect 216528 38898 216570 39134
rect 216806 38898 216848 39134
rect 216528 38866 216848 38898
rect 247248 39454 247568 39486
rect 247248 39218 247290 39454
rect 247526 39218 247568 39454
rect 247248 39134 247568 39218
rect 247248 38898 247290 39134
rect 247526 38898 247568 39134
rect 247248 38866 247568 38898
rect 277968 39454 278288 39486
rect 277968 39218 278010 39454
rect 278246 39218 278288 39454
rect 277968 39134 278288 39218
rect 277968 38898 278010 39134
rect 278246 38898 278288 39134
rect 277968 38866 278288 38898
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 28894 27854 32000
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32000
rect 37794 3454 38414 32000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 32000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 10894 45854 32000
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 32000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 32000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 32000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 32000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32000
rect 73794 3454 74414 32000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 32000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 32000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 32000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 32000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 32000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 32000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32000
rect 109794 3454 110414 32000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 32000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 32000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 32000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 32000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 32000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 32000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32000
rect 145794 3454 146414 32000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 32000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 32000
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 32000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 32000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 32000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 32000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32000
rect 181794 3454 182414 32000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 32000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 32000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 32000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 32000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 32000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 32000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32000
rect 217794 3454 218414 32000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 32000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 32000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 32000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 32000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 32000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 32000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32000
rect 253794 3454 254414 32000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 32000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 32000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 32000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 32000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 32000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 32000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32000
rect 289794 3454 290414 32000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 32000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 32000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 32000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 697262 398414 704282
rect 401514 697262 402134 706202
rect 405234 697262 405854 708122
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 697262 409574 698058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 697262 416414 705242
rect 419514 697262 420134 707162
rect 423234 697262 423854 709082
rect 426954 697262 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 697262 434414 704282
rect 437514 697262 438134 706202
rect 441234 697262 441854 708122
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 697262 445574 698058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 697262 452414 705242
rect 455514 697262 456134 707162
rect 459234 697262 459854 709082
rect 462954 697262 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 697262 470414 704282
rect 473514 697262 474134 706202
rect 477234 697262 477854 708122
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 697262 481574 698058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 697262 488414 705242
rect 491514 697262 492134 707162
rect 495234 697262 495854 709082
rect 498954 697262 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 697262 506414 704282
rect 509514 697262 510134 706202
rect 513234 697262 513854 708122
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 697262 517574 698058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 697262 524414 705242
rect 527514 697262 528134 707162
rect 531234 697262 531854 709082
rect 534954 697262 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 697262 542414 704282
rect 545514 697262 546134 706202
rect 549234 697262 549854 708122
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 697262 553574 698058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 697262 560414 705242
rect 394766 687454 398024 687486
rect 394766 687218 394837 687454
rect 395073 687218 395157 687454
rect 395393 687218 395477 687454
rect 395713 687218 395797 687454
rect 396033 687218 396117 687454
rect 396353 687218 396437 687454
rect 396673 687218 396757 687454
rect 396993 687218 397077 687454
rect 397313 687218 397397 687454
rect 397633 687218 397717 687454
rect 397953 687218 398024 687454
rect 394766 687134 398024 687218
rect 394766 686898 394837 687134
rect 395073 686898 395157 687134
rect 395393 686898 395477 687134
rect 395713 686898 395797 687134
rect 396033 686898 396117 687134
rect 396353 686898 396437 687134
rect 396673 686898 396757 687134
rect 396993 686898 397077 687134
rect 397313 686898 397397 687134
rect 397633 686898 397717 687134
rect 397953 686898 398024 687134
rect 394766 686866 398024 686898
rect 461456 687454 462396 687486
rect 461456 687218 461488 687454
rect 461724 687218 461808 687454
rect 462044 687218 462128 687454
rect 462364 687218 462396 687454
rect 461456 687134 462396 687218
rect 461456 686898 461488 687134
rect 461724 686898 461808 687134
rect 462044 686898 462128 687134
rect 462364 686898 462396 687134
rect 461456 686866 462396 686898
rect 538132 687454 546798 687486
rect 538132 687218 538187 687454
rect 538423 687218 538507 687454
rect 538743 687218 538827 687454
rect 539063 687218 539147 687454
rect 539383 687218 539467 687454
rect 539703 687218 539787 687454
rect 540023 687218 540107 687454
rect 540343 687218 540427 687454
rect 540663 687218 540747 687454
rect 540983 687218 541067 687454
rect 541303 687218 541387 687454
rect 541623 687218 541707 687454
rect 541943 687218 542027 687454
rect 542263 687218 542347 687454
rect 542583 687218 542667 687454
rect 542903 687218 542987 687454
rect 543223 687218 543307 687454
rect 543543 687218 543627 687454
rect 543863 687218 543947 687454
rect 544183 687218 544267 687454
rect 544503 687218 544587 687454
rect 544823 687218 544907 687454
rect 545143 687218 545227 687454
rect 545463 687218 545547 687454
rect 545783 687218 545867 687454
rect 546103 687218 546187 687454
rect 546423 687218 546507 687454
rect 546743 687218 546798 687454
rect 538132 687134 546798 687218
rect 538132 686898 538187 687134
rect 538423 686898 538507 687134
rect 538743 686898 538827 687134
rect 539063 686898 539147 687134
rect 539383 686898 539467 687134
rect 539703 686898 539787 687134
rect 540023 686898 540107 687134
rect 540343 686898 540427 687134
rect 540663 686898 540747 687134
rect 540983 686898 541067 687134
rect 541303 686898 541387 687134
rect 541623 686898 541707 687134
rect 541943 686898 542027 687134
rect 542263 686898 542347 687134
rect 542583 686898 542667 687134
rect 542903 686898 542987 687134
rect 543223 686898 543307 687134
rect 543543 686898 543627 687134
rect 543863 686898 543947 687134
rect 544183 686898 544267 687134
rect 544503 686898 544587 687134
rect 544823 686898 544907 687134
rect 545143 686898 545227 687134
rect 545463 686898 545547 687134
rect 545783 686898 545867 687134
rect 546103 686898 546187 687134
rect 546423 686898 546507 687134
rect 546743 686898 546798 687134
rect 538132 686866 546798 686898
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 399978 669454 403236 669486
rect 399978 669218 400049 669454
rect 400285 669218 400369 669454
rect 400605 669218 400689 669454
rect 400925 669218 401009 669454
rect 401245 669218 401329 669454
rect 401565 669218 401649 669454
rect 401885 669218 401969 669454
rect 402205 669218 402289 669454
rect 402525 669218 402609 669454
rect 402845 669218 402929 669454
rect 403165 669218 403236 669454
rect 399978 669134 403236 669218
rect 399978 668898 400049 669134
rect 400285 668898 400369 669134
rect 400605 668898 400689 669134
rect 400925 668898 401009 669134
rect 401245 668898 401329 669134
rect 401565 668898 401649 669134
rect 401885 668898 401969 669134
rect 402205 668898 402289 669134
rect 402525 668898 402609 669134
rect 402845 668898 402929 669134
rect 403165 668898 403236 669134
rect 399978 668866 403236 668898
rect 549206 669454 555800 669486
rect 549206 669218 549345 669454
rect 549581 669218 549665 669454
rect 549901 669218 549985 669454
rect 550221 669218 550305 669454
rect 550541 669218 550625 669454
rect 550861 669218 550945 669454
rect 551181 669218 551265 669454
rect 551501 669218 551585 669454
rect 551821 669218 551905 669454
rect 552141 669218 552225 669454
rect 552461 669218 552545 669454
rect 552781 669218 552865 669454
rect 553101 669218 553185 669454
rect 553421 669218 553505 669454
rect 553741 669218 553825 669454
rect 554061 669218 554145 669454
rect 554381 669218 554465 669454
rect 554701 669218 554785 669454
rect 555021 669218 555105 669454
rect 555341 669218 555425 669454
rect 555661 669218 555800 669454
rect 549206 669134 555800 669218
rect 549206 668898 549345 669134
rect 549581 668898 549665 669134
rect 549901 668898 549985 669134
rect 550221 668898 550305 669134
rect 550541 668898 550625 669134
rect 550861 668898 550945 669134
rect 551181 668898 551265 669134
rect 551501 668898 551585 669134
rect 551821 668898 551905 669134
rect 552141 668898 552225 669134
rect 552461 668898 552545 669134
rect 552781 668898 552865 669134
rect 553101 668898 553185 669134
rect 553421 668898 553505 669134
rect 553741 668898 553825 669134
rect 554061 668898 554145 669134
rect 554381 668898 554465 669134
rect 554701 668898 554785 669134
rect 555021 668898 555105 669134
rect 555341 668898 555425 669134
rect 555661 668898 555800 669134
rect 549206 668866 555800 668898
rect 394766 651454 398024 651486
rect 394766 651218 394837 651454
rect 395073 651218 395157 651454
rect 395393 651218 395477 651454
rect 395713 651218 395797 651454
rect 396033 651218 396117 651454
rect 396353 651218 396437 651454
rect 396673 651218 396757 651454
rect 396993 651218 397077 651454
rect 397313 651218 397397 651454
rect 397633 651218 397717 651454
rect 397953 651218 398024 651454
rect 394766 651134 398024 651218
rect 394766 650898 394837 651134
rect 395073 650898 395157 651134
rect 395393 650898 395477 651134
rect 395713 650898 395797 651134
rect 396033 650898 396117 651134
rect 396353 650898 396437 651134
rect 396673 650898 396757 651134
rect 396993 650898 397077 651134
rect 397313 650898 397397 651134
rect 397633 650898 397717 651134
rect 397953 650898 398024 651134
rect 394766 650866 398024 650898
rect 538132 651454 546798 651486
rect 538132 651218 538187 651454
rect 538423 651218 538507 651454
rect 538743 651218 538827 651454
rect 539063 651218 539147 651454
rect 539383 651218 539467 651454
rect 539703 651218 539787 651454
rect 540023 651218 540107 651454
rect 540343 651218 540427 651454
rect 540663 651218 540747 651454
rect 540983 651218 541067 651454
rect 541303 651218 541387 651454
rect 541623 651218 541707 651454
rect 541943 651218 542027 651454
rect 542263 651218 542347 651454
rect 542583 651218 542667 651454
rect 542903 651218 542987 651454
rect 543223 651218 543307 651454
rect 543543 651218 543627 651454
rect 543863 651218 543947 651454
rect 544183 651218 544267 651454
rect 544503 651218 544587 651454
rect 544823 651218 544907 651454
rect 545143 651218 545227 651454
rect 545463 651218 545547 651454
rect 545783 651218 545867 651454
rect 546103 651218 546187 651454
rect 546423 651218 546507 651454
rect 546743 651218 546798 651454
rect 538132 651134 546798 651218
rect 538132 650898 538187 651134
rect 538423 650898 538507 651134
rect 538743 650898 538827 651134
rect 539063 650898 539147 651134
rect 539383 650898 539467 651134
rect 539703 650898 539787 651134
rect 540023 650898 540107 651134
rect 540343 650898 540427 651134
rect 540663 650898 540747 651134
rect 540983 650898 541067 651134
rect 541303 650898 541387 651134
rect 541623 650898 541707 651134
rect 541943 650898 542027 651134
rect 542263 650898 542347 651134
rect 542583 650898 542667 651134
rect 542903 650898 542987 651134
rect 543223 650898 543307 651134
rect 543543 650898 543627 651134
rect 543863 650898 543947 651134
rect 544183 650898 544267 651134
rect 544503 650898 544587 651134
rect 544823 650898 544907 651134
rect 545143 650898 545227 651134
rect 545463 650898 545547 651134
rect 545783 650898 545867 651134
rect 546103 650898 546187 651134
rect 546423 650898 546507 651134
rect 546743 650898 546798 651134
rect 538132 650866 546798 650898
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 399978 633454 403236 633486
rect 399978 633218 400049 633454
rect 400285 633218 400369 633454
rect 400605 633218 400689 633454
rect 400925 633218 401009 633454
rect 401245 633218 401329 633454
rect 401565 633218 401649 633454
rect 401885 633218 401969 633454
rect 402205 633218 402289 633454
rect 402525 633218 402609 633454
rect 402845 633218 402929 633454
rect 403165 633218 403236 633454
rect 399978 633134 403236 633218
rect 399978 632898 400049 633134
rect 400285 632898 400369 633134
rect 400605 632898 400689 633134
rect 400925 632898 401009 633134
rect 401245 632898 401329 633134
rect 401565 632898 401649 633134
rect 401885 632898 401969 633134
rect 402205 632898 402289 633134
rect 402525 632898 402609 633134
rect 402845 632898 402929 633134
rect 403165 632898 403236 633134
rect 399978 632866 403236 632898
rect 461364 633454 461712 633486
rect 461364 633218 461420 633454
rect 461656 633218 461712 633454
rect 461364 633134 461712 633218
rect 461364 632898 461420 633134
rect 461656 632898 461712 633134
rect 461364 632866 461712 632898
rect 473666 633454 475598 633486
rect 473666 633218 473714 633454
rect 473950 633218 474034 633454
rect 474270 633218 474354 633454
rect 474590 633218 474674 633454
rect 474910 633218 474994 633454
rect 475230 633218 475314 633454
rect 475550 633218 475598 633454
rect 473666 633134 475598 633218
rect 473666 632898 473714 633134
rect 473950 632898 474034 633134
rect 474270 632898 474354 633134
rect 474590 632898 474674 633134
rect 474910 632898 474994 633134
rect 475230 632898 475314 633134
rect 475550 632898 475598 633134
rect 473666 632866 475598 632898
rect 486280 633454 487936 633486
rect 486280 633218 486350 633454
rect 486586 633218 486670 633454
rect 486906 633218 486990 633454
rect 487226 633218 487310 633454
rect 487546 633218 487630 633454
rect 487866 633218 487936 633454
rect 486280 633134 487936 633218
rect 486280 632898 486350 633134
rect 486586 632898 486670 633134
rect 486906 632898 486990 633134
rect 487226 632898 487310 633134
rect 487546 632898 487630 633134
rect 487866 632898 487936 633134
rect 486280 632866 487936 632898
rect 549206 633454 555800 633486
rect 549206 633218 549345 633454
rect 549581 633218 549665 633454
rect 549901 633218 549985 633454
rect 550221 633218 550305 633454
rect 550541 633218 550625 633454
rect 550861 633218 550945 633454
rect 551181 633218 551265 633454
rect 551501 633218 551585 633454
rect 551821 633218 551905 633454
rect 552141 633218 552225 633454
rect 552461 633218 552545 633454
rect 552781 633218 552865 633454
rect 553101 633218 553185 633454
rect 553421 633218 553505 633454
rect 553741 633218 553825 633454
rect 554061 633218 554145 633454
rect 554381 633218 554465 633454
rect 554701 633218 554785 633454
rect 555021 633218 555105 633454
rect 555341 633218 555425 633454
rect 555661 633218 555800 633454
rect 549206 633134 555800 633218
rect 549206 632898 549345 633134
rect 549581 632898 549665 633134
rect 549901 632898 549985 633134
rect 550221 632898 550305 633134
rect 550541 632898 550625 633134
rect 550861 632898 550945 633134
rect 551181 632898 551265 633134
rect 551501 632898 551585 633134
rect 551821 632898 551905 633134
rect 552141 632898 552225 633134
rect 552461 632898 552545 633134
rect 552781 632898 552865 633134
rect 553101 632898 553185 633134
rect 553421 632898 553505 633134
rect 553741 632898 553825 633134
rect 554061 632898 554145 633134
rect 554381 632898 554465 633134
rect 554701 632898 554785 633134
rect 555021 632898 555105 633134
rect 555341 632898 555425 633134
rect 555661 632898 555800 633134
rect 549206 632866 555800 632898
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 397794 579454 398414 605200
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 569600 398414 578898
rect 401514 583174 402134 605200
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 569600 402134 582618
rect 405234 586894 405854 605200
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 569600 405854 586338
rect 408954 590614 409574 605200
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 569600 409574 590058
rect 415794 597454 416414 605200
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 569600 416414 596898
rect 419514 601174 420134 605200
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 569600 420134 600618
rect 423234 604894 423854 605200
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 569600 423854 604338
rect 426954 572614 427574 605200
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 569600 427574 572058
rect 433794 579454 434414 605200
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 404874 561454 405194 561486
rect 404874 561218 404916 561454
rect 405152 561218 405194 561454
rect 404874 561134 405194 561218
rect 404874 560898 404916 561134
rect 405152 560898 405194 561134
rect 404874 560866 405194 560898
rect 414805 561454 415125 561486
rect 414805 561218 414847 561454
rect 415083 561218 415125 561454
rect 414805 561134 415125 561218
rect 414805 560898 414847 561134
rect 415083 560898 415125 561134
rect 414805 560866 415125 560898
rect 399909 543454 400229 543486
rect 399909 543218 399951 543454
rect 400187 543218 400229 543454
rect 399909 543134 400229 543218
rect 399909 542898 399951 543134
rect 400187 542898 400229 543134
rect 399909 542866 400229 542898
rect 409839 543454 410159 543486
rect 409839 543218 409881 543454
rect 410117 543218 410159 543454
rect 409839 543134 410159 543218
rect 409839 542898 409881 543134
rect 410117 542898 410159 543134
rect 409839 542866 410159 542898
rect 419770 543454 420090 543486
rect 419770 543218 419812 543454
rect 420048 543218 420090 543454
rect 419770 543134 420090 543218
rect 419770 542898 419812 543134
rect 420048 542898 420090 543134
rect 419770 542866 420090 542898
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 507454 398414 533600
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 511174 402134 533600
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 514894 405854 533600
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 518614 409574 533600
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 525454 416414 533600
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 529174 420134 533600
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 532894 423854 533600
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 500614 427574 533600
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 583174 438134 605200
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 586894 441854 605200
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 590614 445574 605200
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 597454 452414 605200
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 601174 456134 605200
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 604894 459854 605200
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 572614 463574 605200
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 579454 470414 605200
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 583174 474134 605200
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 586894 477854 605200
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 590614 481574 605200
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 597454 488414 605200
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 601174 492134 605200
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 604894 495854 605200
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 572614 499574 605200
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 579454 506414 605200
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 583174 510134 605200
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 586894 513854 605200
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 590614 517574 605200
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 597454 524414 605200
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 601174 528134 605200
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 604894 531854 605200
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 572614 535574 605200
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 579454 542414 605200
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 583174 546134 605200
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 586894 549854 605200
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 590614 553574 605200
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 597454 560414 605200
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 55470 651218 55706 651454
rect 55790 651218 56026 651454
rect 56110 651218 56346 651454
rect 56430 651218 56666 651454
rect 56750 651218 56986 651454
rect 57070 651218 57306 651454
rect 57390 651218 57626 651454
rect 57710 651218 57946 651454
rect 58030 651218 58266 651454
rect 58350 651218 58586 651454
rect 58670 651218 58906 651454
rect 58990 651218 59226 651454
rect 59310 651218 59546 651454
rect 59630 651218 59866 651454
rect 59950 651218 60186 651454
rect 60270 651218 60506 651454
rect 60590 651218 60826 651454
rect 60910 651218 61146 651454
rect 55470 650898 55706 651134
rect 55790 650898 56026 651134
rect 56110 650898 56346 651134
rect 56430 650898 56666 651134
rect 56750 650898 56986 651134
rect 57070 650898 57306 651134
rect 57390 650898 57626 651134
rect 57710 650898 57946 651134
rect 58030 650898 58266 651134
rect 58350 650898 58586 651134
rect 58670 650898 58906 651134
rect 58990 650898 59226 651134
rect 59310 650898 59546 651134
rect 59630 650898 59866 651134
rect 59950 650898 60186 651134
rect 60270 650898 60506 651134
rect 60590 650898 60826 651134
rect 60910 650898 61146 651134
rect 286929 651218 287165 651454
rect 287249 651218 287485 651454
rect 287569 651218 287805 651454
rect 287889 651218 288125 651454
rect 288209 651218 288445 651454
rect 288529 651218 288765 651454
rect 288849 651218 289085 651454
rect 289169 651218 289405 651454
rect 289489 651218 289725 651454
rect 289809 651218 290045 651454
rect 290129 651218 290365 651454
rect 290449 651218 290685 651454
rect 290769 651218 291005 651454
rect 291089 651218 291325 651454
rect 291409 651218 291645 651454
rect 286929 650898 287165 651134
rect 287249 650898 287485 651134
rect 287569 650898 287805 651134
rect 287889 650898 288125 651134
rect 288209 650898 288445 651134
rect 288529 650898 288765 651134
rect 288849 650898 289085 651134
rect 289169 650898 289405 651134
rect 289489 650898 289725 651134
rect 289809 650898 290045 651134
rect 290129 650898 290365 651134
rect 290449 650898 290685 651134
rect 290769 650898 291005 651134
rect 291089 650898 291325 651134
rect 291409 650898 291645 651134
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 44959 633218 45195 633454
rect 45279 633218 45515 633454
rect 45599 633218 45835 633454
rect 45919 633218 46155 633454
rect 46239 633218 46475 633454
rect 46559 633218 46795 633454
rect 46879 633218 47115 633454
rect 47199 633218 47435 633454
rect 47519 633218 47755 633454
rect 47839 633218 48075 633454
rect 48159 633218 48395 633454
rect 48479 633218 48715 633454
rect 48799 633218 49035 633454
rect 49119 633218 49355 633454
rect 49439 633218 49675 633454
rect 49759 633218 49995 633454
rect 50079 633218 50315 633454
rect 50399 633218 50635 633454
rect 50719 633218 50955 633454
rect 51039 633218 51275 633454
rect 51359 633218 51595 633454
rect 51679 633218 51915 633454
rect 51999 633218 52235 633454
rect 44959 632898 45195 633134
rect 45279 632898 45515 633134
rect 45599 632898 45835 633134
rect 45919 632898 46155 633134
rect 46239 632898 46475 633134
rect 46559 632898 46795 633134
rect 46879 632898 47115 633134
rect 47199 632898 47435 633134
rect 47519 632898 47755 633134
rect 47839 632898 48075 633134
rect 48159 632898 48395 633134
rect 48479 632898 48715 633134
rect 48799 632898 49035 633134
rect 49119 632898 49355 633134
rect 49439 632898 49675 633134
rect 49759 632898 49995 633134
rect 50079 632898 50315 633134
rect 50399 632898 50635 633134
rect 50719 632898 50955 633134
rect 51039 632898 51275 633134
rect 51359 632898 51595 633134
rect 51679 632898 51915 633134
rect 51999 632898 52235 633134
rect 295141 633218 295377 633454
rect 295461 633218 295697 633454
rect 295781 633218 296017 633454
rect 296101 633218 296337 633454
rect 296421 633218 296657 633454
rect 296741 633218 296977 633454
rect 297061 633218 297297 633454
rect 297381 633218 297617 633454
rect 297701 633218 297937 633454
rect 298021 633218 298257 633454
rect 298341 633218 298577 633454
rect 298661 633218 298897 633454
rect 298981 633218 299217 633454
rect 299301 633218 299537 633454
rect 299621 633218 299857 633454
rect 299941 633218 300177 633454
rect 300261 633218 300497 633454
rect 295141 632898 295377 633134
rect 295461 632898 295697 633134
rect 295781 632898 296017 633134
rect 296101 632898 296337 633134
rect 296421 632898 296657 633134
rect 296741 632898 296977 633134
rect 297061 632898 297297 633134
rect 297381 632898 297617 633134
rect 297701 632898 297937 633134
rect 298021 632898 298257 633134
rect 298341 632898 298577 633134
rect 298661 632898 298897 633134
rect 298981 632898 299217 633134
rect 299301 632898 299537 633134
rect 299621 632898 299857 633134
rect 299941 632898 300177 633134
rect 300261 632898 300497 633134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 55470 615218 55706 615454
rect 55790 615218 56026 615454
rect 56110 615218 56346 615454
rect 56430 615218 56666 615454
rect 56750 615218 56986 615454
rect 57070 615218 57306 615454
rect 57390 615218 57626 615454
rect 57710 615218 57946 615454
rect 58030 615218 58266 615454
rect 58350 615218 58586 615454
rect 58670 615218 58906 615454
rect 58990 615218 59226 615454
rect 59310 615218 59546 615454
rect 59630 615218 59866 615454
rect 59950 615218 60186 615454
rect 60270 615218 60506 615454
rect 60590 615218 60826 615454
rect 60910 615218 61146 615454
rect 55470 614898 55706 615134
rect 55790 614898 56026 615134
rect 56110 614898 56346 615134
rect 56430 614898 56666 615134
rect 56750 614898 56986 615134
rect 57070 614898 57306 615134
rect 57390 614898 57626 615134
rect 57710 614898 57946 615134
rect 58030 614898 58266 615134
rect 58350 614898 58586 615134
rect 58670 614898 58906 615134
rect 58990 614898 59226 615134
rect 59310 614898 59546 615134
rect 59630 614898 59866 615134
rect 59950 614898 60186 615134
rect 60270 614898 60506 615134
rect 60590 614898 60826 615134
rect 60910 614898 61146 615134
rect 286929 615218 287165 615454
rect 287249 615218 287485 615454
rect 287569 615218 287805 615454
rect 287889 615218 288125 615454
rect 288209 615218 288445 615454
rect 288529 615218 288765 615454
rect 288849 615218 289085 615454
rect 289169 615218 289405 615454
rect 289489 615218 289725 615454
rect 289809 615218 290045 615454
rect 290129 615218 290365 615454
rect 290449 615218 290685 615454
rect 290769 615218 291005 615454
rect 291089 615218 291325 615454
rect 291409 615218 291645 615454
rect 286929 614898 287165 615134
rect 287249 614898 287485 615134
rect 287569 614898 287805 615134
rect 287889 614898 288125 615134
rect 288209 614898 288445 615134
rect 288529 614898 288765 615134
rect 288849 614898 289085 615134
rect 289169 614898 289405 615134
rect 289489 614898 289725 615134
rect 289809 614898 290045 615134
rect 290129 614898 290365 615134
rect 290449 614898 290685 615134
rect 290769 614898 291005 615134
rect 291089 614898 291325 615134
rect 291409 614898 291645 615134
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 44959 597218 45195 597454
rect 45279 597218 45515 597454
rect 45599 597218 45835 597454
rect 45919 597218 46155 597454
rect 46239 597218 46475 597454
rect 46559 597218 46795 597454
rect 46879 597218 47115 597454
rect 47199 597218 47435 597454
rect 47519 597218 47755 597454
rect 47839 597218 48075 597454
rect 48159 597218 48395 597454
rect 48479 597218 48715 597454
rect 48799 597218 49035 597454
rect 49119 597218 49355 597454
rect 49439 597218 49675 597454
rect 49759 597218 49995 597454
rect 50079 597218 50315 597454
rect 50399 597218 50635 597454
rect 50719 597218 50955 597454
rect 51039 597218 51275 597454
rect 51359 597218 51595 597454
rect 51679 597218 51915 597454
rect 51999 597218 52235 597454
rect 44959 596898 45195 597134
rect 45279 596898 45515 597134
rect 45599 596898 45835 597134
rect 45919 596898 46155 597134
rect 46239 596898 46475 597134
rect 46559 596898 46795 597134
rect 46879 596898 47115 597134
rect 47199 596898 47435 597134
rect 47519 596898 47755 597134
rect 47839 596898 48075 597134
rect 48159 596898 48395 597134
rect 48479 596898 48715 597134
rect 48799 596898 49035 597134
rect 49119 596898 49355 597134
rect 49439 596898 49675 597134
rect 49759 596898 49995 597134
rect 50079 596898 50315 597134
rect 50399 596898 50635 597134
rect 50719 596898 50955 597134
rect 51039 596898 51275 597134
rect 51359 596898 51595 597134
rect 51679 596898 51915 597134
rect 51999 596898 52235 597134
rect 295141 597218 295377 597454
rect 295461 597218 295697 597454
rect 295781 597218 296017 597454
rect 296101 597218 296337 597454
rect 296421 597218 296657 597454
rect 296741 597218 296977 597454
rect 297061 597218 297297 597454
rect 297381 597218 297617 597454
rect 297701 597218 297937 597454
rect 298021 597218 298257 597454
rect 298341 597218 298577 597454
rect 298661 597218 298897 597454
rect 298981 597218 299217 597454
rect 299301 597218 299537 597454
rect 299621 597218 299857 597454
rect 299941 597218 300177 597454
rect 300261 597218 300497 597454
rect 295141 596898 295377 597134
rect 295461 596898 295697 597134
rect 295781 596898 296017 597134
rect 296101 596898 296337 597134
rect 296421 596898 296657 597134
rect 296741 596898 296977 597134
rect 297061 596898 297297 597134
rect 297381 596898 297617 597134
rect 297701 596898 297937 597134
rect 298021 596898 298257 597134
rect 298341 596898 298577 597134
rect 298661 596898 298897 597134
rect 298981 596898 299217 597134
rect 299301 596898 299537 597134
rect 299621 596898 299857 597134
rect 299941 596898 300177 597134
rect 300261 596898 300497 597134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 286929 579218 287165 579454
rect 287249 579218 287485 579454
rect 287569 579218 287805 579454
rect 287889 579218 288125 579454
rect 288209 579218 288445 579454
rect 288529 579218 288765 579454
rect 288849 579218 289085 579454
rect 289169 579218 289405 579454
rect 289489 579218 289725 579454
rect 289809 579218 290045 579454
rect 290129 579218 290365 579454
rect 290449 579218 290685 579454
rect 290769 579218 291005 579454
rect 291089 579218 291325 579454
rect 291409 579218 291645 579454
rect 286929 578898 287165 579134
rect 287249 578898 287485 579134
rect 287569 578898 287805 579134
rect 287889 578898 288125 579134
rect 288209 578898 288445 579134
rect 288529 578898 288765 579134
rect 288849 578898 289085 579134
rect 289169 578898 289405 579134
rect 289489 578898 289725 579134
rect 289809 578898 290045 579134
rect 290129 578898 290365 579134
rect 290449 578898 290685 579134
rect 290769 578898 291005 579134
rect 291089 578898 291325 579134
rect 291409 578898 291645 579134
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 32250 291218 32486 291454
rect 32250 290898 32486 291134
rect 62970 291218 63206 291454
rect 62970 290898 63206 291134
rect 93690 291218 93926 291454
rect 93690 290898 93926 291134
rect 124410 291218 124646 291454
rect 124410 290898 124646 291134
rect 155130 291218 155366 291454
rect 155130 290898 155366 291134
rect 185850 291218 186086 291454
rect 185850 290898 186086 291134
rect 216570 291218 216806 291454
rect 216570 290898 216806 291134
rect 247290 291218 247526 291454
rect 247290 290898 247526 291134
rect 278010 291218 278246 291454
rect 278010 290898 278246 291134
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 47610 273218 47846 273454
rect 47610 272898 47846 273134
rect 78330 273218 78566 273454
rect 78330 272898 78566 273134
rect 109050 273218 109286 273454
rect 109050 272898 109286 273134
rect 139770 273218 140006 273454
rect 139770 272898 140006 273134
rect 170490 273218 170726 273454
rect 170490 272898 170726 273134
rect 201210 273218 201446 273454
rect 201210 272898 201446 273134
rect 231930 273218 232166 273454
rect 231930 272898 232166 273134
rect 262650 273218 262886 273454
rect 262650 272898 262886 273134
rect 293370 273218 293606 273454
rect 293370 272898 293606 273134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 32250 255218 32486 255454
rect 32250 254898 32486 255134
rect 62970 255218 63206 255454
rect 62970 254898 63206 255134
rect 93690 255218 93926 255454
rect 93690 254898 93926 255134
rect 124410 255218 124646 255454
rect 124410 254898 124646 255134
rect 155130 255218 155366 255454
rect 155130 254898 155366 255134
rect 185850 255218 186086 255454
rect 185850 254898 186086 255134
rect 216570 255218 216806 255454
rect 216570 254898 216806 255134
rect 247290 255218 247526 255454
rect 247290 254898 247526 255134
rect 278010 255218 278246 255454
rect 278010 254898 278246 255134
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 47610 237218 47846 237454
rect 47610 236898 47846 237134
rect 78330 237218 78566 237454
rect 78330 236898 78566 237134
rect 109050 237218 109286 237454
rect 109050 236898 109286 237134
rect 139770 237218 140006 237454
rect 139770 236898 140006 237134
rect 170490 237218 170726 237454
rect 170490 236898 170726 237134
rect 201210 237218 201446 237454
rect 201210 236898 201446 237134
rect 231930 237218 232166 237454
rect 231930 236898 232166 237134
rect 262650 237218 262886 237454
rect 262650 236898 262886 237134
rect 293370 237218 293606 237454
rect 293370 236898 293606 237134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 32250 219218 32486 219454
rect 32250 218898 32486 219134
rect 62970 219218 63206 219454
rect 62970 218898 63206 219134
rect 93690 219218 93926 219454
rect 93690 218898 93926 219134
rect 124410 219218 124646 219454
rect 124410 218898 124646 219134
rect 155130 219218 155366 219454
rect 155130 218898 155366 219134
rect 185850 219218 186086 219454
rect 185850 218898 186086 219134
rect 216570 219218 216806 219454
rect 216570 218898 216806 219134
rect 247290 219218 247526 219454
rect 247290 218898 247526 219134
rect 278010 219218 278246 219454
rect 278010 218898 278246 219134
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 47610 201218 47846 201454
rect 47610 200898 47846 201134
rect 78330 201218 78566 201454
rect 78330 200898 78566 201134
rect 109050 201218 109286 201454
rect 109050 200898 109286 201134
rect 139770 201218 140006 201454
rect 139770 200898 140006 201134
rect 170490 201218 170726 201454
rect 170490 200898 170726 201134
rect 201210 201218 201446 201454
rect 201210 200898 201446 201134
rect 231930 201218 232166 201454
rect 231930 200898 232166 201134
rect 262650 201218 262886 201454
rect 262650 200898 262886 201134
rect 293370 201218 293606 201454
rect 293370 200898 293606 201134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 32250 183218 32486 183454
rect 32250 182898 32486 183134
rect 62970 183218 63206 183454
rect 62970 182898 63206 183134
rect 93690 183218 93926 183454
rect 93690 182898 93926 183134
rect 124410 183218 124646 183454
rect 124410 182898 124646 183134
rect 155130 183218 155366 183454
rect 155130 182898 155366 183134
rect 185850 183218 186086 183454
rect 185850 182898 186086 183134
rect 216570 183218 216806 183454
rect 216570 182898 216806 183134
rect 247290 183218 247526 183454
rect 247290 182898 247526 183134
rect 278010 183218 278246 183454
rect 278010 182898 278246 183134
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 47610 165218 47846 165454
rect 47610 164898 47846 165134
rect 78330 165218 78566 165454
rect 78330 164898 78566 165134
rect 109050 165218 109286 165454
rect 109050 164898 109286 165134
rect 139770 165218 140006 165454
rect 139770 164898 140006 165134
rect 170490 165218 170726 165454
rect 170490 164898 170726 165134
rect 201210 165218 201446 165454
rect 201210 164898 201446 165134
rect 231930 165218 232166 165454
rect 231930 164898 232166 165134
rect 262650 165218 262886 165454
rect 262650 164898 262886 165134
rect 293370 165218 293606 165454
rect 293370 164898 293606 165134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 32250 147218 32486 147454
rect 32250 146898 32486 147134
rect 62970 147218 63206 147454
rect 62970 146898 63206 147134
rect 93690 147218 93926 147454
rect 93690 146898 93926 147134
rect 124410 147218 124646 147454
rect 124410 146898 124646 147134
rect 155130 147218 155366 147454
rect 155130 146898 155366 147134
rect 185850 147218 186086 147454
rect 185850 146898 186086 147134
rect 216570 147218 216806 147454
rect 216570 146898 216806 147134
rect 247290 147218 247526 147454
rect 247290 146898 247526 147134
rect 278010 147218 278246 147454
rect 278010 146898 278246 147134
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 47610 129218 47846 129454
rect 47610 128898 47846 129134
rect 78330 129218 78566 129454
rect 78330 128898 78566 129134
rect 109050 129218 109286 129454
rect 109050 128898 109286 129134
rect 139770 129218 140006 129454
rect 139770 128898 140006 129134
rect 170490 129218 170726 129454
rect 170490 128898 170726 129134
rect 201210 129218 201446 129454
rect 201210 128898 201446 129134
rect 231930 129218 232166 129454
rect 231930 128898 232166 129134
rect 262650 129218 262886 129454
rect 262650 128898 262886 129134
rect 293370 129218 293606 129454
rect 293370 128898 293606 129134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 32250 111218 32486 111454
rect 32250 110898 32486 111134
rect 62970 111218 63206 111454
rect 62970 110898 63206 111134
rect 93690 111218 93926 111454
rect 93690 110898 93926 111134
rect 124410 111218 124646 111454
rect 124410 110898 124646 111134
rect 155130 111218 155366 111454
rect 155130 110898 155366 111134
rect 185850 111218 186086 111454
rect 185850 110898 186086 111134
rect 216570 111218 216806 111454
rect 216570 110898 216806 111134
rect 247290 111218 247526 111454
rect 247290 110898 247526 111134
rect 278010 111218 278246 111454
rect 278010 110898 278246 111134
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 47610 93218 47846 93454
rect 47610 92898 47846 93134
rect 78330 93218 78566 93454
rect 78330 92898 78566 93134
rect 109050 93218 109286 93454
rect 109050 92898 109286 93134
rect 139770 93218 140006 93454
rect 139770 92898 140006 93134
rect 170490 93218 170726 93454
rect 170490 92898 170726 93134
rect 201210 93218 201446 93454
rect 201210 92898 201446 93134
rect 231930 93218 232166 93454
rect 231930 92898 232166 93134
rect 262650 93218 262886 93454
rect 262650 92898 262886 93134
rect 293370 93218 293606 93454
rect 293370 92898 293606 93134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 32250 75218 32486 75454
rect 32250 74898 32486 75134
rect 62970 75218 63206 75454
rect 62970 74898 63206 75134
rect 93690 75218 93926 75454
rect 93690 74898 93926 75134
rect 124410 75218 124646 75454
rect 124410 74898 124646 75134
rect 155130 75218 155366 75454
rect 155130 74898 155366 75134
rect 185850 75218 186086 75454
rect 185850 74898 186086 75134
rect 216570 75218 216806 75454
rect 216570 74898 216806 75134
rect 247290 75218 247526 75454
rect 247290 74898 247526 75134
rect 278010 75218 278246 75454
rect 278010 74898 278246 75134
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 47610 57218 47846 57454
rect 47610 56898 47846 57134
rect 78330 57218 78566 57454
rect 78330 56898 78566 57134
rect 109050 57218 109286 57454
rect 109050 56898 109286 57134
rect 139770 57218 140006 57454
rect 139770 56898 140006 57134
rect 170490 57218 170726 57454
rect 170490 56898 170726 57134
rect 201210 57218 201446 57454
rect 201210 56898 201446 57134
rect 231930 57218 232166 57454
rect 231930 56898 232166 57134
rect 262650 57218 262886 57454
rect 262650 56898 262886 57134
rect 293370 57218 293606 57454
rect 293370 56898 293606 57134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 32250 39218 32486 39454
rect 32250 38898 32486 39134
rect 62970 39218 63206 39454
rect 62970 38898 63206 39134
rect 93690 39218 93926 39454
rect 93690 38898 93926 39134
rect 124410 39218 124646 39454
rect 124410 38898 124646 39134
rect 155130 39218 155366 39454
rect 155130 38898 155366 39134
rect 185850 39218 186086 39454
rect 185850 38898 186086 39134
rect 216570 39218 216806 39454
rect 216570 38898 216806 39134
rect 247290 39218 247526 39454
rect 247290 38898 247526 39134
rect 278010 39218 278246 39454
rect 278010 38898 278246 39134
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 394837 687218 395073 687454
rect 395157 687218 395393 687454
rect 395477 687218 395713 687454
rect 395797 687218 396033 687454
rect 396117 687218 396353 687454
rect 396437 687218 396673 687454
rect 396757 687218 396993 687454
rect 397077 687218 397313 687454
rect 397397 687218 397633 687454
rect 397717 687218 397953 687454
rect 394837 686898 395073 687134
rect 395157 686898 395393 687134
rect 395477 686898 395713 687134
rect 395797 686898 396033 687134
rect 396117 686898 396353 687134
rect 396437 686898 396673 687134
rect 396757 686898 396993 687134
rect 397077 686898 397313 687134
rect 397397 686898 397633 687134
rect 397717 686898 397953 687134
rect 461488 687218 461724 687454
rect 461808 687218 462044 687454
rect 462128 687218 462364 687454
rect 461488 686898 461724 687134
rect 461808 686898 462044 687134
rect 462128 686898 462364 687134
rect 538187 687218 538423 687454
rect 538507 687218 538743 687454
rect 538827 687218 539063 687454
rect 539147 687218 539383 687454
rect 539467 687218 539703 687454
rect 539787 687218 540023 687454
rect 540107 687218 540343 687454
rect 540427 687218 540663 687454
rect 540747 687218 540983 687454
rect 541067 687218 541303 687454
rect 541387 687218 541623 687454
rect 541707 687218 541943 687454
rect 542027 687218 542263 687454
rect 542347 687218 542583 687454
rect 542667 687218 542903 687454
rect 542987 687218 543223 687454
rect 543307 687218 543543 687454
rect 543627 687218 543863 687454
rect 543947 687218 544183 687454
rect 544267 687218 544503 687454
rect 544587 687218 544823 687454
rect 544907 687218 545143 687454
rect 545227 687218 545463 687454
rect 545547 687218 545783 687454
rect 545867 687218 546103 687454
rect 546187 687218 546423 687454
rect 546507 687218 546743 687454
rect 538187 686898 538423 687134
rect 538507 686898 538743 687134
rect 538827 686898 539063 687134
rect 539147 686898 539383 687134
rect 539467 686898 539703 687134
rect 539787 686898 540023 687134
rect 540107 686898 540343 687134
rect 540427 686898 540663 687134
rect 540747 686898 540983 687134
rect 541067 686898 541303 687134
rect 541387 686898 541623 687134
rect 541707 686898 541943 687134
rect 542027 686898 542263 687134
rect 542347 686898 542583 687134
rect 542667 686898 542903 687134
rect 542987 686898 543223 687134
rect 543307 686898 543543 687134
rect 543627 686898 543863 687134
rect 543947 686898 544183 687134
rect 544267 686898 544503 687134
rect 544587 686898 544823 687134
rect 544907 686898 545143 687134
rect 545227 686898 545463 687134
rect 545547 686898 545783 687134
rect 545867 686898 546103 687134
rect 546187 686898 546423 687134
rect 546507 686898 546743 687134
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 400049 669218 400285 669454
rect 400369 669218 400605 669454
rect 400689 669218 400925 669454
rect 401009 669218 401245 669454
rect 401329 669218 401565 669454
rect 401649 669218 401885 669454
rect 401969 669218 402205 669454
rect 402289 669218 402525 669454
rect 402609 669218 402845 669454
rect 402929 669218 403165 669454
rect 400049 668898 400285 669134
rect 400369 668898 400605 669134
rect 400689 668898 400925 669134
rect 401009 668898 401245 669134
rect 401329 668898 401565 669134
rect 401649 668898 401885 669134
rect 401969 668898 402205 669134
rect 402289 668898 402525 669134
rect 402609 668898 402845 669134
rect 402929 668898 403165 669134
rect 549345 669218 549581 669454
rect 549665 669218 549901 669454
rect 549985 669218 550221 669454
rect 550305 669218 550541 669454
rect 550625 669218 550861 669454
rect 550945 669218 551181 669454
rect 551265 669218 551501 669454
rect 551585 669218 551821 669454
rect 551905 669218 552141 669454
rect 552225 669218 552461 669454
rect 552545 669218 552781 669454
rect 552865 669218 553101 669454
rect 553185 669218 553421 669454
rect 553505 669218 553741 669454
rect 553825 669218 554061 669454
rect 554145 669218 554381 669454
rect 554465 669218 554701 669454
rect 554785 669218 555021 669454
rect 555105 669218 555341 669454
rect 555425 669218 555661 669454
rect 549345 668898 549581 669134
rect 549665 668898 549901 669134
rect 549985 668898 550221 669134
rect 550305 668898 550541 669134
rect 550625 668898 550861 669134
rect 550945 668898 551181 669134
rect 551265 668898 551501 669134
rect 551585 668898 551821 669134
rect 551905 668898 552141 669134
rect 552225 668898 552461 669134
rect 552545 668898 552781 669134
rect 552865 668898 553101 669134
rect 553185 668898 553421 669134
rect 553505 668898 553741 669134
rect 553825 668898 554061 669134
rect 554145 668898 554381 669134
rect 554465 668898 554701 669134
rect 554785 668898 555021 669134
rect 555105 668898 555341 669134
rect 555425 668898 555661 669134
rect 394837 651218 395073 651454
rect 395157 651218 395393 651454
rect 395477 651218 395713 651454
rect 395797 651218 396033 651454
rect 396117 651218 396353 651454
rect 396437 651218 396673 651454
rect 396757 651218 396993 651454
rect 397077 651218 397313 651454
rect 397397 651218 397633 651454
rect 397717 651218 397953 651454
rect 394837 650898 395073 651134
rect 395157 650898 395393 651134
rect 395477 650898 395713 651134
rect 395797 650898 396033 651134
rect 396117 650898 396353 651134
rect 396437 650898 396673 651134
rect 396757 650898 396993 651134
rect 397077 650898 397313 651134
rect 397397 650898 397633 651134
rect 397717 650898 397953 651134
rect 538187 651218 538423 651454
rect 538507 651218 538743 651454
rect 538827 651218 539063 651454
rect 539147 651218 539383 651454
rect 539467 651218 539703 651454
rect 539787 651218 540023 651454
rect 540107 651218 540343 651454
rect 540427 651218 540663 651454
rect 540747 651218 540983 651454
rect 541067 651218 541303 651454
rect 541387 651218 541623 651454
rect 541707 651218 541943 651454
rect 542027 651218 542263 651454
rect 542347 651218 542583 651454
rect 542667 651218 542903 651454
rect 542987 651218 543223 651454
rect 543307 651218 543543 651454
rect 543627 651218 543863 651454
rect 543947 651218 544183 651454
rect 544267 651218 544503 651454
rect 544587 651218 544823 651454
rect 544907 651218 545143 651454
rect 545227 651218 545463 651454
rect 545547 651218 545783 651454
rect 545867 651218 546103 651454
rect 546187 651218 546423 651454
rect 546507 651218 546743 651454
rect 538187 650898 538423 651134
rect 538507 650898 538743 651134
rect 538827 650898 539063 651134
rect 539147 650898 539383 651134
rect 539467 650898 539703 651134
rect 539787 650898 540023 651134
rect 540107 650898 540343 651134
rect 540427 650898 540663 651134
rect 540747 650898 540983 651134
rect 541067 650898 541303 651134
rect 541387 650898 541623 651134
rect 541707 650898 541943 651134
rect 542027 650898 542263 651134
rect 542347 650898 542583 651134
rect 542667 650898 542903 651134
rect 542987 650898 543223 651134
rect 543307 650898 543543 651134
rect 543627 650898 543863 651134
rect 543947 650898 544183 651134
rect 544267 650898 544503 651134
rect 544587 650898 544823 651134
rect 544907 650898 545143 651134
rect 545227 650898 545463 651134
rect 545547 650898 545783 651134
rect 545867 650898 546103 651134
rect 546187 650898 546423 651134
rect 546507 650898 546743 651134
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 400049 633218 400285 633454
rect 400369 633218 400605 633454
rect 400689 633218 400925 633454
rect 401009 633218 401245 633454
rect 401329 633218 401565 633454
rect 401649 633218 401885 633454
rect 401969 633218 402205 633454
rect 402289 633218 402525 633454
rect 402609 633218 402845 633454
rect 402929 633218 403165 633454
rect 400049 632898 400285 633134
rect 400369 632898 400605 633134
rect 400689 632898 400925 633134
rect 401009 632898 401245 633134
rect 401329 632898 401565 633134
rect 401649 632898 401885 633134
rect 401969 632898 402205 633134
rect 402289 632898 402525 633134
rect 402609 632898 402845 633134
rect 402929 632898 403165 633134
rect 461420 633218 461656 633454
rect 461420 632898 461656 633134
rect 473714 633218 473950 633454
rect 474034 633218 474270 633454
rect 474354 633218 474590 633454
rect 474674 633218 474910 633454
rect 474994 633218 475230 633454
rect 475314 633218 475550 633454
rect 473714 632898 473950 633134
rect 474034 632898 474270 633134
rect 474354 632898 474590 633134
rect 474674 632898 474910 633134
rect 474994 632898 475230 633134
rect 475314 632898 475550 633134
rect 486350 633218 486586 633454
rect 486670 633218 486906 633454
rect 486990 633218 487226 633454
rect 487310 633218 487546 633454
rect 487630 633218 487866 633454
rect 486350 632898 486586 633134
rect 486670 632898 486906 633134
rect 486990 632898 487226 633134
rect 487310 632898 487546 633134
rect 487630 632898 487866 633134
rect 549345 633218 549581 633454
rect 549665 633218 549901 633454
rect 549985 633218 550221 633454
rect 550305 633218 550541 633454
rect 550625 633218 550861 633454
rect 550945 633218 551181 633454
rect 551265 633218 551501 633454
rect 551585 633218 551821 633454
rect 551905 633218 552141 633454
rect 552225 633218 552461 633454
rect 552545 633218 552781 633454
rect 552865 633218 553101 633454
rect 553185 633218 553421 633454
rect 553505 633218 553741 633454
rect 553825 633218 554061 633454
rect 554145 633218 554381 633454
rect 554465 633218 554701 633454
rect 554785 633218 555021 633454
rect 555105 633218 555341 633454
rect 555425 633218 555661 633454
rect 549345 632898 549581 633134
rect 549665 632898 549901 633134
rect 549985 632898 550221 633134
rect 550305 632898 550541 633134
rect 550625 632898 550861 633134
rect 550945 632898 551181 633134
rect 551265 632898 551501 633134
rect 551585 632898 551821 633134
rect 551905 632898 552141 633134
rect 552225 632898 552461 633134
rect 552545 632898 552781 633134
rect 552865 632898 553101 633134
rect 553185 632898 553421 633134
rect 553505 632898 553741 633134
rect 553825 632898 554061 633134
rect 554145 632898 554381 633134
rect 554465 632898 554701 633134
rect 554785 632898 555021 633134
rect 555105 632898 555341 633134
rect 555425 632898 555661 633134
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 404916 561218 405152 561454
rect 404916 560898 405152 561134
rect 414847 561218 415083 561454
rect 414847 560898 415083 561134
rect 399951 543218 400187 543454
rect 399951 542898 400187 543134
rect 409881 543218 410117 543454
rect 409881 542898 410117 543134
rect 419812 543218 420048 543454
rect 419812 542898 420048 543134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 394837 687454
rect 395073 687218 395157 687454
rect 395393 687218 395477 687454
rect 395713 687218 395797 687454
rect 396033 687218 396117 687454
rect 396353 687218 396437 687454
rect 396673 687218 396757 687454
rect 396993 687218 397077 687454
rect 397313 687218 397397 687454
rect 397633 687218 397717 687454
rect 397953 687218 461488 687454
rect 461724 687218 461808 687454
rect 462044 687218 462128 687454
rect 462364 687218 538187 687454
rect 538423 687218 538507 687454
rect 538743 687218 538827 687454
rect 539063 687218 539147 687454
rect 539383 687218 539467 687454
rect 539703 687218 539787 687454
rect 540023 687218 540107 687454
rect 540343 687218 540427 687454
rect 540663 687218 540747 687454
rect 540983 687218 541067 687454
rect 541303 687218 541387 687454
rect 541623 687218 541707 687454
rect 541943 687218 542027 687454
rect 542263 687218 542347 687454
rect 542583 687218 542667 687454
rect 542903 687218 542987 687454
rect 543223 687218 543307 687454
rect 543543 687218 543627 687454
rect 543863 687218 543947 687454
rect 544183 687218 544267 687454
rect 544503 687218 544587 687454
rect 544823 687218 544907 687454
rect 545143 687218 545227 687454
rect 545463 687218 545547 687454
rect 545783 687218 545867 687454
rect 546103 687218 546187 687454
rect 546423 687218 546507 687454
rect 546743 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 394837 687134
rect 395073 686898 395157 687134
rect 395393 686898 395477 687134
rect 395713 686898 395797 687134
rect 396033 686898 396117 687134
rect 396353 686898 396437 687134
rect 396673 686898 396757 687134
rect 396993 686898 397077 687134
rect 397313 686898 397397 687134
rect 397633 686898 397717 687134
rect 397953 686898 461488 687134
rect 461724 686898 461808 687134
rect 462044 686898 462128 687134
rect 462364 686898 538187 687134
rect 538423 686898 538507 687134
rect 538743 686898 538827 687134
rect 539063 686898 539147 687134
rect 539383 686898 539467 687134
rect 539703 686898 539787 687134
rect 540023 686898 540107 687134
rect 540343 686898 540427 687134
rect 540663 686898 540747 687134
rect 540983 686898 541067 687134
rect 541303 686898 541387 687134
rect 541623 686898 541707 687134
rect 541943 686898 542027 687134
rect 542263 686898 542347 687134
rect 542583 686898 542667 687134
rect 542903 686898 542987 687134
rect 543223 686898 543307 687134
rect 543543 686898 543627 687134
rect 543863 686898 543947 687134
rect 544183 686898 544267 687134
rect 544503 686898 544587 687134
rect 544823 686898 544907 687134
rect 545143 686898 545227 687134
rect 545463 686898 545547 687134
rect 545783 686898 545867 687134
rect 546103 686898 546187 687134
rect 546423 686898 546507 687134
rect 546743 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 400049 669454
rect 400285 669218 400369 669454
rect 400605 669218 400689 669454
rect 400925 669218 401009 669454
rect 401245 669218 401329 669454
rect 401565 669218 401649 669454
rect 401885 669218 401969 669454
rect 402205 669218 402289 669454
rect 402525 669218 402609 669454
rect 402845 669218 402929 669454
rect 403165 669218 549345 669454
rect 549581 669218 549665 669454
rect 549901 669218 549985 669454
rect 550221 669218 550305 669454
rect 550541 669218 550625 669454
rect 550861 669218 550945 669454
rect 551181 669218 551265 669454
rect 551501 669218 551585 669454
rect 551821 669218 551905 669454
rect 552141 669218 552225 669454
rect 552461 669218 552545 669454
rect 552781 669218 552865 669454
rect 553101 669218 553185 669454
rect 553421 669218 553505 669454
rect 553741 669218 553825 669454
rect 554061 669218 554145 669454
rect 554381 669218 554465 669454
rect 554701 669218 554785 669454
rect 555021 669218 555105 669454
rect 555341 669218 555425 669454
rect 555661 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 400049 669134
rect 400285 668898 400369 669134
rect 400605 668898 400689 669134
rect 400925 668898 401009 669134
rect 401245 668898 401329 669134
rect 401565 668898 401649 669134
rect 401885 668898 401969 669134
rect 402205 668898 402289 669134
rect 402525 668898 402609 669134
rect 402845 668898 402929 669134
rect 403165 668898 549345 669134
rect 549581 668898 549665 669134
rect 549901 668898 549985 669134
rect 550221 668898 550305 669134
rect 550541 668898 550625 669134
rect 550861 668898 550945 669134
rect 551181 668898 551265 669134
rect 551501 668898 551585 669134
rect 551821 668898 551905 669134
rect 552141 668898 552225 669134
rect 552461 668898 552545 669134
rect 552781 668898 552865 669134
rect 553101 668898 553185 669134
rect 553421 668898 553505 669134
rect 553741 668898 553825 669134
rect 554061 668898 554145 669134
rect 554381 668898 554465 669134
rect 554701 668898 554785 669134
rect 555021 668898 555105 669134
rect 555341 668898 555425 669134
rect 555661 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 55470 651454
rect 55706 651218 55790 651454
rect 56026 651218 56110 651454
rect 56346 651218 56430 651454
rect 56666 651218 56750 651454
rect 56986 651218 57070 651454
rect 57306 651218 57390 651454
rect 57626 651218 57710 651454
rect 57946 651218 58030 651454
rect 58266 651218 58350 651454
rect 58586 651218 58670 651454
rect 58906 651218 58990 651454
rect 59226 651218 59310 651454
rect 59546 651218 59630 651454
rect 59866 651218 59950 651454
rect 60186 651218 60270 651454
rect 60506 651218 60590 651454
rect 60826 651218 60910 651454
rect 61146 651218 286929 651454
rect 287165 651218 287249 651454
rect 287485 651218 287569 651454
rect 287805 651218 287889 651454
rect 288125 651218 288209 651454
rect 288445 651218 288529 651454
rect 288765 651218 288849 651454
rect 289085 651218 289169 651454
rect 289405 651218 289489 651454
rect 289725 651218 289809 651454
rect 290045 651218 290129 651454
rect 290365 651218 290449 651454
rect 290685 651218 290769 651454
rect 291005 651218 291089 651454
rect 291325 651218 291409 651454
rect 291645 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 394837 651454
rect 395073 651218 395157 651454
rect 395393 651218 395477 651454
rect 395713 651218 395797 651454
rect 396033 651218 396117 651454
rect 396353 651218 396437 651454
rect 396673 651218 396757 651454
rect 396993 651218 397077 651454
rect 397313 651218 397397 651454
rect 397633 651218 397717 651454
rect 397953 651218 538187 651454
rect 538423 651218 538507 651454
rect 538743 651218 538827 651454
rect 539063 651218 539147 651454
rect 539383 651218 539467 651454
rect 539703 651218 539787 651454
rect 540023 651218 540107 651454
rect 540343 651218 540427 651454
rect 540663 651218 540747 651454
rect 540983 651218 541067 651454
rect 541303 651218 541387 651454
rect 541623 651218 541707 651454
rect 541943 651218 542027 651454
rect 542263 651218 542347 651454
rect 542583 651218 542667 651454
rect 542903 651218 542987 651454
rect 543223 651218 543307 651454
rect 543543 651218 543627 651454
rect 543863 651218 543947 651454
rect 544183 651218 544267 651454
rect 544503 651218 544587 651454
rect 544823 651218 544907 651454
rect 545143 651218 545227 651454
rect 545463 651218 545547 651454
rect 545783 651218 545867 651454
rect 546103 651218 546187 651454
rect 546423 651218 546507 651454
rect 546743 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 55470 651134
rect 55706 650898 55790 651134
rect 56026 650898 56110 651134
rect 56346 650898 56430 651134
rect 56666 650898 56750 651134
rect 56986 650898 57070 651134
rect 57306 650898 57390 651134
rect 57626 650898 57710 651134
rect 57946 650898 58030 651134
rect 58266 650898 58350 651134
rect 58586 650898 58670 651134
rect 58906 650898 58990 651134
rect 59226 650898 59310 651134
rect 59546 650898 59630 651134
rect 59866 650898 59950 651134
rect 60186 650898 60270 651134
rect 60506 650898 60590 651134
rect 60826 650898 60910 651134
rect 61146 650898 286929 651134
rect 287165 650898 287249 651134
rect 287485 650898 287569 651134
rect 287805 650898 287889 651134
rect 288125 650898 288209 651134
rect 288445 650898 288529 651134
rect 288765 650898 288849 651134
rect 289085 650898 289169 651134
rect 289405 650898 289489 651134
rect 289725 650898 289809 651134
rect 290045 650898 290129 651134
rect 290365 650898 290449 651134
rect 290685 650898 290769 651134
rect 291005 650898 291089 651134
rect 291325 650898 291409 651134
rect 291645 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 394837 651134
rect 395073 650898 395157 651134
rect 395393 650898 395477 651134
rect 395713 650898 395797 651134
rect 396033 650898 396117 651134
rect 396353 650898 396437 651134
rect 396673 650898 396757 651134
rect 396993 650898 397077 651134
rect 397313 650898 397397 651134
rect 397633 650898 397717 651134
rect 397953 650898 538187 651134
rect 538423 650898 538507 651134
rect 538743 650898 538827 651134
rect 539063 650898 539147 651134
rect 539383 650898 539467 651134
rect 539703 650898 539787 651134
rect 540023 650898 540107 651134
rect 540343 650898 540427 651134
rect 540663 650898 540747 651134
rect 540983 650898 541067 651134
rect 541303 650898 541387 651134
rect 541623 650898 541707 651134
rect 541943 650898 542027 651134
rect 542263 650898 542347 651134
rect 542583 650898 542667 651134
rect 542903 650898 542987 651134
rect 543223 650898 543307 651134
rect 543543 650898 543627 651134
rect 543863 650898 543947 651134
rect 544183 650898 544267 651134
rect 544503 650898 544587 651134
rect 544823 650898 544907 651134
rect 545143 650898 545227 651134
rect 545463 650898 545547 651134
rect 545783 650898 545867 651134
rect 546103 650898 546187 651134
rect 546423 650898 546507 651134
rect 546743 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 44959 633454
rect 45195 633218 45279 633454
rect 45515 633218 45599 633454
rect 45835 633218 45919 633454
rect 46155 633218 46239 633454
rect 46475 633218 46559 633454
rect 46795 633218 46879 633454
rect 47115 633218 47199 633454
rect 47435 633218 47519 633454
rect 47755 633218 47839 633454
rect 48075 633218 48159 633454
rect 48395 633218 48479 633454
rect 48715 633218 48799 633454
rect 49035 633218 49119 633454
rect 49355 633218 49439 633454
rect 49675 633218 49759 633454
rect 49995 633218 50079 633454
rect 50315 633218 50399 633454
rect 50635 633218 50719 633454
rect 50955 633218 51039 633454
rect 51275 633218 51359 633454
rect 51595 633218 51679 633454
rect 51915 633218 51999 633454
rect 52235 633218 295141 633454
rect 295377 633218 295461 633454
rect 295697 633218 295781 633454
rect 296017 633218 296101 633454
rect 296337 633218 296421 633454
rect 296657 633218 296741 633454
rect 296977 633218 297061 633454
rect 297297 633218 297381 633454
rect 297617 633218 297701 633454
rect 297937 633218 298021 633454
rect 298257 633218 298341 633454
rect 298577 633218 298661 633454
rect 298897 633218 298981 633454
rect 299217 633218 299301 633454
rect 299537 633218 299621 633454
rect 299857 633218 299941 633454
rect 300177 633218 300261 633454
rect 300497 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 400049 633454
rect 400285 633218 400369 633454
rect 400605 633218 400689 633454
rect 400925 633218 401009 633454
rect 401245 633218 401329 633454
rect 401565 633218 401649 633454
rect 401885 633218 401969 633454
rect 402205 633218 402289 633454
rect 402525 633218 402609 633454
rect 402845 633218 402929 633454
rect 403165 633218 461420 633454
rect 461656 633218 473714 633454
rect 473950 633218 474034 633454
rect 474270 633218 474354 633454
rect 474590 633218 474674 633454
rect 474910 633218 474994 633454
rect 475230 633218 475314 633454
rect 475550 633218 486350 633454
rect 486586 633218 486670 633454
rect 486906 633218 486990 633454
rect 487226 633218 487310 633454
rect 487546 633218 487630 633454
rect 487866 633218 549345 633454
rect 549581 633218 549665 633454
rect 549901 633218 549985 633454
rect 550221 633218 550305 633454
rect 550541 633218 550625 633454
rect 550861 633218 550945 633454
rect 551181 633218 551265 633454
rect 551501 633218 551585 633454
rect 551821 633218 551905 633454
rect 552141 633218 552225 633454
rect 552461 633218 552545 633454
rect 552781 633218 552865 633454
rect 553101 633218 553185 633454
rect 553421 633218 553505 633454
rect 553741 633218 553825 633454
rect 554061 633218 554145 633454
rect 554381 633218 554465 633454
rect 554701 633218 554785 633454
rect 555021 633218 555105 633454
rect 555341 633218 555425 633454
rect 555661 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 44959 633134
rect 45195 632898 45279 633134
rect 45515 632898 45599 633134
rect 45835 632898 45919 633134
rect 46155 632898 46239 633134
rect 46475 632898 46559 633134
rect 46795 632898 46879 633134
rect 47115 632898 47199 633134
rect 47435 632898 47519 633134
rect 47755 632898 47839 633134
rect 48075 632898 48159 633134
rect 48395 632898 48479 633134
rect 48715 632898 48799 633134
rect 49035 632898 49119 633134
rect 49355 632898 49439 633134
rect 49675 632898 49759 633134
rect 49995 632898 50079 633134
rect 50315 632898 50399 633134
rect 50635 632898 50719 633134
rect 50955 632898 51039 633134
rect 51275 632898 51359 633134
rect 51595 632898 51679 633134
rect 51915 632898 51999 633134
rect 52235 632898 295141 633134
rect 295377 632898 295461 633134
rect 295697 632898 295781 633134
rect 296017 632898 296101 633134
rect 296337 632898 296421 633134
rect 296657 632898 296741 633134
rect 296977 632898 297061 633134
rect 297297 632898 297381 633134
rect 297617 632898 297701 633134
rect 297937 632898 298021 633134
rect 298257 632898 298341 633134
rect 298577 632898 298661 633134
rect 298897 632898 298981 633134
rect 299217 632898 299301 633134
rect 299537 632898 299621 633134
rect 299857 632898 299941 633134
rect 300177 632898 300261 633134
rect 300497 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 400049 633134
rect 400285 632898 400369 633134
rect 400605 632898 400689 633134
rect 400925 632898 401009 633134
rect 401245 632898 401329 633134
rect 401565 632898 401649 633134
rect 401885 632898 401969 633134
rect 402205 632898 402289 633134
rect 402525 632898 402609 633134
rect 402845 632898 402929 633134
rect 403165 632898 461420 633134
rect 461656 632898 473714 633134
rect 473950 632898 474034 633134
rect 474270 632898 474354 633134
rect 474590 632898 474674 633134
rect 474910 632898 474994 633134
rect 475230 632898 475314 633134
rect 475550 632898 486350 633134
rect 486586 632898 486670 633134
rect 486906 632898 486990 633134
rect 487226 632898 487310 633134
rect 487546 632898 487630 633134
rect 487866 632898 549345 633134
rect 549581 632898 549665 633134
rect 549901 632898 549985 633134
rect 550221 632898 550305 633134
rect 550541 632898 550625 633134
rect 550861 632898 550945 633134
rect 551181 632898 551265 633134
rect 551501 632898 551585 633134
rect 551821 632898 551905 633134
rect 552141 632898 552225 633134
rect 552461 632898 552545 633134
rect 552781 632898 552865 633134
rect 553101 632898 553185 633134
rect 553421 632898 553505 633134
rect 553741 632898 553825 633134
rect 554061 632898 554145 633134
rect 554381 632898 554465 633134
rect 554701 632898 554785 633134
rect 555021 632898 555105 633134
rect 555341 632898 555425 633134
rect 555661 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 55470 615454
rect 55706 615218 55790 615454
rect 56026 615218 56110 615454
rect 56346 615218 56430 615454
rect 56666 615218 56750 615454
rect 56986 615218 57070 615454
rect 57306 615218 57390 615454
rect 57626 615218 57710 615454
rect 57946 615218 58030 615454
rect 58266 615218 58350 615454
rect 58586 615218 58670 615454
rect 58906 615218 58990 615454
rect 59226 615218 59310 615454
rect 59546 615218 59630 615454
rect 59866 615218 59950 615454
rect 60186 615218 60270 615454
rect 60506 615218 60590 615454
rect 60826 615218 60910 615454
rect 61146 615218 286929 615454
rect 287165 615218 287249 615454
rect 287485 615218 287569 615454
rect 287805 615218 287889 615454
rect 288125 615218 288209 615454
rect 288445 615218 288529 615454
rect 288765 615218 288849 615454
rect 289085 615218 289169 615454
rect 289405 615218 289489 615454
rect 289725 615218 289809 615454
rect 290045 615218 290129 615454
rect 290365 615218 290449 615454
rect 290685 615218 290769 615454
rect 291005 615218 291089 615454
rect 291325 615218 291409 615454
rect 291645 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 55470 615134
rect 55706 614898 55790 615134
rect 56026 614898 56110 615134
rect 56346 614898 56430 615134
rect 56666 614898 56750 615134
rect 56986 614898 57070 615134
rect 57306 614898 57390 615134
rect 57626 614898 57710 615134
rect 57946 614898 58030 615134
rect 58266 614898 58350 615134
rect 58586 614898 58670 615134
rect 58906 614898 58990 615134
rect 59226 614898 59310 615134
rect 59546 614898 59630 615134
rect 59866 614898 59950 615134
rect 60186 614898 60270 615134
rect 60506 614898 60590 615134
rect 60826 614898 60910 615134
rect 61146 614898 286929 615134
rect 287165 614898 287249 615134
rect 287485 614898 287569 615134
rect 287805 614898 287889 615134
rect 288125 614898 288209 615134
rect 288445 614898 288529 615134
rect 288765 614898 288849 615134
rect 289085 614898 289169 615134
rect 289405 614898 289489 615134
rect 289725 614898 289809 615134
rect 290045 614898 290129 615134
rect 290365 614898 290449 615134
rect 290685 614898 290769 615134
rect 291005 614898 291089 615134
rect 291325 614898 291409 615134
rect 291645 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 44959 597454
rect 45195 597218 45279 597454
rect 45515 597218 45599 597454
rect 45835 597218 45919 597454
rect 46155 597218 46239 597454
rect 46475 597218 46559 597454
rect 46795 597218 46879 597454
rect 47115 597218 47199 597454
rect 47435 597218 47519 597454
rect 47755 597218 47839 597454
rect 48075 597218 48159 597454
rect 48395 597218 48479 597454
rect 48715 597218 48799 597454
rect 49035 597218 49119 597454
rect 49355 597218 49439 597454
rect 49675 597218 49759 597454
rect 49995 597218 50079 597454
rect 50315 597218 50399 597454
rect 50635 597218 50719 597454
rect 50955 597218 51039 597454
rect 51275 597218 51359 597454
rect 51595 597218 51679 597454
rect 51915 597218 51999 597454
rect 52235 597218 295141 597454
rect 295377 597218 295461 597454
rect 295697 597218 295781 597454
rect 296017 597218 296101 597454
rect 296337 597218 296421 597454
rect 296657 597218 296741 597454
rect 296977 597218 297061 597454
rect 297297 597218 297381 597454
rect 297617 597218 297701 597454
rect 297937 597218 298021 597454
rect 298257 597218 298341 597454
rect 298577 597218 298661 597454
rect 298897 597218 298981 597454
rect 299217 597218 299301 597454
rect 299537 597218 299621 597454
rect 299857 597218 299941 597454
rect 300177 597218 300261 597454
rect 300497 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 44959 597134
rect 45195 596898 45279 597134
rect 45515 596898 45599 597134
rect 45835 596898 45919 597134
rect 46155 596898 46239 597134
rect 46475 596898 46559 597134
rect 46795 596898 46879 597134
rect 47115 596898 47199 597134
rect 47435 596898 47519 597134
rect 47755 596898 47839 597134
rect 48075 596898 48159 597134
rect 48395 596898 48479 597134
rect 48715 596898 48799 597134
rect 49035 596898 49119 597134
rect 49355 596898 49439 597134
rect 49675 596898 49759 597134
rect 49995 596898 50079 597134
rect 50315 596898 50399 597134
rect 50635 596898 50719 597134
rect 50955 596898 51039 597134
rect 51275 596898 51359 597134
rect 51595 596898 51679 597134
rect 51915 596898 51999 597134
rect 52235 596898 295141 597134
rect 295377 596898 295461 597134
rect 295697 596898 295781 597134
rect 296017 596898 296101 597134
rect 296337 596898 296421 597134
rect 296657 596898 296741 597134
rect 296977 596898 297061 597134
rect 297297 596898 297381 597134
rect 297617 596898 297701 597134
rect 297937 596898 298021 597134
rect 298257 596898 298341 597134
rect 298577 596898 298661 597134
rect 298897 596898 298981 597134
rect 299217 596898 299301 597134
rect 299537 596898 299621 597134
rect 299857 596898 299941 597134
rect 300177 596898 300261 597134
rect 300497 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 286929 579454
rect 287165 579218 287249 579454
rect 287485 579218 287569 579454
rect 287805 579218 287889 579454
rect 288125 579218 288209 579454
rect 288445 579218 288529 579454
rect 288765 579218 288849 579454
rect 289085 579218 289169 579454
rect 289405 579218 289489 579454
rect 289725 579218 289809 579454
rect 290045 579218 290129 579454
rect 290365 579218 290449 579454
rect 290685 579218 290769 579454
rect 291005 579218 291089 579454
rect 291325 579218 291409 579454
rect 291645 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 286929 579134
rect 287165 578898 287249 579134
rect 287485 578898 287569 579134
rect 287805 578898 287889 579134
rect 288125 578898 288209 579134
rect 288445 578898 288529 579134
rect 288765 578898 288849 579134
rect 289085 578898 289169 579134
rect 289405 578898 289489 579134
rect 289725 578898 289809 579134
rect 290045 578898 290129 579134
rect 290365 578898 290449 579134
rect 290685 578898 290769 579134
rect 291005 578898 291089 579134
rect 291325 578898 291409 579134
rect 291645 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 404916 561454
rect 405152 561218 414847 561454
rect 415083 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 404916 561134
rect 405152 560898 414847 561134
rect 415083 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 399951 543454
rect 400187 543218 409881 543454
rect 410117 543218 419812 543454
rect 420048 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 399951 543134
rect 400187 542898 409881 543134
rect 410117 542898 419812 543134
rect 420048 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 32250 291454
rect 32486 291218 62970 291454
rect 63206 291218 93690 291454
rect 93926 291218 124410 291454
rect 124646 291218 155130 291454
rect 155366 291218 185850 291454
rect 186086 291218 216570 291454
rect 216806 291218 247290 291454
rect 247526 291218 278010 291454
rect 278246 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 32250 291134
rect 32486 290898 62970 291134
rect 63206 290898 93690 291134
rect 93926 290898 124410 291134
rect 124646 290898 155130 291134
rect 155366 290898 185850 291134
rect 186086 290898 216570 291134
rect 216806 290898 247290 291134
rect 247526 290898 278010 291134
rect 278246 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 47610 273454
rect 47846 273218 78330 273454
rect 78566 273218 109050 273454
rect 109286 273218 139770 273454
rect 140006 273218 170490 273454
rect 170726 273218 201210 273454
rect 201446 273218 231930 273454
rect 232166 273218 262650 273454
rect 262886 273218 293370 273454
rect 293606 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 47610 273134
rect 47846 272898 78330 273134
rect 78566 272898 109050 273134
rect 109286 272898 139770 273134
rect 140006 272898 170490 273134
rect 170726 272898 201210 273134
rect 201446 272898 231930 273134
rect 232166 272898 262650 273134
rect 262886 272898 293370 273134
rect 293606 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 32250 255454
rect 32486 255218 62970 255454
rect 63206 255218 93690 255454
rect 93926 255218 124410 255454
rect 124646 255218 155130 255454
rect 155366 255218 185850 255454
rect 186086 255218 216570 255454
rect 216806 255218 247290 255454
rect 247526 255218 278010 255454
rect 278246 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 32250 255134
rect 32486 254898 62970 255134
rect 63206 254898 93690 255134
rect 93926 254898 124410 255134
rect 124646 254898 155130 255134
rect 155366 254898 185850 255134
rect 186086 254898 216570 255134
rect 216806 254898 247290 255134
rect 247526 254898 278010 255134
rect 278246 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 47610 237454
rect 47846 237218 78330 237454
rect 78566 237218 109050 237454
rect 109286 237218 139770 237454
rect 140006 237218 170490 237454
rect 170726 237218 201210 237454
rect 201446 237218 231930 237454
rect 232166 237218 262650 237454
rect 262886 237218 293370 237454
rect 293606 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 47610 237134
rect 47846 236898 78330 237134
rect 78566 236898 109050 237134
rect 109286 236898 139770 237134
rect 140006 236898 170490 237134
rect 170726 236898 201210 237134
rect 201446 236898 231930 237134
rect 232166 236898 262650 237134
rect 262886 236898 293370 237134
rect 293606 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 32250 219454
rect 32486 219218 62970 219454
rect 63206 219218 93690 219454
rect 93926 219218 124410 219454
rect 124646 219218 155130 219454
rect 155366 219218 185850 219454
rect 186086 219218 216570 219454
rect 216806 219218 247290 219454
rect 247526 219218 278010 219454
rect 278246 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 32250 219134
rect 32486 218898 62970 219134
rect 63206 218898 93690 219134
rect 93926 218898 124410 219134
rect 124646 218898 155130 219134
rect 155366 218898 185850 219134
rect 186086 218898 216570 219134
rect 216806 218898 247290 219134
rect 247526 218898 278010 219134
rect 278246 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 47610 201454
rect 47846 201218 78330 201454
rect 78566 201218 109050 201454
rect 109286 201218 139770 201454
rect 140006 201218 170490 201454
rect 170726 201218 201210 201454
rect 201446 201218 231930 201454
rect 232166 201218 262650 201454
rect 262886 201218 293370 201454
rect 293606 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 47610 201134
rect 47846 200898 78330 201134
rect 78566 200898 109050 201134
rect 109286 200898 139770 201134
rect 140006 200898 170490 201134
rect 170726 200898 201210 201134
rect 201446 200898 231930 201134
rect 232166 200898 262650 201134
rect 262886 200898 293370 201134
rect 293606 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 32250 183454
rect 32486 183218 62970 183454
rect 63206 183218 93690 183454
rect 93926 183218 124410 183454
rect 124646 183218 155130 183454
rect 155366 183218 185850 183454
rect 186086 183218 216570 183454
rect 216806 183218 247290 183454
rect 247526 183218 278010 183454
rect 278246 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 32250 183134
rect 32486 182898 62970 183134
rect 63206 182898 93690 183134
rect 93926 182898 124410 183134
rect 124646 182898 155130 183134
rect 155366 182898 185850 183134
rect 186086 182898 216570 183134
rect 216806 182898 247290 183134
rect 247526 182898 278010 183134
rect 278246 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 47610 165454
rect 47846 165218 78330 165454
rect 78566 165218 109050 165454
rect 109286 165218 139770 165454
rect 140006 165218 170490 165454
rect 170726 165218 201210 165454
rect 201446 165218 231930 165454
rect 232166 165218 262650 165454
rect 262886 165218 293370 165454
rect 293606 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 47610 165134
rect 47846 164898 78330 165134
rect 78566 164898 109050 165134
rect 109286 164898 139770 165134
rect 140006 164898 170490 165134
rect 170726 164898 201210 165134
rect 201446 164898 231930 165134
rect 232166 164898 262650 165134
rect 262886 164898 293370 165134
rect 293606 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 32250 147454
rect 32486 147218 62970 147454
rect 63206 147218 93690 147454
rect 93926 147218 124410 147454
rect 124646 147218 155130 147454
rect 155366 147218 185850 147454
rect 186086 147218 216570 147454
rect 216806 147218 247290 147454
rect 247526 147218 278010 147454
rect 278246 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 32250 147134
rect 32486 146898 62970 147134
rect 63206 146898 93690 147134
rect 93926 146898 124410 147134
rect 124646 146898 155130 147134
rect 155366 146898 185850 147134
rect 186086 146898 216570 147134
rect 216806 146898 247290 147134
rect 247526 146898 278010 147134
rect 278246 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 47610 129454
rect 47846 129218 78330 129454
rect 78566 129218 109050 129454
rect 109286 129218 139770 129454
rect 140006 129218 170490 129454
rect 170726 129218 201210 129454
rect 201446 129218 231930 129454
rect 232166 129218 262650 129454
rect 262886 129218 293370 129454
rect 293606 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 47610 129134
rect 47846 128898 78330 129134
rect 78566 128898 109050 129134
rect 109286 128898 139770 129134
rect 140006 128898 170490 129134
rect 170726 128898 201210 129134
rect 201446 128898 231930 129134
rect 232166 128898 262650 129134
rect 262886 128898 293370 129134
rect 293606 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 32250 111454
rect 32486 111218 62970 111454
rect 63206 111218 93690 111454
rect 93926 111218 124410 111454
rect 124646 111218 155130 111454
rect 155366 111218 185850 111454
rect 186086 111218 216570 111454
rect 216806 111218 247290 111454
rect 247526 111218 278010 111454
rect 278246 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 32250 111134
rect 32486 110898 62970 111134
rect 63206 110898 93690 111134
rect 93926 110898 124410 111134
rect 124646 110898 155130 111134
rect 155366 110898 185850 111134
rect 186086 110898 216570 111134
rect 216806 110898 247290 111134
rect 247526 110898 278010 111134
rect 278246 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 47610 93454
rect 47846 93218 78330 93454
rect 78566 93218 109050 93454
rect 109286 93218 139770 93454
rect 140006 93218 170490 93454
rect 170726 93218 201210 93454
rect 201446 93218 231930 93454
rect 232166 93218 262650 93454
rect 262886 93218 293370 93454
rect 293606 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 47610 93134
rect 47846 92898 78330 93134
rect 78566 92898 109050 93134
rect 109286 92898 139770 93134
rect 140006 92898 170490 93134
rect 170726 92898 201210 93134
rect 201446 92898 231930 93134
rect 232166 92898 262650 93134
rect 262886 92898 293370 93134
rect 293606 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 32250 75454
rect 32486 75218 62970 75454
rect 63206 75218 93690 75454
rect 93926 75218 124410 75454
rect 124646 75218 155130 75454
rect 155366 75218 185850 75454
rect 186086 75218 216570 75454
rect 216806 75218 247290 75454
rect 247526 75218 278010 75454
rect 278246 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 32250 75134
rect 32486 74898 62970 75134
rect 63206 74898 93690 75134
rect 93926 74898 124410 75134
rect 124646 74898 155130 75134
rect 155366 74898 185850 75134
rect 186086 74898 216570 75134
rect 216806 74898 247290 75134
rect 247526 74898 278010 75134
rect 278246 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 47610 57454
rect 47846 57218 78330 57454
rect 78566 57218 109050 57454
rect 109286 57218 139770 57454
rect 140006 57218 170490 57454
rect 170726 57218 201210 57454
rect 201446 57218 231930 57454
rect 232166 57218 262650 57454
rect 262886 57218 293370 57454
rect 293606 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 47610 57134
rect 47846 56898 78330 57134
rect 78566 56898 109050 57134
rect 109286 56898 139770 57134
rect 140006 56898 170490 57134
rect 170726 56898 201210 57134
rect 201446 56898 231930 57134
rect 232166 56898 262650 57134
rect 262886 56898 293370 57134
rect 293606 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 32250 39454
rect 32486 39218 62970 39454
rect 63206 39218 93690 39454
rect 93926 39218 124410 39454
rect 124646 39218 155130 39454
rect 155366 39218 185850 39454
rect 186086 39218 216570 39454
rect 216806 39218 247290 39454
rect 247526 39218 278010 39454
rect 278246 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 32250 39134
rect 32486 38898 62970 39134
rect 63206 38898 93690 39134
rect 93926 38898 124410 39134
rect 124646 38898 155130 39134
rect 155366 38898 185850 39134
rect 186086 38898 216570 39134
rect 216806 38898 247290 39134
rect 247526 38898 278010 39134
rect 278246 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use LVDT  temp3
timestamp 1638096800
transform 1 0 66022 0 1 579250
box -26022 -21250 234618 98114
use temp_digital  temp2
timestamp 1638096800
transform 1 0 394000 0 1 535600
box 0 0 32000 32000
use analog_macro  temp1
timestamp 1638096800
transform 1 0 401554 0 1 616054
box -7554 -8854 157400 79208
use user_proj_example  mprj
timestamp 1638096800
transform 1 0 28000 0 1 34000
box 289 0 274238 276712
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 533600 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 312712 38414 556000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 312712 74414 556000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 312712 110414 556000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 312712 146414 556000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 312712 182414 556000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 312712 218414 556000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 312712 254414 556000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 312712 290414 556000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 569600 398414 605200 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 605200 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 605200 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 605200 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 605200 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 679364 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 679364 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 679364 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 679364 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 679364 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 679364 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 679364 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 679364 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 697262 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 697262 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 697262 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 697262 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 697262 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 32000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 32000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 32000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 32000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 32000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 32000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 32000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 32000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 533600 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 312712 42134 556000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 312712 78134 556000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 312712 114134 556000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 312712 150134 556000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 312712 186134 556000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 312712 222134 556000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 312712 258134 556000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 312712 294134 556000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 569600 402134 605200 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 605200 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 605200 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 605200 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 605200 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 679364 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 679364 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 679364 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 679364 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 679364 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 679364 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 679364 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 679364 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 697262 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 697262 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 697262 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 697262 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 697262 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 32000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 32000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 32000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 32000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 32000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 32000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 32000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 32000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 533600 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 312712 45854 556000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 312712 81854 556000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 312712 117854 556000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 312712 153854 556000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 312712 189854 556000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 312712 225854 556000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 312712 261854 556000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 312712 297854 556000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 569600 405854 605200 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 605200 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 605200 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 605200 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 605200 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 679364 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 679364 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 679364 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 679364 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 679364 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 679364 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 679364 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 679364 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 697262 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 697262 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 697262 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 697262 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 697262 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 32000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 32000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 32000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 32000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 32000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 32000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 32000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 32000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 533600 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 312712 49574 556000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 312712 85574 556000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 312712 121574 556000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 312712 157574 556000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 312712 193574 556000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 312712 229574 556000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 312712 265574 556000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 312712 301574 556000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 569600 409574 605200 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 605200 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 605200 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 605200 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 605200 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 679364 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 679364 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 679364 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 679364 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 679364 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 679364 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 679364 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 679364 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 697262 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 697262 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 697262 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 697262 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 697262 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 32000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 32000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 32000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 32000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 32000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 32000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 32000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 32000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 533600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 312712 63854 556000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 312712 99854 556000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 312712 135854 556000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 312712 171854 556000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 312712 207854 556000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 312712 243854 556000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 312712 279854 556000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 569600 423854 605200 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 605200 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 605200 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 605200 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 312712 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 679364 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 679364 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 679364 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 679364 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 679364 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 679364 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 679364 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 697262 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 697262 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 697262 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 697262 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 32000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 32000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 32000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 32000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 32000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 32000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 32000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 32000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 533600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 312712 67574 556000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 312712 103574 556000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 312712 139574 556000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 312712 175574 556000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 312712 211574 556000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 312712 247574 556000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 312712 283574 556000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 569600 427574 605200 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 605200 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 605200 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 605200 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 312712 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 679364 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 679364 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 679364 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 679364 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 679364 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 679364 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 679364 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 697262 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 697262 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 697262 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 697262 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 32000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 32000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 32000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 32000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 32000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 32000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 32000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 533600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 312712 56414 556000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 312712 92414 556000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 312712 128414 556000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 312712 164414 556000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 312712 200414 556000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 312712 236414 556000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 312712 272414 556000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 569600 416414 605200 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 605200 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 605200 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 605200 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 605200 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 679364 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 679364 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 679364 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 679364 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 679364 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 679364 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 679364 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 697262 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 697262 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 697262 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 697262 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 697262 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 32000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 32000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 32000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 32000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 32000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 32000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 32000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 533600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 312712 60134 556000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 312712 96134 556000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 312712 132134 556000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 312712 168134 556000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 312712 204134 556000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 312712 240134 556000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 312712 276134 556000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 569600 420134 605200 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 605200 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 605200 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 605200 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 679364 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 679364 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 679364 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 679364 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 679364 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 679364 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 679364 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 697262 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 697262 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 697262 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 697262 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
