VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LVDT
  CLASS BLOCK ;
  FOREIGN LVDT ;
  ORIGIN 130.110 106.250 ;
  SIZE 1303.200 BY 596.820 ;
  PIN Iin
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 50.000000 ;
    ANTENNADIFFAREA 30.449999 ;
    PORT
      LAYER li1 ;
        RECT -96.070 354.130 -95.900 355.750 ;
        RECT -93.490 354.130 -93.320 355.750 ;
        RECT -90.910 354.130 -90.740 355.750 ;
        RECT -88.330 354.130 -88.160 355.750 ;
        RECT -85.750 354.130 -85.580 355.750 ;
        RECT -83.170 354.130 -83.000 355.750 ;
        RECT -80.590 354.130 -80.420 355.750 ;
        RECT -78.010 354.130 -77.840 355.750 ;
        RECT -75.430 354.130 -75.260 355.750 ;
        RECT -72.850 354.130 -72.680 355.750 ;
        RECT -51.130 353.915 -50.960 355.535 ;
        RECT -48.550 353.915 -48.380 355.535 ;
        RECT -45.970 353.915 -45.800 355.535 ;
        RECT -43.390 353.915 -43.220 355.535 ;
        RECT -40.810 353.915 -40.640 355.535 ;
        RECT -38.230 353.915 -38.060 355.535 ;
        RECT -35.650 353.915 -35.480 355.535 ;
        RECT -33.070 353.915 -32.900 355.535 ;
        RECT -30.490 353.915 -30.320 355.535 ;
        RECT -27.910 353.915 -27.740 355.535 ;
        RECT 866.030 320.450 866.200 320.870 ;
        RECT 866.030 318.980 866.200 319.400 ;
        RECT 866.030 317.510 866.200 317.930 ;
        RECT 866.030 316.040 866.200 316.460 ;
        RECT 866.030 314.570 866.200 314.990 ;
        RECT 865.150 313.520 865.740 314.150 ;
      LAYER mcon ;
        RECT -96.070 355.395 -95.900 355.565 ;
        RECT -96.070 355.035 -95.900 355.205 ;
        RECT -96.070 354.675 -95.900 354.845 ;
        RECT -96.070 354.315 -95.900 354.485 ;
        RECT -93.490 355.395 -93.320 355.565 ;
        RECT -93.490 355.035 -93.320 355.205 ;
        RECT -93.490 354.675 -93.320 354.845 ;
        RECT -93.490 354.315 -93.320 354.485 ;
        RECT -90.910 355.395 -90.740 355.565 ;
        RECT -90.910 355.035 -90.740 355.205 ;
        RECT -90.910 354.675 -90.740 354.845 ;
        RECT -90.910 354.315 -90.740 354.485 ;
        RECT -88.330 355.395 -88.160 355.565 ;
        RECT -88.330 355.035 -88.160 355.205 ;
        RECT -88.330 354.675 -88.160 354.845 ;
        RECT -88.330 354.315 -88.160 354.485 ;
        RECT -85.750 355.395 -85.580 355.565 ;
        RECT -85.750 355.035 -85.580 355.205 ;
        RECT -85.750 354.675 -85.580 354.845 ;
        RECT -85.750 354.315 -85.580 354.485 ;
        RECT -83.170 355.395 -83.000 355.565 ;
        RECT -83.170 355.035 -83.000 355.205 ;
        RECT -83.170 354.675 -83.000 354.845 ;
        RECT -83.170 354.315 -83.000 354.485 ;
        RECT -80.590 355.395 -80.420 355.565 ;
        RECT -80.590 355.035 -80.420 355.205 ;
        RECT -80.590 354.675 -80.420 354.845 ;
        RECT -80.590 354.315 -80.420 354.485 ;
        RECT -78.010 355.395 -77.840 355.565 ;
        RECT -78.010 355.035 -77.840 355.205 ;
        RECT -78.010 354.675 -77.840 354.845 ;
        RECT -78.010 354.315 -77.840 354.485 ;
        RECT -75.430 355.395 -75.260 355.565 ;
        RECT -75.430 355.035 -75.260 355.205 ;
        RECT -75.430 354.675 -75.260 354.845 ;
        RECT -75.430 354.315 -75.260 354.485 ;
        RECT -72.850 355.395 -72.680 355.565 ;
        RECT -72.850 355.035 -72.680 355.205 ;
        RECT -72.850 354.675 -72.680 354.845 ;
        RECT -72.850 354.315 -72.680 354.485 ;
        RECT -51.130 355.180 -50.960 355.350 ;
        RECT -51.130 354.820 -50.960 354.990 ;
        RECT -51.130 354.460 -50.960 354.630 ;
        RECT -51.130 354.100 -50.960 354.270 ;
        RECT -48.550 355.180 -48.380 355.350 ;
        RECT -48.550 354.820 -48.380 354.990 ;
        RECT -48.550 354.460 -48.380 354.630 ;
        RECT -48.550 354.100 -48.380 354.270 ;
        RECT -45.970 355.180 -45.800 355.350 ;
        RECT -45.970 354.820 -45.800 354.990 ;
        RECT -45.970 354.460 -45.800 354.630 ;
        RECT -45.970 354.100 -45.800 354.270 ;
        RECT -43.390 355.180 -43.220 355.350 ;
        RECT -43.390 354.820 -43.220 354.990 ;
        RECT -43.390 354.460 -43.220 354.630 ;
        RECT -43.390 354.100 -43.220 354.270 ;
        RECT -40.810 355.180 -40.640 355.350 ;
        RECT -40.810 354.820 -40.640 354.990 ;
        RECT -40.810 354.460 -40.640 354.630 ;
        RECT -40.810 354.100 -40.640 354.270 ;
        RECT -38.230 355.180 -38.060 355.350 ;
        RECT -38.230 354.820 -38.060 354.990 ;
        RECT -38.230 354.460 -38.060 354.630 ;
        RECT -38.230 354.100 -38.060 354.270 ;
        RECT -35.650 355.180 -35.480 355.350 ;
        RECT -35.650 354.820 -35.480 354.990 ;
        RECT -35.650 354.460 -35.480 354.630 ;
        RECT -35.650 354.100 -35.480 354.270 ;
        RECT -33.070 355.180 -32.900 355.350 ;
        RECT -33.070 354.820 -32.900 354.990 ;
        RECT -33.070 354.460 -32.900 354.630 ;
        RECT -33.070 354.100 -32.900 354.270 ;
        RECT -30.490 355.180 -30.320 355.350 ;
        RECT -30.490 354.820 -30.320 354.990 ;
        RECT -30.490 354.460 -30.320 354.630 ;
        RECT -30.490 354.100 -30.320 354.270 ;
        RECT -27.910 355.180 -27.740 355.350 ;
        RECT -27.910 354.820 -27.740 354.990 ;
        RECT -27.910 354.460 -27.740 354.630 ;
        RECT -27.910 354.100 -27.740 354.270 ;
        RECT 866.030 320.575 866.200 320.745 ;
        RECT 866.030 319.105 866.200 319.275 ;
        RECT 866.030 317.635 866.200 317.805 ;
        RECT 866.030 316.165 866.200 316.335 ;
        RECT 866.030 314.695 866.200 314.865 ;
        RECT 865.335 313.725 865.505 313.895 ;
      LAYER met1 ;
        RECT -75.475 356.850 -75.245 359.065 ;
        RECT -96.210 356.200 -72.210 356.850 ;
        RECT -96.105 355.730 -95.895 356.200 ;
        RECT -93.525 355.730 -93.315 356.200 ;
        RECT -90.955 355.730 -90.745 356.200 ;
        RECT -88.395 355.730 -88.185 356.200 ;
        RECT -85.755 355.730 -85.545 356.200 ;
        RECT -96.105 355.395 -95.870 355.730 ;
        RECT -93.525 355.435 -93.290 355.730 ;
        RECT -90.955 355.435 -90.710 355.730 ;
        RECT -96.100 354.150 -95.870 355.395 ;
        RECT -93.520 354.150 -93.290 355.435 ;
        RECT -90.940 354.150 -90.710 355.435 ;
        RECT -88.395 355.415 -88.130 355.730 ;
        RECT -88.360 354.150 -88.130 355.415 ;
        RECT -85.780 355.395 -85.545 355.730 ;
        RECT -83.215 355.730 -83.005 356.200 ;
        RECT -80.575 355.730 -80.365 356.200 ;
        RECT -78.025 355.730 -77.815 356.200 ;
        RECT -75.465 355.730 -75.255 356.200 ;
        RECT -72.845 355.730 -72.635 356.200 ;
        RECT -85.780 354.150 -85.550 355.395 ;
        RECT -83.215 355.365 -82.970 355.730 ;
        RECT -83.200 354.150 -82.970 355.365 ;
        RECT -80.620 355.265 -80.365 355.730 ;
        RECT -80.620 354.150 -80.390 355.265 ;
        RECT -78.040 354.150 -77.810 355.730 ;
        RECT -75.465 355.305 -75.230 355.730 ;
        RECT -75.460 354.150 -75.230 355.305 ;
        RECT -72.880 355.395 -72.635 355.730 ;
        RECT -72.880 354.150 -72.650 355.395 ;
        RECT -51.160 354.190 -50.930 355.515 ;
        RECT -51.165 353.280 -50.925 354.190 ;
        RECT -48.580 354.110 -48.350 355.515 ;
        RECT -46.000 354.130 -45.770 355.515 ;
        RECT -43.420 354.190 -43.190 355.515 ;
        RECT -48.605 353.935 -48.350 354.110 ;
        RECT -48.605 353.280 -48.365 353.935 ;
        RECT -46.005 353.280 -45.765 354.130 ;
        RECT -43.445 353.935 -43.190 354.190 ;
        RECT -40.840 354.150 -40.610 355.515 ;
        RECT -38.260 354.190 -38.030 355.515 ;
        RECT -40.865 353.935 -40.610 354.150 ;
        RECT -43.445 353.280 -43.205 353.935 ;
        RECT -40.865 353.280 -40.625 353.935 ;
        RECT -38.265 353.280 -38.025 354.190 ;
        RECT -35.680 354.170 -35.450 355.515 ;
        RECT -35.685 353.280 -35.445 354.170 ;
        RECT -33.100 354.110 -32.870 355.515 ;
        RECT -30.520 354.150 -30.290 355.515 ;
        RECT -33.105 353.280 -32.865 354.110 ;
        RECT -30.545 353.935 -30.290 354.150 ;
        RECT -27.940 354.130 -27.710 355.515 ;
        RECT -27.940 353.935 -27.655 354.130 ;
        RECT -30.545 353.280 -30.305 353.935 ;
        RECT -27.895 353.280 -27.655 353.935 ;
        RECT -51.270 352.640 -27.450 353.280 ;
        RECT -27.965 350.650 -27.655 352.640 ;
        RECT 866.000 320.630 866.230 320.850 ;
        RECT 866.000 314.930 866.270 320.630 ;
        RECT 863.580 313.850 864.360 314.230 ;
        RECT 865.150 314.030 865.740 314.150 ;
        RECT 865.970 314.030 866.320 314.930 ;
        RECT 865.150 313.920 866.320 314.030 ;
        RECT 865.150 313.850 866.260 313.920 ;
        RECT 863.580 313.790 866.260 313.850 ;
        RECT 863.580 313.620 865.740 313.790 ;
        RECT 863.580 313.380 864.360 313.620 ;
        RECT 865.150 313.520 865.740 313.620 ;
      LAYER via ;
        RECT -96.020 356.235 -72.400 356.815 ;
        RECT -51.170 352.670 -27.550 353.250 ;
        RECT 863.680 313.515 864.260 314.095 ;
      LAYER met2 ;
        RECT -97.420 356.900 -95.420 356.980 ;
        RECT -97.420 356.150 -60.790 356.900 ;
        RECT -97.420 356.140 -95.420 356.150 ;
        RECT -61.660 353.330 -60.900 356.150 ;
        RECT -61.660 352.590 -27.500 353.330 ;
        RECT -61.660 352.580 -46.950 352.590 ;
        RECT 863.630 313.330 864.310 314.280 ;
      LAYER via2 ;
        RECT -97.360 356.220 -95.480 356.900 ;
        RECT -51.100 352.820 -50.820 353.100 ;
        RECT -50.700 352.820 -50.420 353.100 ;
        RECT -50.300 352.820 -50.020 353.100 ;
        RECT -49.900 352.820 -49.620 353.100 ;
        RECT -49.500 352.820 -49.220 353.100 ;
        RECT -49.100 352.820 -48.820 353.100 ;
        RECT -48.700 352.820 -48.420 353.100 ;
        RECT -48.300 352.820 -48.020 353.100 ;
        RECT -47.900 352.820 -47.620 353.100 ;
        RECT -47.500 352.820 -47.220 353.100 ;
        RECT -47.100 352.820 -46.820 353.100 ;
        RECT -46.700 352.820 -46.420 353.100 ;
        RECT -46.300 352.820 -46.020 353.100 ;
        RECT -45.900 352.820 -45.620 353.100 ;
        RECT -45.500 352.820 -45.220 353.100 ;
        RECT -45.100 352.820 -44.820 353.100 ;
        RECT -44.700 352.820 -44.420 353.100 ;
        RECT -44.300 352.820 -44.020 353.100 ;
        RECT -43.900 352.820 -43.620 353.100 ;
        RECT -43.500 352.820 -43.220 353.100 ;
        RECT -43.100 352.820 -42.820 353.100 ;
        RECT -42.700 352.820 -42.420 353.100 ;
        RECT -42.300 352.820 -42.020 353.100 ;
        RECT -41.900 352.820 -41.620 353.100 ;
        RECT -41.500 352.820 -41.220 353.100 ;
        RECT -41.100 352.820 -40.820 353.100 ;
        RECT -40.700 352.820 -40.420 353.100 ;
        RECT -40.300 352.820 -40.020 353.100 ;
        RECT -39.900 352.820 -39.620 353.100 ;
        RECT -39.500 352.820 -39.220 353.100 ;
        RECT -39.100 352.820 -38.820 353.100 ;
        RECT -38.700 352.820 -38.420 353.100 ;
        RECT -38.300 352.820 -38.020 353.100 ;
        RECT -37.900 352.820 -37.620 353.100 ;
        RECT -37.500 352.820 -37.220 353.100 ;
        RECT -37.100 352.820 -36.820 353.100 ;
        RECT -36.700 352.820 -36.420 353.100 ;
        RECT -36.300 352.820 -36.020 353.100 ;
        RECT -35.900 352.820 -35.620 353.100 ;
        RECT -35.500 352.820 -35.220 353.100 ;
        RECT -35.100 352.820 -34.820 353.100 ;
        RECT -34.700 352.820 -34.420 353.100 ;
        RECT -34.300 352.820 -34.020 353.100 ;
        RECT -33.900 352.820 -33.620 353.100 ;
        RECT -33.500 352.820 -33.220 353.100 ;
        RECT -33.100 352.820 -32.820 353.100 ;
        RECT -32.700 352.820 -32.420 353.100 ;
        RECT -32.300 352.820 -32.020 353.100 ;
        RECT -31.900 352.820 -31.620 353.100 ;
        RECT -31.500 352.820 -31.220 353.100 ;
        RECT -31.100 352.820 -30.820 353.100 ;
        RECT -30.700 352.820 -30.420 353.100 ;
        RECT -30.300 352.820 -30.020 353.100 ;
        RECT -29.900 352.820 -29.620 353.100 ;
        RECT -29.500 352.820 -29.220 353.100 ;
        RECT -29.100 352.820 -28.820 353.100 ;
        RECT -28.700 352.820 -28.420 353.100 ;
        RECT -28.300 352.820 -28.020 353.100 ;
        RECT -27.900 352.820 -27.620 353.100 ;
        RECT 863.630 313.465 864.310 314.145 ;
      LAYER met3 ;
        RECT -130.110 356.955 -96.650 357.550 ;
        RECT -130.110 356.165 -95.370 356.955 ;
        RECT -130.110 355.100 -96.650 356.165 ;
        RECT -5.410 353.380 -1.220 356.550 ;
        RECT -28.390 353.305 -1.220 353.380 ;
        RECT -51.270 352.615 -1.220 353.305 ;
        RECT -28.390 352.570 -1.220 352.615 ;
        RECT -5.410 351.280 -1.220 352.570 ;
        RECT 710.390 313.820 712.520 314.360 ;
        RECT 863.580 313.820 864.360 314.255 ;
        RECT 710.390 313.730 748.990 313.820 ;
        RECT 777.350 313.760 795.380 313.810 ;
        RECT 812.240 313.800 830.270 313.810 ;
        RECT 847.380 313.800 864.360 313.820 ;
        RECT 812.240 313.760 864.360 313.800 ;
        RECT 760.020 313.730 864.360 313.760 ;
        RECT 710.390 313.410 864.360 313.730 ;
        RECT 710.390 313.360 847.880 313.410 ;
        RECT 710.390 313.310 778.050 313.360 ;
        RECT 794.480 313.310 812.510 313.360 ;
        RECT 829.850 313.350 847.880 313.360 ;
        RECT 863.580 313.355 864.360 313.410 ;
        RECT 710.390 313.280 766.000 313.310 ;
        RECT 710.390 313.220 748.990 313.280 ;
        RECT 710.390 312.650 712.520 313.220 ;
      LAYER via3 ;
        RECT -5.275 351.355 -1.355 356.475 ;
        RECT 710.495 312.745 712.415 314.265 ;
      LAYER met4 ;
        RECT -5.365 356.130 -1.265 356.555 ;
        RECT 545.930 356.130 561.860 356.230 ;
        RECT -5.365 352.420 561.860 356.130 ;
        RECT -5.365 352.400 545.770 352.420 ;
        RECT -5.365 351.275 -1.265 352.400 ;
        RECT 558.850 351.920 561.860 352.420 ;
        RECT 558.860 314.030 561.860 351.920 ;
        RECT 710.435 314.030 712.475 314.365 ;
        RECT 558.860 312.770 712.475 314.030 ;
        RECT 562.090 312.730 712.475 312.770 ;
        RECT 710.435 312.645 712.475 312.730 ;
    END
  END Iin
  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1836.000000 ;
    ANTENNADIFFAREA 485.750000 ;
    PORT
      LAYER li1 ;
        RECT 103.290 271.960 104.120 273.360 ;
        RECT 116.390 271.830 117.070 273.900 ;
        RECT -96.560 232.930 -96.390 234.550 ;
        RECT -93.980 232.930 -93.810 234.550 ;
        RECT -91.400 232.930 -91.230 234.550 ;
        RECT -88.820 232.930 -88.650 234.550 ;
        RECT -86.240 232.930 -86.070 234.550 ;
        RECT -83.660 232.930 -83.490 234.550 ;
        RECT -81.080 232.930 -80.910 234.550 ;
        RECT -78.500 232.930 -78.330 234.550 ;
        RECT -75.920 232.930 -75.750 234.550 ;
        RECT -73.340 232.930 -73.170 234.550 ;
        RECT -51.120 232.535 -50.950 234.155 ;
        RECT -48.540 232.535 -48.370 234.155 ;
        RECT -45.960 232.535 -45.790 234.155 ;
        RECT -43.380 232.535 -43.210 234.155 ;
        RECT -40.800 232.535 -40.630 234.155 ;
        RECT -38.220 232.535 -38.050 234.155 ;
        RECT -35.640 232.535 -35.470 234.155 ;
        RECT -33.060 232.535 -32.890 234.155 ;
        RECT -30.480 232.535 -30.310 234.155 ;
        RECT -27.900 232.535 -27.730 234.155 ;
        RECT 104.710 216.600 106.970 218.170 ;
        RECT 107.270 216.650 107.610 216.700 ;
        RECT 117.790 216.650 118.130 216.730 ;
        RECT 128.410 216.660 128.750 216.810 ;
        RECT 139.880 216.730 140.220 216.780 ;
        RECT 150.400 216.730 150.740 216.810 ;
        RECT 161.020 216.770 161.360 216.890 ;
        RECT 172.430 216.770 172.770 216.810 ;
        RECT 173.060 216.770 174.360 216.860 ;
        RECT 160.850 216.760 175.400 216.770 ;
        RECT 182.950 216.760 183.290 216.840 ;
        RECT 193.570 216.760 193.910 216.920 ;
        RECT 160.850 216.730 193.910 216.760 ;
        RECT 139.880 216.720 193.910 216.730 ;
        RECT 139.880 216.680 193.960 216.720 ;
        RECT 139.190 216.660 193.960 216.680 ;
        RECT 128.300 216.650 193.960 216.660 ;
        RECT 107.270 216.600 193.960 216.650 ;
        RECT 104.710 216.280 193.960 216.600 ;
        RECT 104.710 216.230 160.640 216.280 ;
        RECT 160.850 216.260 193.960 216.280 ;
        RECT 104.710 216.200 141.200 216.230 ;
        RECT 104.710 216.150 128.030 216.200 ;
        RECT 104.710 215.370 106.970 216.150 ;
        RECT 107.270 214.750 107.610 216.150 ;
        RECT 117.790 215.080 118.130 216.150 ;
        RECT 128.300 215.970 141.200 216.200 ;
        RECT 117.790 214.820 118.160 215.080 ;
        RECT 107.270 213.720 107.510 214.750 ;
        RECT 107.270 209.870 107.500 213.720 ;
        RECT 107.270 208.250 107.510 209.870 ;
        RECT 107.270 204.400 107.500 208.250 ;
        RECT 107.270 202.780 107.510 204.400 ;
        RECT 107.270 198.930 107.500 202.780 ;
        RECT 107.270 197.310 107.510 198.930 ;
        RECT 107.270 193.580 107.500 197.310 ;
        RECT 107.130 187.570 107.790 193.580 ;
        RECT 117.870 193.090 118.100 214.820 ;
        RECT 128.370 214.800 128.790 215.970 ;
        RECT 139.880 214.830 140.220 215.970 ;
        RECT 150.400 215.160 150.740 216.230 ;
        RECT 160.850 215.810 175.400 216.260 ;
        RECT 150.400 214.900 150.770 215.160 ;
        RECT 128.470 193.230 128.700 214.800 ;
        RECT 139.880 213.800 140.120 214.830 ;
        RECT 139.880 209.950 140.110 213.800 ;
        RECT 139.880 208.330 140.120 209.950 ;
        RECT 139.880 204.480 140.110 208.330 ;
        RECT 139.880 202.860 140.120 204.480 ;
        RECT 139.880 199.010 140.110 202.860 ;
        RECT 139.880 197.390 140.120 199.010 ;
        RECT 139.880 193.990 140.110 197.390 ;
        RECT 117.920 191.840 118.090 193.090 ;
        RECT 128.500 191.840 128.670 193.230 ;
        RECT 117.790 187.570 118.130 187.650 ;
        RECT 128.410 187.570 128.750 187.730 ;
        RECT 139.850 187.650 140.510 193.990 ;
        RECT 150.480 193.170 150.710 214.900 ;
        RECT 160.980 214.880 161.400 215.810 ;
        RECT 161.080 193.310 161.310 214.880 ;
        RECT 172.430 214.860 172.770 215.810 ;
        RECT 182.950 215.190 183.290 216.260 ;
        RECT 192.310 215.810 193.960 216.260 ;
        RECT 182.950 214.930 183.320 215.190 ;
        RECT 172.430 213.830 172.670 214.860 ;
        RECT 172.430 209.980 172.660 213.830 ;
        RECT 172.430 208.360 172.670 209.980 ;
        RECT 172.430 204.510 172.660 208.360 ;
        RECT 172.430 202.890 172.670 204.510 ;
        RECT 172.430 199.040 172.660 202.890 ;
        RECT 172.430 197.420 172.670 199.040 ;
        RECT 172.430 193.590 172.660 197.420 ;
        RECT 150.530 191.920 150.700 193.170 ;
        RECT 161.110 191.920 161.280 193.310 ;
        RECT 172.220 192.550 172.830 193.590 ;
        RECT 183.030 193.200 183.260 214.930 ;
        RECT 193.530 214.910 193.950 215.810 ;
        RECT 193.630 193.340 193.860 214.910 ;
        RECT 172.220 192.310 172.880 192.550 ;
        RECT 150.400 187.650 150.740 187.730 ;
        RECT 161.020 187.650 161.360 187.810 ;
        RECT 139.850 187.600 161.360 187.650 ;
        RECT 172.250 187.680 172.880 192.310 ;
        RECT 183.080 191.950 183.250 193.200 ;
        RECT 193.660 191.950 193.830 193.340 ;
        RECT 182.950 187.680 183.290 187.760 ;
        RECT 193.570 187.680 193.910 187.840 ;
        RECT 172.250 187.630 193.910 187.680 ;
        RECT 107.130 187.520 128.750 187.570 ;
        RECT 106.580 187.300 128.750 187.520 ;
        RECT 139.190 187.380 161.360 187.600 ;
        RECT 171.740 187.410 193.910 187.630 ;
        RECT 106.580 187.120 128.790 187.300 ;
        RECT 139.190 187.200 161.400 187.380 ;
        RECT 139.190 187.150 160.640 187.200 ;
        RECT 106.580 187.070 128.030 187.120 ;
        RECT 107.130 186.540 107.790 187.070 ;
        RECT 107.270 185.670 107.610 186.540 ;
        RECT 117.790 186.000 118.130 187.070 ;
        RECT 117.790 185.740 118.160 186.000 ;
        RECT 107.270 184.640 107.510 185.670 ;
        RECT 107.270 180.790 107.500 184.640 ;
        RECT 107.270 179.170 107.510 180.790 ;
        RECT 107.270 175.320 107.500 179.170 ;
        RECT 107.270 173.700 107.510 175.320 ;
        RECT 107.270 169.850 107.500 173.700 ;
        RECT 107.270 168.230 107.510 169.850 ;
        RECT 107.270 164.580 107.500 168.230 ;
        RECT 107.200 158.400 107.860 164.580 ;
        RECT 117.870 164.010 118.100 185.740 ;
        RECT 128.370 185.720 128.790 187.120 ;
        RECT 139.850 186.950 140.510 187.150 ;
        RECT 139.880 185.750 140.220 186.950 ;
        RECT 150.400 186.080 150.740 187.150 ;
        RECT 150.400 185.820 150.770 186.080 ;
        RECT 128.470 164.150 128.700 185.720 ;
        RECT 139.880 184.720 140.120 185.750 ;
        RECT 139.880 180.870 140.110 184.720 ;
        RECT 139.880 179.250 140.120 180.870 ;
        RECT 139.880 175.400 140.110 179.250 ;
        RECT 139.880 173.780 140.120 175.400 ;
        RECT 139.880 169.930 140.110 173.780 ;
        RECT 139.880 168.310 140.120 169.930 ;
        RECT 139.880 164.770 140.110 168.310 ;
        RECT 117.920 162.760 118.090 164.010 ;
        RECT 128.500 162.760 128.670 164.150 ;
        RECT 117.790 158.400 118.130 158.480 ;
        RECT 128.410 158.400 128.750 158.560 ;
        RECT 139.740 158.480 140.400 164.770 ;
        RECT 150.480 164.090 150.710 185.820 ;
        RECT 160.980 185.800 161.400 187.200 ;
        RECT 171.740 187.230 193.950 187.410 ;
        RECT 171.740 187.180 193.190 187.230 ;
        RECT 161.080 164.230 161.310 185.800 ;
        RECT 172.250 185.630 172.880 187.180 ;
        RECT 182.950 186.110 183.290 187.180 ;
        RECT 182.950 185.850 183.320 186.110 ;
        RECT 172.430 184.750 172.670 185.630 ;
        RECT 172.430 180.900 172.660 184.750 ;
        RECT 172.430 179.280 172.670 180.900 ;
        RECT 172.430 175.430 172.660 179.280 ;
        RECT 172.430 173.810 172.670 175.430 ;
        RECT 172.430 169.960 172.660 173.810 ;
        RECT 172.430 168.340 172.670 169.960 ;
        RECT 172.430 164.490 172.660 168.340 ;
        RECT 150.530 162.840 150.700 164.090 ;
        RECT 161.110 162.840 161.280 164.230 ;
        RECT 172.430 164.120 172.670 164.490 ;
        RECT 183.030 164.120 183.260 185.850 ;
        RECT 193.530 185.830 193.950 187.230 ;
        RECT 193.630 164.260 193.860 185.830 ;
        RECT 172.500 163.860 172.670 164.120 ;
        RECT 150.400 158.480 150.740 158.560 ;
        RECT 161.020 158.480 161.360 158.640 ;
        RECT 139.740 158.430 161.360 158.480 ;
        RECT 172.250 158.510 172.880 163.860 ;
        RECT 183.080 162.870 183.250 164.120 ;
        RECT 193.660 162.870 193.830 164.260 ;
        RECT 182.950 158.510 183.290 158.590 ;
        RECT 193.570 158.510 193.910 158.670 ;
        RECT 172.250 158.460 193.910 158.510 ;
        RECT 107.200 158.350 128.750 158.400 ;
        RECT 106.580 158.130 128.750 158.350 ;
        RECT 139.190 158.210 161.360 158.430 ;
        RECT 171.740 158.240 193.910 158.460 ;
        RECT 106.580 157.950 128.790 158.130 ;
        RECT 139.190 158.030 161.400 158.210 ;
        RECT 139.190 157.980 160.640 158.030 ;
        RECT 106.580 157.900 128.030 157.950 ;
        RECT 107.200 157.540 107.860 157.900 ;
        RECT 107.270 156.500 107.610 157.540 ;
        RECT 117.790 156.830 118.130 157.900 ;
        RECT 117.790 156.570 118.160 156.830 ;
        RECT 107.270 155.470 107.510 156.500 ;
        RECT 107.270 151.620 107.500 155.470 ;
        RECT 107.270 150.000 107.510 151.620 ;
        RECT 107.270 146.150 107.500 150.000 ;
        RECT 107.270 144.530 107.510 146.150 ;
        RECT 107.270 140.680 107.500 144.530 ;
        RECT 107.270 139.060 107.510 140.680 ;
        RECT 107.270 135.360 107.500 139.060 ;
        RECT 107.050 129.220 107.710 135.360 ;
        RECT 117.870 134.840 118.100 156.570 ;
        RECT 128.370 156.550 128.790 157.950 ;
        RECT 139.740 157.730 140.400 157.980 ;
        RECT 139.880 156.580 140.220 157.730 ;
        RECT 150.400 156.910 150.740 157.980 ;
        RECT 150.400 156.650 150.770 156.910 ;
        RECT 128.470 134.980 128.700 156.550 ;
        RECT 139.880 155.550 140.120 156.580 ;
        RECT 139.880 151.700 140.110 155.550 ;
        RECT 139.880 150.080 140.120 151.700 ;
        RECT 139.880 146.230 140.110 150.080 ;
        RECT 139.880 144.610 140.120 146.230 ;
        RECT 139.880 140.760 140.110 144.610 ;
        RECT 139.880 139.140 140.120 140.760 ;
        RECT 139.880 135.400 140.110 139.140 ;
        RECT 117.920 133.590 118.090 134.840 ;
        RECT 128.500 133.590 128.670 134.980 ;
        RECT 117.790 129.220 118.130 129.300 ;
        RECT 128.410 129.220 128.750 129.380 ;
        RECT 139.820 129.300 140.480 135.400 ;
        RECT 150.480 134.920 150.710 156.650 ;
        RECT 160.980 156.630 161.400 158.030 ;
        RECT 171.740 158.060 193.950 158.240 ;
        RECT 171.740 158.010 193.190 158.060 ;
        RECT 172.250 156.940 172.880 158.010 ;
        RECT 182.950 156.940 183.290 158.010 ;
        RECT 161.080 135.060 161.310 156.630 ;
        RECT 172.430 156.610 172.770 156.940 ;
        RECT 182.950 156.680 183.320 156.940 ;
        RECT 172.430 155.580 172.670 156.610 ;
        RECT 172.430 151.730 172.660 155.580 ;
        RECT 172.430 150.110 172.670 151.730 ;
        RECT 172.430 146.260 172.660 150.110 ;
        RECT 172.430 144.640 172.670 146.260 ;
        RECT 172.430 140.790 172.660 144.640 ;
        RECT 172.430 139.170 172.670 140.790 ;
        RECT 172.430 135.320 172.660 139.170 ;
        RECT 150.530 133.670 150.700 134.920 ;
        RECT 161.110 133.670 161.280 135.060 ;
        RECT 172.430 134.950 172.670 135.320 ;
        RECT 183.030 134.950 183.260 156.680 ;
        RECT 193.530 156.660 193.950 158.060 ;
        RECT 193.630 135.090 193.860 156.660 ;
        RECT 172.500 134.680 172.670 134.950 ;
        RECT 150.400 129.300 150.740 129.380 ;
        RECT 161.020 129.300 161.360 129.460 ;
        RECT 139.820 129.250 161.360 129.300 ;
        RECT 172.250 129.330 172.880 134.680 ;
        RECT 183.080 133.700 183.250 134.950 ;
        RECT 193.660 133.700 193.830 135.090 ;
        RECT 182.950 129.330 183.290 129.410 ;
        RECT 193.570 129.330 193.910 129.490 ;
        RECT 172.250 129.280 193.910 129.330 ;
        RECT 107.050 129.170 128.750 129.220 ;
        RECT 106.580 128.950 128.750 129.170 ;
        RECT 139.190 129.030 161.360 129.250 ;
        RECT 171.740 129.060 193.910 129.280 ;
        RECT 106.580 128.770 128.790 128.950 ;
        RECT 139.190 128.850 161.400 129.030 ;
        RECT 139.190 128.800 160.640 128.850 ;
        RECT 106.580 128.720 128.030 128.770 ;
        RECT 107.050 128.320 107.710 128.720 ;
        RECT 107.270 127.320 107.610 128.320 ;
        RECT 117.790 127.650 118.130 128.720 ;
        RECT 117.790 127.390 118.160 127.650 ;
        RECT 107.270 126.290 107.510 127.320 ;
        RECT 107.270 122.440 107.500 126.290 ;
        RECT 107.270 120.820 107.510 122.440 ;
        RECT 107.270 116.970 107.500 120.820 ;
        RECT 107.270 115.350 107.510 116.970 ;
        RECT 107.270 111.500 107.500 115.350 ;
        RECT 107.270 109.880 107.510 111.500 ;
        RECT 107.270 106.030 107.500 109.880 ;
        RECT 107.270 105.670 107.510 106.030 ;
        RECT 107.050 99.900 107.710 105.670 ;
        RECT 117.870 105.660 118.100 127.390 ;
        RECT 128.370 127.370 128.790 128.770 ;
        RECT 139.820 128.360 140.480 128.800 ;
        RECT 139.880 127.400 140.220 128.360 ;
        RECT 150.400 127.730 150.740 128.800 ;
        RECT 150.400 127.470 150.770 127.730 ;
        RECT 128.470 105.800 128.700 127.370 ;
        RECT 139.880 126.370 140.120 127.400 ;
        RECT 139.880 122.520 140.110 126.370 ;
        RECT 139.880 120.900 140.120 122.520 ;
        RECT 139.880 117.050 140.110 120.900 ;
        RECT 139.880 115.430 140.120 117.050 ;
        RECT 139.880 111.580 140.110 115.430 ;
        RECT 139.880 109.960 140.120 111.580 ;
        RECT 139.880 106.290 140.110 109.960 ;
        RECT 117.920 104.410 118.090 105.660 ;
        RECT 128.500 104.410 128.670 105.800 ;
        RECT 117.790 99.900 118.130 99.980 ;
        RECT 128.410 99.900 128.750 100.060 ;
        RECT 139.630 99.980 140.290 106.290 ;
        RECT 150.480 105.740 150.710 127.470 ;
        RECT 160.980 127.450 161.400 128.850 ;
        RECT 171.740 128.880 193.950 129.060 ;
        RECT 171.740 128.830 193.190 128.880 ;
        RECT 172.250 127.760 172.880 128.830 ;
        RECT 182.950 127.760 183.290 128.830 ;
        RECT 161.080 105.880 161.310 127.450 ;
        RECT 172.430 127.430 172.770 127.760 ;
        RECT 182.950 127.500 183.320 127.760 ;
        RECT 172.430 126.400 172.670 127.430 ;
        RECT 172.430 122.550 172.660 126.400 ;
        RECT 172.430 120.930 172.670 122.550 ;
        RECT 172.430 117.080 172.660 120.930 ;
        RECT 172.430 115.460 172.670 117.080 ;
        RECT 172.430 111.610 172.660 115.460 ;
        RECT 172.430 109.990 172.670 111.610 ;
        RECT 172.430 106.140 172.660 109.990 ;
        RECT 150.530 104.490 150.700 105.740 ;
        RECT 161.110 104.490 161.280 105.880 ;
        RECT 172.430 105.850 172.670 106.140 ;
        RECT 150.400 99.980 150.740 100.060 ;
        RECT 161.020 99.980 161.360 100.140 ;
        RECT 139.630 99.930 161.360 99.980 ;
        RECT 172.330 100.010 172.960 105.850 ;
        RECT 183.030 105.770 183.260 127.500 ;
        RECT 193.530 127.480 193.950 128.880 ;
        RECT 193.630 105.910 193.860 127.480 ;
        RECT 183.080 104.520 183.250 105.770 ;
        RECT 193.660 104.520 193.830 105.910 ;
        RECT 182.950 100.010 183.290 100.090 ;
        RECT 193.570 100.010 193.910 100.170 ;
        RECT 172.330 99.960 193.910 100.010 ;
        RECT 107.050 99.850 128.750 99.900 ;
        RECT 106.580 99.630 128.750 99.850 ;
        RECT 139.190 99.710 161.360 99.930 ;
        RECT 171.740 99.740 193.910 99.960 ;
        RECT 106.580 99.450 128.790 99.630 ;
        RECT 139.190 99.530 161.400 99.710 ;
        RECT 139.190 99.480 160.640 99.530 ;
        RECT 106.580 99.400 128.030 99.450 ;
        RECT 107.050 98.460 107.710 99.400 ;
        RECT 107.270 98.000 107.610 98.460 ;
        RECT 117.790 98.330 118.130 99.400 ;
        RECT 117.790 98.070 118.160 98.330 ;
        RECT 107.270 96.970 107.510 98.000 ;
        RECT 107.270 93.120 107.500 96.970 ;
        RECT 107.270 91.500 107.510 93.120 ;
        RECT 107.270 87.650 107.500 91.500 ;
        RECT 107.270 86.030 107.510 87.650 ;
        RECT 107.270 82.180 107.500 86.030 ;
        RECT 107.270 80.560 107.510 82.180 ;
        RECT 107.270 76.710 107.500 80.560 ;
        RECT 107.270 76.650 107.510 76.710 ;
        RECT 107.200 70.620 107.860 76.650 ;
        RECT 117.870 76.340 118.100 98.070 ;
        RECT 128.370 98.050 128.790 99.450 ;
        RECT 139.630 99.250 140.290 99.480 ;
        RECT 139.880 98.080 140.220 99.250 ;
        RECT 150.400 98.410 150.740 99.480 ;
        RECT 150.400 98.150 150.770 98.410 ;
        RECT 128.470 76.480 128.700 98.050 ;
        RECT 139.880 97.050 140.120 98.080 ;
        RECT 139.880 93.200 140.110 97.050 ;
        RECT 139.880 91.580 140.120 93.200 ;
        RECT 139.880 87.730 140.110 91.580 ;
        RECT 139.880 86.110 140.120 87.730 ;
        RECT 139.880 82.260 140.110 86.110 ;
        RECT 139.880 80.640 140.120 82.260 ;
        RECT 139.880 76.880 140.110 80.640 ;
        RECT 117.920 75.090 118.090 76.340 ;
        RECT 128.500 75.090 128.670 76.480 ;
        RECT 117.840 70.620 118.180 70.700 ;
        RECT 128.460 70.620 128.800 70.780 ;
        RECT 139.850 70.700 140.510 76.880 ;
        RECT 150.480 76.420 150.710 98.150 ;
        RECT 160.980 98.130 161.400 99.530 ;
        RECT 171.740 99.560 193.950 99.740 ;
        RECT 171.740 99.510 193.190 99.560 ;
        RECT 172.330 98.930 172.960 99.510 ;
        RECT 161.080 76.560 161.310 98.130 ;
        RECT 172.430 98.110 172.770 98.930 ;
        RECT 182.950 98.440 183.290 99.510 ;
        RECT 182.950 98.180 183.320 98.440 ;
        RECT 172.430 97.080 172.670 98.110 ;
        RECT 172.430 93.230 172.660 97.080 ;
        RECT 172.430 91.610 172.670 93.230 ;
        RECT 172.430 87.760 172.660 91.610 ;
        RECT 172.430 86.140 172.670 87.760 ;
        RECT 172.430 82.290 172.660 86.140 ;
        RECT 172.430 80.670 172.670 82.290 ;
        RECT 172.430 76.820 172.660 80.670 ;
        RECT 150.530 75.170 150.700 76.420 ;
        RECT 161.110 75.170 161.280 76.560 ;
        RECT 172.430 76.450 172.670 76.820 ;
        RECT 183.030 76.450 183.260 98.180 ;
        RECT 193.530 98.160 193.950 99.560 ;
        RECT 193.630 76.590 193.860 98.160 ;
        RECT 172.500 76.240 172.670 76.450 ;
        RECT 150.450 70.700 150.790 70.780 ;
        RECT 161.070 70.700 161.410 70.860 ;
        RECT 139.850 70.650 161.410 70.700 ;
        RECT 172.250 70.730 172.880 76.240 ;
        RECT 183.080 75.200 183.250 76.450 ;
        RECT 193.660 75.200 193.830 76.590 ;
        RECT 183.000 70.730 183.340 70.810 ;
        RECT 193.620 70.730 193.960 70.890 ;
        RECT 172.250 70.680 193.960 70.730 ;
        RECT 107.200 70.570 128.800 70.620 ;
        RECT 106.630 70.350 128.800 70.570 ;
        RECT 139.240 70.430 161.410 70.650 ;
        RECT 171.790 70.460 193.960 70.680 ;
        RECT 106.630 70.170 128.840 70.350 ;
        RECT 139.240 70.250 161.450 70.430 ;
        RECT 139.240 70.200 160.690 70.250 ;
        RECT 106.630 70.120 128.080 70.170 ;
        RECT 107.200 69.610 107.860 70.120 ;
        RECT 107.320 68.720 107.660 69.610 ;
        RECT 117.840 69.050 118.180 70.120 ;
        RECT 117.840 68.790 118.210 69.050 ;
        RECT 107.320 67.690 107.560 68.720 ;
        RECT 107.320 63.840 107.550 67.690 ;
        RECT 107.320 62.220 107.560 63.840 ;
        RECT 107.320 58.370 107.550 62.220 ;
        RECT 107.320 56.750 107.560 58.370 ;
        RECT 107.320 52.900 107.550 56.750 ;
        RECT 107.320 51.280 107.560 52.900 ;
        RECT 107.320 47.430 107.550 51.280 ;
        RECT 107.320 47.080 107.560 47.430 ;
        RECT 107.270 46.910 107.620 47.080 ;
        RECT 117.920 47.060 118.150 68.790 ;
        RECT 128.420 68.770 128.840 70.170 ;
        RECT 139.850 69.840 140.510 70.200 ;
        RECT 139.930 68.800 140.270 69.840 ;
        RECT 150.450 69.130 150.790 70.200 ;
        RECT 150.450 68.870 150.820 69.130 ;
        RECT 128.520 47.200 128.750 68.770 ;
        RECT 139.930 67.770 140.170 68.800 ;
        RECT 139.930 63.920 140.160 67.770 ;
        RECT 139.930 62.300 140.170 63.920 ;
        RECT 139.930 58.450 140.160 62.300 ;
        RECT 139.930 56.830 140.170 58.450 ;
        RECT 139.930 52.980 140.160 56.830 ;
        RECT 139.930 51.360 140.170 52.980 ;
        RECT 139.930 47.510 140.160 51.360 ;
        RECT 139.930 47.500 140.170 47.510 ;
        RECT 107.270 41.080 107.930 46.910 ;
        RECT 117.970 45.810 118.140 47.060 ;
        RECT 128.550 45.810 128.720 47.200 ;
        RECT 139.870 46.950 140.340 47.500 ;
        RECT 150.530 47.140 150.760 68.870 ;
        RECT 161.030 68.850 161.450 70.250 ;
        RECT 171.790 70.280 194.000 70.460 ;
        RECT 171.790 70.230 193.240 70.280 ;
        RECT 172.250 69.320 172.880 70.230 ;
        RECT 161.130 47.280 161.360 68.850 ;
        RECT 172.480 68.830 172.820 69.320 ;
        RECT 183.000 69.160 183.340 70.230 ;
        RECT 183.000 68.900 183.370 69.160 ;
        RECT 172.480 67.800 172.720 68.830 ;
        RECT 172.480 63.950 172.710 67.800 ;
        RECT 172.480 62.330 172.720 63.950 ;
        RECT 172.480 58.480 172.710 62.330 ;
        RECT 172.480 56.860 172.720 58.480 ;
        RECT 172.480 53.010 172.710 56.860 ;
        RECT 172.480 51.390 172.720 53.010 ;
        RECT 172.480 47.540 172.710 51.390 ;
        RECT 117.930 41.080 118.270 41.160 ;
        RECT 128.550 41.080 128.890 41.240 ;
        RECT 139.820 41.160 140.480 46.950 ;
        RECT 150.580 45.890 150.750 47.140 ;
        RECT 161.160 45.890 161.330 47.280 ;
        RECT 172.480 47.170 172.720 47.540 ;
        RECT 183.080 47.170 183.310 68.900 ;
        RECT 193.580 68.880 194.000 70.280 ;
        RECT 193.680 47.310 193.910 68.880 ;
        RECT 172.550 46.710 172.720 47.170 ;
        RECT 150.540 41.160 150.880 41.240 ;
        RECT 161.160 41.160 161.500 41.320 ;
        RECT 139.820 41.110 161.500 41.160 ;
        RECT 172.330 41.190 172.960 46.710 ;
        RECT 183.130 45.920 183.300 47.170 ;
        RECT 193.710 45.920 193.880 47.310 ;
        RECT 183.090 41.190 183.430 41.270 ;
        RECT 193.710 41.190 194.050 41.350 ;
        RECT 172.330 41.140 194.050 41.190 ;
        RECT 107.270 41.030 128.890 41.080 ;
        RECT 106.720 40.810 128.890 41.030 ;
        RECT 139.330 40.890 161.500 41.110 ;
        RECT 171.880 40.920 194.050 41.140 ;
        RECT 106.720 40.630 128.930 40.810 ;
        RECT 139.330 40.710 161.540 40.890 ;
        RECT 139.330 40.660 160.780 40.710 ;
        RECT 106.720 40.580 128.170 40.630 ;
        RECT 107.270 39.870 107.930 40.580 ;
        RECT 107.410 39.180 107.750 39.870 ;
        RECT 117.930 39.510 118.270 40.580 ;
        RECT 117.930 39.250 118.300 39.510 ;
        RECT 107.410 38.150 107.650 39.180 ;
        RECT 107.410 34.300 107.640 38.150 ;
        RECT 107.410 32.680 107.650 34.300 ;
        RECT 107.410 28.830 107.640 32.680 ;
        RECT 107.410 27.210 107.650 28.830 ;
        RECT 107.410 23.360 107.640 27.210 ;
        RECT 107.410 21.740 107.650 23.360 ;
        RECT 107.410 17.890 107.640 21.740 ;
        RECT 107.410 17.520 107.650 17.890 ;
        RECT 118.010 17.520 118.240 39.250 ;
        RECT 128.510 39.230 128.930 40.630 ;
        RECT 139.820 39.910 140.480 40.660 ;
        RECT 140.020 39.260 140.360 39.910 ;
        RECT 150.540 39.590 150.880 40.660 ;
        RECT 150.540 39.330 150.910 39.590 ;
        RECT 128.610 17.660 128.840 39.230 ;
        RECT 140.020 38.230 140.260 39.260 ;
        RECT 140.020 34.380 140.250 38.230 ;
        RECT 140.020 32.760 140.260 34.380 ;
        RECT 140.020 28.910 140.250 32.760 ;
        RECT 140.020 27.290 140.260 28.910 ;
        RECT 140.020 23.440 140.250 27.290 ;
        RECT 140.020 21.820 140.260 23.440 ;
        RECT 140.020 17.970 140.250 21.820 ;
        RECT 107.480 16.270 107.650 17.520 ;
        RECT 118.060 16.270 118.230 17.520 ;
        RECT 128.640 16.270 128.810 17.660 ;
        RECT 140.020 17.600 140.260 17.970 ;
        RECT 150.620 17.600 150.850 39.330 ;
        RECT 161.120 39.310 161.540 40.710 ;
        RECT 171.880 40.740 194.090 40.920 ;
        RECT 171.880 40.690 193.330 40.740 ;
        RECT 172.330 39.790 172.960 40.690 ;
        RECT 161.220 17.740 161.450 39.310 ;
        RECT 172.570 39.290 172.910 39.790 ;
        RECT 183.090 39.620 183.430 40.690 ;
        RECT 183.090 39.360 183.460 39.620 ;
        RECT 172.570 38.260 172.810 39.290 ;
        RECT 172.570 34.410 172.800 38.260 ;
        RECT 172.570 32.790 172.810 34.410 ;
        RECT 172.570 28.940 172.800 32.790 ;
        RECT 172.570 27.320 172.810 28.940 ;
        RECT 172.570 23.470 172.800 27.320 ;
        RECT 172.570 21.850 172.810 23.470 ;
        RECT 172.570 18.000 172.800 21.850 ;
        RECT 140.090 16.350 140.260 17.600 ;
        RECT 150.670 16.350 150.840 17.600 ;
        RECT 161.250 16.350 161.420 17.740 ;
        RECT 172.570 17.630 172.810 18.000 ;
        RECT 183.170 17.630 183.400 39.360 ;
        RECT 193.670 39.340 194.090 40.740 ;
        RECT 193.770 17.770 194.000 39.340 ;
        RECT 172.640 16.380 172.810 17.630 ;
        RECT 183.220 16.380 183.390 17.630 ;
        RECT 193.800 16.380 193.970 17.770 ;
      LAYER mcon ;
        RECT 116.640 273.385 116.810 273.555 ;
        RECT 103.565 272.795 103.735 272.965 ;
        RECT 103.565 272.435 103.735 272.605 ;
        RECT 116.640 273.025 116.810 273.195 ;
        RECT 116.640 272.665 116.810 272.835 ;
        RECT 116.640 272.305 116.810 272.475 ;
        RECT -96.560 234.195 -96.390 234.365 ;
        RECT -96.560 233.835 -96.390 234.005 ;
        RECT -96.560 233.475 -96.390 233.645 ;
        RECT -96.560 233.115 -96.390 233.285 ;
        RECT -93.980 234.195 -93.810 234.365 ;
        RECT -93.980 233.835 -93.810 234.005 ;
        RECT -93.980 233.475 -93.810 233.645 ;
        RECT -93.980 233.115 -93.810 233.285 ;
        RECT -91.400 234.195 -91.230 234.365 ;
        RECT -91.400 233.835 -91.230 234.005 ;
        RECT -91.400 233.475 -91.230 233.645 ;
        RECT -91.400 233.115 -91.230 233.285 ;
        RECT -88.820 234.195 -88.650 234.365 ;
        RECT -88.820 233.835 -88.650 234.005 ;
        RECT -88.820 233.475 -88.650 233.645 ;
        RECT -88.820 233.115 -88.650 233.285 ;
        RECT -86.240 234.195 -86.070 234.365 ;
        RECT -86.240 233.835 -86.070 234.005 ;
        RECT -86.240 233.475 -86.070 233.645 ;
        RECT -86.240 233.115 -86.070 233.285 ;
        RECT -83.660 234.195 -83.490 234.365 ;
        RECT -83.660 233.835 -83.490 234.005 ;
        RECT -83.660 233.475 -83.490 233.645 ;
        RECT -83.660 233.115 -83.490 233.285 ;
        RECT -81.080 234.195 -80.910 234.365 ;
        RECT -81.080 233.835 -80.910 234.005 ;
        RECT -81.080 233.475 -80.910 233.645 ;
        RECT -81.080 233.115 -80.910 233.285 ;
        RECT -78.500 234.195 -78.330 234.365 ;
        RECT -78.500 233.835 -78.330 234.005 ;
        RECT -78.500 233.475 -78.330 233.645 ;
        RECT -78.500 233.115 -78.330 233.285 ;
        RECT -75.920 234.195 -75.750 234.365 ;
        RECT -75.920 233.835 -75.750 234.005 ;
        RECT -75.920 233.475 -75.750 233.645 ;
        RECT -75.920 233.115 -75.750 233.285 ;
        RECT -73.340 234.195 -73.170 234.365 ;
        RECT -73.340 233.835 -73.170 234.005 ;
        RECT -73.340 233.475 -73.170 233.645 ;
        RECT -73.340 233.115 -73.170 233.285 ;
        RECT -51.120 233.800 -50.950 233.970 ;
        RECT -51.120 233.440 -50.950 233.610 ;
        RECT -51.120 233.080 -50.950 233.250 ;
        RECT -51.120 232.720 -50.950 232.890 ;
        RECT -48.540 233.800 -48.370 233.970 ;
        RECT -48.540 233.440 -48.370 233.610 ;
        RECT -48.540 233.080 -48.370 233.250 ;
        RECT -48.540 232.720 -48.370 232.890 ;
        RECT -45.960 233.800 -45.790 233.970 ;
        RECT -45.960 233.440 -45.790 233.610 ;
        RECT -45.960 233.080 -45.790 233.250 ;
        RECT -45.960 232.720 -45.790 232.890 ;
        RECT -43.380 233.800 -43.210 233.970 ;
        RECT -43.380 233.440 -43.210 233.610 ;
        RECT -43.380 233.080 -43.210 233.250 ;
        RECT -43.380 232.720 -43.210 232.890 ;
        RECT -40.800 233.800 -40.630 233.970 ;
        RECT -40.800 233.440 -40.630 233.610 ;
        RECT -40.800 233.080 -40.630 233.250 ;
        RECT -40.800 232.720 -40.630 232.890 ;
        RECT -38.220 233.800 -38.050 233.970 ;
        RECT -38.220 233.440 -38.050 233.610 ;
        RECT -38.220 233.080 -38.050 233.250 ;
        RECT -38.220 232.720 -38.050 232.890 ;
        RECT -35.640 233.800 -35.470 233.970 ;
        RECT -35.640 233.440 -35.470 233.610 ;
        RECT -35.640 233.080 -35.470 233.250 ;
        RECT -35.640 232.720 -35.470 232.890 ;
        RECT -33.060 233.800 -32.890 233.970 ;
        RECT -33.060 233.440 -32.890 233.610 ;
        RECT -33.060 233.080 -32.890 233.250 ;
        RECT -33.060 232.720 -32.890 232.890 ;
        RECT -30.480 233.800 -30.310 233.970 ;
        RECT -30.480 233.440 -30.310 233.610 ;
        RECT -30.480 233.080 -30.310 233.250 ;
        RECT -30.480 232.720 -30.310 232.890 ;
        RECT -27.900 233.800 -27.730 233.970 ;
        RECT -27.900 233.440 -27.730 233.610 ;
        RECT -27.900 233.080 -27.730 233.250 ;
        RECT -27.900 232.720 -27.730 232.890 ;
        RECT 107.340 214.985 107.510 215.155 ;
        RECT 117.920 214.985 118.090 215.155 ;
        RECT 128.500 214.985 128.670 215.155 ;
        RECT 107.340 214.625 107.510 214.795 ;
        RECT 139.950 215.065 140.120 215.235 ;
        RECT 150.530 215.065 150.700 215.235 ;
        RECT 161.110 215.065 161.280 215.235 ;
        RECT 107.340 214.265 107.510 214.435 ;
        RECT 107.340 213.905 107.510 214.075 ;
        RECT 117.920 214.625 118.090 214.795 ;
        RECT 117.920 214.265 118.090 214.435 ;
        RECT 117.920 213.905 118.090 214.075 ;
        RECT 107.340 209.515 107.510 209.685 ;
        RECT 107.340 209.155 107.510 209.325 ;
        RECT 107.340 208.795 107.510 208.965 ;
        RECT 107.340 208.435 107.510 208.605 ;
        RECT 117.920 209.515 118.090 209.685 ;
        RECT 117.920 209.155 118.090 209.325 ;
        RECT 117.920 208.795 118.090 208.965 ;
        RECT 117.920 208.435 118.090 208.605 ;
        RECT 107.340 204.045 107.510 204.215 ;
        RECT 107.340 203.685 107.510 203.855 ;
        RECT 107.340 203.325 107.510 203.495 ;
        RECT 107.340 202.965 107.510 203.135 ;
        RECT 117.920 204.045 118.090 204.215 ;
        RECT 117.920 203.685 118.090 203.855 ;
        RECT 117.920 203.325 118.090 203.495 ;
        RECT 117.920 202.965 118.090 203.135 ;
        RECT 107.340 198.575 107.510 198.745 ;
        RECT 107.340 198.215 107.510 198.385 ;
        RECT 107.340 197.855 107.510 198.025 ;
        RECT 107.340 197.495 107.510 197.665 ;
        RECT 117.920 198.575 118.090 198.745 ;
        RECT 117.920 198.215 118.090 198.385 ;
        RECT 117.920 197.855 118.090 198.025 ;
        RECT 117.920 197.495 118.090 197.665 ;
        RECT 107.340 193.105 107.510 193.275 ;
        RECT 117.920 193.105 118.090 193.275 ;
        RECT 128.500 214.625 128.670 214.795 ;
        RECT 128.500 214.265 128.670 214.435 ;
        RECT 128.500 213.905 128.670 214.075 ;
        RECT 128.500 209.515 128.670 209.685 ;
        RECT 128.500 209.155 128.670 209.325 ;
        RECT 128.500 208.795 128.670 208.965 ;
        RECT 128.500 208.435 128.670 208.605 ;
        RECT 128.500 204.045 128.670 204.215 ;
        RECT 128.500 203.685 128.670 203.855 ;
        RECT 128.500 203.325 128.670 203.495 ;
        RECT 128.500 202.965 128.670 203.135 ;
        RECT 128.500 198.575 128.670 198.745 ;
        RECT 128.500 198.215 128.670 198.385 ;
        RECT 128.500 197.855 128.670 198.025 ;
        RECT 128.500 197.495 128.670 197.665 ;
        RECT 139.950 214.705 140.120 214.875 ;
        RECT 172.500 215.095 172.670 215.265 ;
        RECT 183.080 215.095 183.250 215.265 ;
        RECT 193.660 215.095 193.830 215.265 ;
        RECT 139.950 214.345 140.120 214.515 ;
        RECT 139.950 213.985 140.120 214.155 ;
        RECT 150.530 214.705 150.700 214.875 ;
        RECT 150.530 214.345 150.700 214.515 ;
        RECT 150.530 213.985 150.700 214.155 ;
        RECT 139.950 209.595 140.120 209.765 ;
        RECT 139.950 209.235 140.120 209.405 ;
        RECT 139.950 208.875 140.120 209.045 ;
        RECT 139.950 208.515 140.120 208.685 ;
        RECT 150.530 209.595 150.700 209.765 ;
        RECT 150.530 209.235 150.700 209.405 ;
        RECT 150.530 208.875 150.700 209.045 ;
        RECT 150.530 208.515 150.700 208.685 ;
        RECT 139.950 204.125 140.120 204.295 ;
        RECT 139.950 203.765 140.120 203.935 ;
        RECT 139.950 203.405 140.120 203.575 ;
        RECT 139.950 203.045 140.120 203.215 ;
        RECT 150.530 204.125 150.700 204.295 ;
        RECT 150.530 203.765 150.700 203.935 ;
        RECT 150.530 203.405 150.700 203.575 ;
        RECT 150.530 203.045 150.700 203.215 ;
        RECT 139.950 198.655 140.120 198.825 ;
        RECT 139.950 198.295 140.120 198.465 ;
        RECT 139.950 197.935 140.120 198.105 ;
        RECT 139.950 197.575 140.120 197.745 ;
        RECT 150.530 198.655 150.700 198.825 ;
        RECT 150.530 198.295 150.700 198.465 ;
        RECT 150.530 197.935 150.700 198.105 ;
        RECT 150.530 197.575 150.700 197.745 ;
        RECT 128.500 193.105 128.670 193.275 ;
        RECT 107.340 192.745 107.510 192.915 ;
        RECT 107.340 192.385 107.510 192.555 ;
        RECT 107.340 192.025 107.510 192.195 ;
        RECT 117.920 192.745 118.090 192.915 ;
        RECT 117.920 192.385 118.090 192.555 ;
        RECT 117.920 192.025 118.090 192.195 ;
        RECT 128.500 192.745 128.670 192.915 ;
        RECT 128.500 192.385 128.670 192.555 ;
        RECT 128.500 192.025 128.670 192.195 ;
        RECT 139.950 193.185 140.120 193.355 ;
        RECT 150.530 193.185 150.700 193.355 ;
        RECT 161.110 214.705 161.280 214.875 ;
        RECT 161.110 214.345 161.280 214.515 ;
        RECT 161.110 213.985 161.280 214.155 ;
        RECT 161.110 209.595 161.280 209.765 ;
        RECT 161.110 209.235 161.280 209.405 ;
        RECT 161.110 208.875 161.280 209.045 ;
        RECT 161.110 208.515 161.280 208.685 ;
        RECT 161.110 204.125 161.280 204.295 ;
        RECT 161.110 203.765 161.280 203.935 ;
        RECT 161.110 203.405 161.280 203.575 ;
        RECT 161.110 203.045 161.280 203.215 ;
        RECT 161.110 198.655 161.280 198.825 ;
        RECT 161.110 198.295 161.280 198.465 ;
        RECT 161.110 197.935 161.280 198.105 ;
        RECT 161.110 197.575 161.280 197.745 ;
        RECT 172.500 214.735 172.670 214.905 ;
        RECT 172.500 214.375 172.670 214.545 ;
        RECT 172.500 214.015 172.670 214.185 ;
        RECT 183.080 214.735 183.250 214.905 ;
        RECT 183.080 214.375 183.250 214.545 ;
        RECT 183.080 214.015 183.250 214.185 ;
        RECT 172.500 209.625 172.670 209.795 ;
        RECT 172.500 209.265 172.670 209.435 ;
        RECT 172.500 208.905 172.670 209.075 ;
        RECT 172.500 208.545 172.670 208.715 ;
        RECT 183.080 209.625 183.250 209.795 ;
        RECT 183.080 209.265 183.250 209.435 ;
        RECT 183.080 208.905 183.250 209.075 ;
        RECT 183.080 208.545 183.250 208.715 ;
        RECT 172.500 204.155 172.670 204.325 ;
        RECT 172.500 203.795 172.670 203.965 ;
        RECT 172.500 203.435 172.670 203.605 ;
        RECT 172.500 203.075 172.670 203.245 ;
        RECT 183.080 204.155 183.250 204.325 ;
        RECT 183.080 203.795 183.250 203.965 ;
        RECT 183.080 203.435 183.250 203.605 ;
        RECT 183.080 203.075 183.250 203.245 ;
        RECT 172.500 198.685 172.670 198.855 ;
        RECT 172.500 198.325 172.670 198.495 ;
        RECT 172.500 197.965 172.670 198.135 ;
        RECT 172.500 197.605 172.670 197.775 ;
        RECT 183.080 198.685 183.250 198.855 ;
        RECT 183.080 198.325 183.250 198.495 ;
        RECT 183.080 197.965 183.250 198.135 ;
        RECT 183.080 197.605 183.250 197.775 ;
        RECT 161.110 193.185 161.280 193.355 ;
        RECT 139.950 192.825 140.120 192.995 ;
        RECT 139.950 192.465 140.120 192.635 ;
        RECT 139.950 192.105 140.120 192.275 ;
        RECT 150.530 192.825 150.700 192.995 ;
        RECT 150.530 192.465 150.700 192.635 ;
        RECT 150.530 192.105 150.700 192.275 ;
        RECT 161.110 192.825 161.280 192.995 ;
        RECT 161.110 192.465 161.280 192.635 ;
        RECT 172.500 193.215 172.670 193.385 ;
        RECT 183.080 193.215 183.250 193.385 ;
        RECT 193.660 214.735 193.830 214.905 ;
        RECT 193.660 214.375 193.830 214.545 ;
        RECT 193.660 214.015 193.830 214.185 ;
        RECT 193.660 209.625 193.830 209.795 ;
        RECT 193.660 209.265 193.830 209.435 ;
        RECT 193.660 208.905 193.830 209.075 ;
        RECT 193.660 208.545 193.830 208.715 ;
        RECT 193.660 204.155 193.830 204.325 ;
        RECT 193.660 203.795 193.830 203.965 ;
        RECT 193.660 203.435 193.830 203.605 ;
        RECT 193.660 203.075 193.830 203.245 ;
        RECT 193.660 198.685 193.830 198.855 ;
        RECT 193.660 198.325 193.830 198.495 ;
        RECT 193.660 197.965 193.830 198.135 ;
        RECT 193.660 197.605 193.830 197.775 ;
        RECT 193.660 193.215 193.830 193.385 ;
        RECT 172.500 192.855 172.670 193.025 ;
        RECT 172.500 192.495 172.670 192.665 ;
        RECT 183.080 192.855 183.250 193.025 ;
        RECT 161.110 192.105 161.280 192.275 ;
        RECT 172.500 192.135 172.670 192.305 ;
        RECT 183.080 192.495 183.250 192.665 ;
        RECT 183.080 192.135 183.250 192.305 ;
        RECT 193.660 192.855 193.830 193.025 ;
        RECT 193.660 192.495 193.830 192.665 ;
        RECT 193.660 192.135 193.830 192.305 ;
        RECT 107.340 185.905 107.510 186.075 ;
        RECT 117.920 185.905 118.090 186.075 ;
        RECT 128.500 185.905 128.670 186.075 ;
        RECT 107.340 185.545 107.510 185.715 ;
        RECT 139.950 185.985 140.120 186.155 ;
        RECT 150.530 185.985 150.700 186.155 ;
        RECT 161.110 185.985 161.280 186.155 ;
        RECT 107.340 185.185 107.510 185.355 ;
        RECT 107.340 184.825 107.510 184.995 ;
        RECT 117.920 185.545 118.090 185.715 ;
        RECT 117.920 185.185 118.090 185.355 ;
        RECT 117.920 184.825 118.090 184.995 ;
        RECT 107.340 180.435 107.510 180.605 ;
        RECT 107.340 180.075 107.510 180.245 ;
        RECT 107.340 179.715 107.510 179.885 ;
        RECT 107.340 179.355 107.510 179.525 ;
        RECT 117.920 180.435 118.090 180.605 ;
        RECT 117.920 180.075 118.090 180.245 ;
        RECT 117.920 179.715 118.090 179.885 ;
        RECT 117.920 179.355 118.090 179.525 ;
        RECT 107.340 174.965 107.510 175.135 ;
        RECT 107.340 174.605 107.510 174.775 ;
        RECT 107.340 174.245 107.510 174.415 ;
        RECT 107.340 173.885 107.510 174.055 ;
        RECT 117.920 174.965 118.090 175.135 ;
        RECT 117.920 174.605 118.090 174.775 ;
        RECT 117.920 174.245 118.090 174.415 ;
        RECT 117.920 173.885 118.090 174.055 ;
        RECT 107.340 169.495 107.510 169.665 ;
        RECT 107.340 169.135 107.510 169.305 ;
        RECT 107.340 168.775 107.510 168.945 ;
        RECT 107.340 168.415 107.510 168.585 ;
        RECT 117.920 169.495 118.090 169.665 ;
        RECT 117.920 169.135 118.090 169.305 ;
        RECT 117.920 168.775 118.090 168.945 ;
        RECT 117.920 168.415 118.090 168.585 ;
        RECT 107.340 164.025 107.510 164.195 ;
        RECT 117.920 164.025 118.090 164.195 ;
        RECT 128.500 185.545 128.670 185.715 ;
        RECT 128.500 185.185 128.670 185.355 ;
        RECT 128.500 184.825 128.670 184.995 ;
        RECT 128.500 180.435 128.670 180.605 ;
        RECT 128.500 180.075 128.670 180.245 ;
        RECT 128.500 179.715 128.670 179.885 ;
        RECT 128.500 179.355 128.670 179.525 ;
        RECT 128.500 174.965 128.670 175.135 ;
        RECT 128.500 174.605 128.670 174.775 ;
        RECT 128.500 174.245 128.670 174.415 ;
        RECT 128.500 173.885 128.670 174.055 ;
        RECT 128.500 169.495 128.670 169.665 ;
        RECT 128.500 169.135 128.670 169.305 ;
        RECT 128.500 168.775 128.670 168.945 ;
        RECT 128.500 168.415 128.670 168.585 ;
        RECT 139.950 185.625 140.120 185.795 ;
        RECT 172.500 186.015 172.670 186.185 ;
        RECT 183.080 186.015 183.250 186.185 ;
        RECT 193.660 186.015 193.830 186.185 ;
        RECT 139.950 185.265 140.120 185.435 ;
        RECT 139.950 184.905 140.120 185.075 ;
        RECT 150.530 185.625 150.700 185.795 ;
        RECT 150.530 185.265 150.700 185.435 ;
        RECT 150.530 184.905 150.700 185.075 ;
        RECT 139.950 180.515 140.120 180.685 ;
        RECT 139.950 180.155 140.120 180.325 ;
        RECT 139.950 179.795 140.120 179.965 ;
        RECT 139.950 179.435 140.120 179.605 ;
        RECT 150.530 180.515 150.700 180.685 ;
        RECT 150.530 180.155 150.700 180.325 ;
        RECT 150.530 179.795 150.700 179.965 ;
        RECT 150.530 179.435 150.700 179.605 ;
        RECT 139.950 175.045 140.120 175.215 ;
        RECT 139.950 174.685 140.120 174.855 ;
        RECT 139.950 174.325 140.120 174.495 ;
        RECT 139.950 173.965 140.120 174.135 ;
        RECT 150.530 175.045 150.700 175.215 ;
        RECT 150.530 174.685 150.700 174.855 ;
        RECT 150.530 174.325 150.700 174.495 ;
        RECT 150.530 173.965 150.700 174.135 ;
        RECT 139.950 169.575 140.120 169.745 ;
        RECT 139.950 169.215 140.120 169.385 ;
        RECT 139.950 168.855 140.120 169.025 ;
        RECT 139.950 168.495 140.120 168.665 ;
        RECT 150.530 169.575 150.700 169.745 ;
        RECT 150.530 169.215 150.700 169.385 ;
        RECT 150.530 168.855 150.700 169.025 ;
        RECT 150.530 168.495 150.700 168.665 ;
        RECT 128.500 164.025 128.670 164.195 ;
        RECT 107.340 163.665 107.510 163.835 ;
        RECT 107.340 163.305 107.510 163.475 ;
        RECT 107.340 162.945 107.510 163.115 ;
        RECT 117.920 163.665 118.090 163.835 ;
        RECT 117.920 163.305 118.090 163.475 ;
        RECT 117.920 162.945 118.090 163.115 ;
        RECT 128.500 163.665 128.670 163.835 ;
        RECT 128.500 163.305 128.670 163.475 ;
        RECT 128.500 162.945 128.670 163.115 ;
        RECT 139.950 164.105 140.120 164.275 ;
        RECT 150.530 164.105 150.700 164.275 ;
        RECT 161.110 185.625 161.280 185.795 ;
        RECT 172.500 185.655 172.670 185.825 ;
        RECT 183.080 185.655 183.250 185.825 ;
        RECT 161.110 185.265 161.280 185.435 ;
        RECT 161.110 184.905 161.280 185.075 ;
        RECT 161.110 180.515 161.280 180.685 ;
        RECT 161.110 180.155 161.280 180.325 ;
        RECT 161.110 179.795 161.280 179.965 ;
        RECT 161.110 179.435 161.280 179.605 ;
        RECT 161.110 175.045 161.280 175.215 ;
        RECT 161.110 174.685 161.280 174.855 ;
        RECT 161.110 174.325 161.280 174.495 ;
        RECT 161.110 173.965 161.280 174.135 ;
        RECT 161.110 169.575 161.280 169.745 ;
        RECT 161.110 169.215 161.280 169.385 ;
        RECT 161.110 168.855 161.280 169.025 ;
        RECT 161.110 168.495 161.280 168.665 ;
        RECT 161.110 164.105 161.280 164.275 ;
        RECT 172.500 185.295 172.670 185.465 ;
        RECT 172.500 184.935 172.670 185.105 ;
        RECT 183.080 185.295 183.250 185.465 ;
        RECT 183.080 184.935 183.250 185.105 ;
        RECT 172.500 180.545 172.670 180.715 ;
        RECT 172.500 180.185 172.670 180.355 ;
        RECT 172.500 179.825 172.670 179.995 ;
        RECT 172.500 179.465 172.670 179.635 ;
        RECT 183.080 180.545 183.250 180.715 ;
        RECT 183.080 180.185 183.250 180.355 ;
        RECT 183.080 179.825 183.250 179.995 ;
        RECT 183.080 179.465 183.250 179.635 ;
        RECT 172.500 175.075 172.670 175.245 ;
        RECT 172.500 174.715 172.670 174.885 ;
        RECT 172.500 174.355 172.670 174.525 ;
        RECT 172.500 173.995 172.670 174.165 ;
        RECT 183.080 175.075 183.250 175.245 ;
        RECT 183.080 174.715 183.250 174.885 ;
        RECT 183.080 174.355 183.250 174.525 ;
        RECT 183.080 173.995 183.250 174.165 ;
        RECT 172.500 169.605 172.670 169.775 ;
        RECT 172.500 169.245 172.670 169.415 ;
        RECT 172.500 168.885 172.670 169.055 ;
        RECT 172.500 168.525 172.670 168.695 ;
        RECT 183.080 169.605 183.250 169.775 ;
        RECT 183.080 169.245 183.250 169.415 ;
        RECT 183.080 168.885 183.250 169.055 ;
        RECT 183.080 168.525 183.250 168.695 ;
        RECT 172.500 164.135 172.670 164.305 ;
        RECT 183.080 164.135 183.250 164.305 ;
        RECT 193.660 185.655 193.830 185.825 ;
        RECT 193.660 185.295 193.830 185.465 ;
        RECT 193.660 184.935 193.830 185.105 ;
        RECT 193.660 180.545 193.830 180.715 ;
        RECT 193.660 180.185 193.830 180.355 ;
        RECT 193.660 179.825 193.830 179.995 ;
        RECT 193.660 179.465 193.830 179.635 ;
        RECT 193.660 175.075 193.830 175.245 ;
        RECT 193.660 174.715 193.830 174.885 ;
        RECT 193.660 174.355 193.830 174.525 ;
        RECT 193.660 173.995 193.830 174.165 ;
        RECT 193.660 169.605 193.830 169.775 ;
        RECT 193.660 169.245 193.830 169.415 ;
        RECT 193.660 168.885 193.830 169.055 ;
        RECT 193.660 168.525 193.830 168.695 ;
        RECT 193.660 164.135 193.830 164.305 ;
        RECT 139.950 163.745 140.120 163.915 ;
        RECT 139.950 163.385 140.120 163.555 ;
        RECT 139.950 163.025 140.120 163.195 ;
        RECT 150.530 163.745 150.700 163.915 ;
        RECT 150.530 163.385 150.700 163.555 ;
        RECT 150.530 163.025 150.700 163.195 ;
        RECT 161.110 163.745 161.280 163.915 ;
        RECT 161.110 163.385 161.280 163.555 ;
        RECT 161.110 163.025 161.280 163.195 ;
        RECT 172.500 163.775 172.670 163.945 ;
        RECT 172.500 163.415 172.670 163.585 ;
        RECT 172.500 163.055 172.670 163.225 ;
        RECT 183.080 163.775 183.250 163.945 ;
        RECT 183.080 163.415 183.250 163.585 ;
        RECT 183.080 163.055 183.250 163.225 ;
        RECT 193.660 163.775 193.830 163.945 ;
        RECT 193.660 163.415 193.830 163.585 ;
        RECT 193.660 163.055 193.830 163.225 ;
        RECT 107.340 156.735 107.510 156.905 ;
        RECT 117.920 156.735 118.090 156.905 ;
        RECT 128.500 156.735 128.670 156.905 ;
        RECT 107.340 156.375 107.510 156.545 ;
        RECT 139.950 156.815 140.120 156.985 ;
        RECT 150.530 156.815 150.700 156.985 ;
        RECT 161.110 156.815 161.280 156.985 ;
        RECT 107.340 156.015 107.510 156.185 ;
        RECT 107.340 155.655 107.510 155.825 ;
        RECT 117.920 156.375 118.090 156.545 ;
        RECT 117.920 156.015 118.090 156.185 ;
        RECT 117.920 155.655 118.090 155.825 ;
        RECT 107.340 151.265 107.510 151.435 ;
        RECT 107.340 150.905 107.510 151.075 ;
        RECT 107.340 150.545 107.510 150.715 ;
        RECT 107.340 150.185 107.510 150.355 ;
        RECT 117.920 151.265 118.090 151.435 ;
        RECT 117.920 150.905 118.090 151.075 ;
        RECT 117.920 150.545 118.090 150.715 ;
        RECT 117.920 150.185 118.090 150.355 ;
        RECT 107.340 145.795 107.510 145.965 ;
        RECT 107.340 145.435 107.510 145.605 ;
        RECT 107.340 145.075 107.510 145.245 ;
        RECT 107.340 144.715 107.510 144.885 ;
        RECT 117.920 145.795 118.090 145.965 ;
        RECT 117.920 145.435 118.090 145.605 ;
        RECT 117.920 145.075 118.090 145.245 ;
        RECT 117.920 144.715 118.090 144.885 ;
        RECT 107.340 140.325 107.510 140.495 ;
        RECT 107.340 139.965 107.510 140.135 ;
        RECT 107.340 139.605 107.510 139.775 ;
        RECT 107.340 139.245 107.510 139.415 ;
        RECT 117.920 140.325 118.090 140.495 ;
        RECT 117.920 139.965 118.090 140.135 ;
        RECT 117.920 139.605 118.090 139.775 ;
        RECT 117.920 139.245 118.090 139.415 ;
        RECT 107.340 134.855 107.510 135.025 ;
        RECT 117.920 134.855 118.090 135.025 ;
        RECT 128.500 156.375 128.670 156.545 ;
        RECT 128.500 156.015 128.670 156.185 ;
        RECT 128.500 155.655 128.670 155.825 ;
        RECT 128.500 151.265 128.670 151.435 ;
        RECT 128.500 150.905 128.670 151.075 ;
        RECT 128.500 150.545 128.670 150.715 ;
        RECT 128.500 150.185 128.670 150.355 ;
        RECT 128.500 145.795 128.670 145.965 ;
        RECT 128.500 145.435 128.670 145.605 ;
        RECT 128.500 145.075 128.670 145.245 ;
        RECT 128.500 144.715 128.670 144.885 ;
        RECT 128.500 140.325 128.670 140.495 ;
        RECT 128.500 139.965 128.670 140.135 ;
        RECT 128.500 139.605 128.670 139.775 ;
        RECT 128.500 139.245 128.670 139.415 ;
        RECT 139.950 156.455 140.120 156.625 ;
        RECT 172.500 156.845 172.670 157.015 ;
        RECT 183.080 156.845 183.250 157.015 ;
        RECT 193.660 156.845 193.830 157.015 ;
        RECT 139.950 156.095 140.120 156.265 ;
        RECT 139.950 155.735 140.120 155.905 ;
        RECT 150.530 156.455 150.700 156.625 ;
        RECT 150.530 156.095 150.700 156.265 ;
        RECT 150.530 155.735 150.700 155.905 ;
        RECT 139.950 151.345 140.120 151.515 ;
        RECT 139.950 150.985 140.120 151.155 ;
        RECT 139.950 150.625 140.120 150.795 ;
        RECT 139.950 150.265 140.120 150.435 ;
        RECT 150.530 151.345 150.700 151.515 ;
        RECT 150.530 150.985 150.700 151.155 ;
        RECT 150.530 150.625 150.700 150.795 ;
        RECT 150.530 150.265 150.700 150.435 ;
        RECT 139.950 145.875 140.120 146.045 ;
        RECT 139.950 145.515 140.120 145.685 ;
        RECT 139.950 145.155 140.120 145.325 ;
        RECT 139.950 144.795 140.120 144.965 ;
        RECT 150.530 145.875 150.700 146.045 ;
        RECT 150.530 145.515 150.700 145.685 ;
        RECT 150.530 145.155 150.700 145.325 ;
        RECT 150.530 144.795 150.700 144.965 ;
        RECT 139.950 140.405 140.120 140.575 ;
        RECT 139.950 140.045 140.120 140.215 ;
        RECT 139.950 139.685 140.120 139.855 ;
        RECT 139.950 139.325 140.120 139.495 ;
        RECT 150.530 140.405 150.700 140.575 ;
        RECT 150.530 140.045 150.700 140.215 ;
        RECT 150.530 139.685 150.700 139.855 ;
        RECT 150.530 139.325 150.700 139.495 ;
        RECT 128.500 134.855 128.670 135.025 ;
        RECT 107.340 134.495 107.510 134.665 ;
        RECT 107.340 134.135 107.510 134.305 ;
        RECT 107.340 133.775 107.510 133.945 ;
        RECT 117.920 134.495 118.090 134.665 ;
        RECT 117.920 134.135 118.090 134.305 ;
        RECT 117.920 133.775 118.090 133.945 ;
        RECT 128.500 134.495 128.670 134.665 ;
        RECT 128.500 134.135 128.670 134.305 ;
        RECT 128.500 133.775 128.670 133.945 ;
        RECT 139.950 134.935 140.120 135.105 ;
        RECT 150.530 134.935 150.700 135.105 ;
        RECT 161.110 156.455 161.280 156.625 ;
        RECT 161.110 156.095 161.280 156.265 ;
        RECT 161.110 155.735 161.280 155.905 ;
        RECT 161.110 151.345 161.280 151.515 ;
        RECT 161.110 150.985 161.280 151.155 ;
        RECT 161.110 150.625 161.280 150.795 ;
        RECT 161.110 150.265 161.280 150.435 ;
        RECT 161.110 145.875 161.280 146.045 ;
        RECT 161.110 145.515 161.280 145.685 ;
        RECT 161.110 145.155 161.280 145.325 ;
        RECT 161.110 144.795 161.280 144.965 ;
        RECT 161.110 140.405 161.280 140.575 ;
        RECT 161.110 140.045 161.280 140.215 ;
        RECT 161.110 139.685 161.280 139.855 ;
        RECT 161.110 139.325 161.280 139.495 ;
        RECT 161.110 134.935 161.280 135.105 ;
        RECT 172.500 156.485 172.670 156.655 ;
        RECT 172.500 156.125 172.670 156.295 ;
        RECT 172.500 155.765 172.670 155.935 ;
        RECT 183.080 156.485 183.250 156.655 ;
        RECT 183.080 156.125 183.250 156.295 ;
        RECT 183.080 155.765 183.250 155.935 ;
        RECT 172.500 151.375 172.670 151.545 ;
        RECT 172.500 151.015 172.670 151.185 ;
        RECT 172.500 150.655 172.670 150.825 ;
        RECT 172.500 150.295 172.670 150.465 ;
        RECT 183.080 151.375 183.250 151.545 ;
        RECT 183.080 151.015 183.250 151.185 ;
        RECT 183.080 150.655 183.250 150.825 ;
        RECT 183.080 150.295 183.250 150.465 ;
        RECT 172.500 145.905 172.670 146.075 ;
        RECT 172.500 145.545 172.670 145.715 ;
        RECT 172.500 145.185 172.670 145.355 ;
        RECT 172.500 144.825 172.670 144.995 ;
        RECT 183.080 145.905 183.250 146.075 ;
        RECT 183.080 145.545 183.250 145.715 ;
        RECT 183.080 145.185 183.250 145.355 ;
        RECT 183.080 144.825 183.250 144.995 ;
        RECT 172.500 140.435 172.670 140.605 ;
        RECT 172.500 140.075 172.670 140.245 ;
        RECT 172.500 139.715 172.670 139.885 ;
        RECT 172.500 139.355 172.670 139.525 ;
        RECT 183.080 140.435 183.250 140.605 ;
        RECT 183.080 140.075 183.250 140.245 ;
        RECT 183.080 139.715 183.250 139.885 ;
        RECT 183.080 139.355 183.250 139.525 ;
        RECT 172.500 134.965 172.670 135.135 ;
        RECT 183.080 134.965 183.250 135.135 ;
        RECT 193.660 156.485 193.830 156.655 ;
        RECT 193.660 156.125 193.830 156.295 ;
        RECT 193.660 155.765 193.830 155.935 ;
        RECT 193.660 151.375 193.830 151.545 ;
        RECT 193.660 151.015 193.830 151.185 ;
        RECT 193.660 150.655 193.830 150.825 ;
        RECT 193.660 150.295 193.830 150.465 ;
        RECT 193.660 145.905 193.830 146.075 ;
        RECT 193.660 145.545 193.830 145.715 ;
        RECT 193.660 145.185 193.830 145.355 ;
        RECT 193.660 144.825 193.830 144.995 ;
        RECT 193.660 140.435 193.830 140.605 ;
        RECT 193.660 140.075 193.830 140.245 ;
        RECT 193.660 139.715 193.830 139.885 ;
        RECT 193.660 139.355 193.830 139.525 ;
        RECT 193.660 134.965 193.830 135.135 ;
        RECT 139.950 134.575 140.120 134.745 ;
        RECT 139.950 134.215 140.120 134.385 ;
        RECT 139.950 133.855 140.120 134.025 ;
        RECT 150.530 134.575 150.700 134.745 ;
        RECT 150.530 134.215 150.700 134.385 ;
        RECT 150.530 133.855 150.700 134.025 ;
        RECT 161.110 134.575 161.280 134.745 ;
        RECT 161.110 134.215 161.280 134.385 ;
        RECT 161.110 133.855 161.280 134.025 ;
        RECT 172.500 134.605 172.670 134.775 ;
        RECT 172.500 134.245 172.670 134.415 ;
        RECT 172.500 133.885 172.670 134.055 ;
        RECT 183.080 134.605 183.250 134.775 ;
        RECT 183.080 134.245 183.250 134.415 ;
        RECT 183.080 133.885 183.250 134.055 ;
        RECT 193.660 134.605 193.830 134.775 ;
        RECT 193.660 134.245 193.830 134.415 ;
        RECT 193.660 133.885 193.830 134.055 ;
        RECT 107.340 127.555 107.510 127.725 ;
        RECT 117.920 127.555 118.090 127.725 ;
        RECT 128.500 127.555 128.670 127.725 ;
        RECT 107.340 127.195 107.510 127.365 ;
        RECT 139.950 127.635 140.120 127.805 ;
        RECT 150.530 127.635 150.700 127.805 ;
        RECT 161.110 127.635 161.280 127.805 ;
        RECT 107.340 126.835 107.510 127.005 ;
        RECT 107.340 126.475 107.510 126.645 ;
        RECT 117.920 127.195 118.090 127.365 ;
        RECT 117.920 126.835 118.090 127.005 ;
        RECT 117.920 126.475 118.090 126.645 ;
        RECT 107.340 122.085 107.510 122.255 ;
        RECT 107.340 121.725 107.510 121.895 ;
        RECT 107.340 121.365 107.510 121.535 ;
        RECT 107.340 121.005 107.510 121.175 ;
        RECT 117.920 122.085 118.090 122.255 ;
        RECT 117.920 121.725 118.090 121.895 ;
        RECT 117.920 121.365 118.090 121.535 ;
        RECT 117.920 121.005 118.090 121.175 ;
        RECT 107.340 116.615 107.510 116.785 ;
        RECT 107.340 116.255 107.510 116.425 ;
        RECT 107.340 115.895 107.510 116.065 ;
        RECT 107.340 115.535 107.510 115.705 ;
        RECT 117.920 116.615 118.090 116.785 ;
        RECT 117.920 116.255 118.090 116.425 ;
        RECT 117.920 115.895 118.090 116.065 ;
        RECT 117.920 115.535 118.090 115.705 ;
        RECT 107.340 111.145 107.510 111.315 ;
        RECT 107.340 110.785 107.510 110.955 ;
        RECT 107.340 110.425 107.510 110.595 ;
        RECT 107.340 110.065 107.510 110.235 ;
        RECT 117.920 111.145 118.090 111.315 ;
        RECT 117.920 110.785 118.090 110.955 ;
        RECT 117.920 110.425 118.090 110.595 ;
        RECT 117.920 110.065 118.090 110.235 ;
        RECT 107.340 105.675 107.510 105.845 ;
        RECT 117.920 105.675 118.090 105.845 ;
        RECT 128.500 127.195 128.670 127.365 ;
        RECT 128.500 126.835 128.670 127.005 ;
        RECT 128.500 126.475 128.670 126.645 ;
        RECT 128.500 122.085 128.670 122.255 ;
        RECT 128.500 121.725 128.670 121.895 ;
        RECT 128.500 121.365 128.670 121.535 ;
        RECT 128.500 121.005 128.670 121.175 ;
        RECT 128.500 116.615 128.670 116.785 ;
        RECT 128.500 116.255 128.670 116.425 ;
        RECT 128.500 115.895 128.670 116.065 ;
        RECT 128.500 115.535 128.670 115.705 ;
        RECT 128.500 111.145 128.670 111.315 ;
        RECT 128.500 110.785 128.670 110.955 ;
        RECT 128.500 110.425 128.670 110.595 ;
        RECT 128.500 110.065 128.670 110.235 ;
        RECT 139.950 127.275 140.120 127.445 ;
        RECT 172.500 127.665 172.670 127.835 ;
        RECT 183.080 127.665 183.250 127.835 ;
        RECT 193.660 127.665 193.830 127.835 ;
        RECT 139.950 126.915 140.120 127.085 ;
        RECT 139.950 126.555 140.120 126.725 ;
        RECT 150.530 127.275 150.700 127.445 ;
        RECT 150.530 126.915 150.700 127.085 ;
        RECT 150.530 126.555 150.700 126.725 ;
        RECT 139.950 122.165 140.120 122.335 ;
        RECT 139.950 121.805 140.120 121.975 ;
        RECT 139.950 121.445 140.120 121.615 ;
        RECT 139.950 121.085 140.120 121.255 ;
        RECT 150.530 122.165 150.700 122.335 ;
        RECT 150.530 121.805 150.700 121.975 ;
        RECT 150.530 121.445 150.700 121.615 ;
        RECT 150.530 121.085 150.700 121.255 ;
        RECT 139.950 116.695 140.120 116.865 ;
        RECT 139.950 116.335 140.120 116.505 ;
        RECT 139.950 115.975 140.120 116.145 ;
        RECT 139.950 115.615 140.120 115.785 ;
        RECT 150.530 116.695 150.700 116.865 ;
        RECT 150.530 116.335 150.700 116.505 ;
        RECT 150.530 115.975 150.700 116.145 ;
        RECT 150.530 115.615 150.700 115.785 ;
        RECT 139.950 111.225 140.120 111.395 ;
        RECT 139.950 110.865 140.120 111.035 ;
        RECT 139.950 110.505 140.120 110.675 ;
        RECT 139.950 110.145 140.120 110.315 ;
        RECT 150.530 111.225 150.700 111.395 ;
        RECT 150.530 110.865 150.700 111.035 ;
        RECT 150.530 110.505 150.700 110.675 ;
        RECT 150.530 110.145 150.700 110.315 ;
        RECT 128.500 105.675 128.670 105.845 ;
        RECT 107.340 105.315 107.510 105.485 ;
        RECT 107.340 104.955 107.510 105.125 ;
        RECT 107.340 104.595 107.510 104.765 ;
        RECT 117.920 105.315 118.090 105.485 ;
        RECT 117.920 104.955 118.090 105.125 ;
        RECT 117.920 104.595 118.090 104.765 ;
        RECT 128.500 105.315 128.670 105.485 ;
        RECT 128.500 104.955 128.670 105.125 ;
        RECT 128.500 104.595 128.670 104.765 ;
        RECT 139.950 105.755 140.120 105.925 ;
        RECT 150.530 105.755 150.700 105.925 ;
        RECT 161.110 127.275 161.280 127.445 ;
        RECT 161.110 126.915 161.280 127.085 ;
        RECT 161.110 126.555 161.280 126.725 ;
        RECT 161.110 122.165 161.280 122.335 ;
        RECT 161.110 121.805 161.280 121.975 ;
        RECT 161.110 121.445 161.280 121.615 ;
        RECT 161.110 121.085 161.280 121.255 ;
        RECT 161.110 116.695 161.280 116.865 ;
        RECT 161.110 116.335 161.280 116.505 ;
        RECT 161.110 115.975 161.280 116.145 ;
        RECT 161.110 115.615 161.280 115.785 ;
        RECT 161.110 111.225 161.280 111.395 ;
        RECT 161.110 110.865 161.280 111.035 ;
        RECT 161.110 110.505 161.280 110.675 ;
        RECT 161.110 110.145 161.280 110.315 ;
        RECT 161.110 105.755 161.280 105.925 ;
        RECT 172.500 127.305 172.670 127.475 ;
        RECT 172.500 126.945 172.670 127.115 ;
        RECT 172.500 126.585 172.670 126.755 ;
        RECT 183.080 127.305 183.250 127.475 ;
        RECT 183.080 126.945 183.250 127.115 ;
        RECT 183.080 126.585 183.250 126.755 ;
        RECT 172.500 122.195 172.670 122.365 ;
        RECT 172.500 121.835 172.670 122.005 ;
        RECT 172.500 121.475 172.670 121.645 ;
        RECT 172.500 121.115 172.670 121.285 ;
        RECT 183.080 122.195 183.250 122.365 ;
        RECT 183.080 121.835 183.250 122.005 ;
        RECT 183.080 121.475 183.250 121.645 ;
        RECT 183.080 121.115 183.250 121.285 ;
        RECT 172.500 116.725 172.670 116.895 ;
        RECT 172.500 116.365 172.670 116.535 ;
        RECT 172.500 116.005 172.670 116.175 ;
        RECT 172.500 115.645 172.670 115.815 ;
        RECT 183.080 116.725 183.250 116.895 ;
        RECT 183.080 116.365 183.250 116.535 ;
        RECT 183.080 116.005 183.250 116.175 ;
        RECT 183.080 115.645 183.250 115.815 ;
        RECT 172.500 111.255 172.670 111.425 ;
        RECT 172.500 110.895 172.670 111.065 ;
        RECT 172.500 110.535 172.670 110.705 ;
        RECT 172.500 110.175 172.670 110.345 ;
        RECT 183.080 111.255 183.250 111.425 ;
        RECT 183.080 110.895 183.250 111.065 ;
        RECT 183.080 110.535 183.250 110.705 ;
        RECT 183.080 110.175 183.250 110.345 ;
        RECT 139.950 105.395 140.120 105.565 ;
        RECT 139.950 105.035 140.120 105.205 ;
        RECT 139.950 104.675 140.120 104.845 ;
        RECT 150.530 105.395 150.700 105.565 ;
        RECT 150.530 105.035 150.700 105.205 ;
        RECT 150.530 104.675 150.700 104.845 ;
        RECT 161.110 105.395 161.280 105.565 ;
        RECT 161.110 105.035 161.280 105.205 ;
        RECT 161.110 104.675 161.280 104.845 ;
        RECT 172.500 105.785 172.670 105.955 ;
        RECT 183.080 105.785 183.250 105.955 ;
        RECT 193.660 127.305 193.830 127.475 ;
        RECT 193.660 126.945 193.830 127.115 ;
        RECT 193.660 126.585 193.830 126.755 ;
        RECT 193.660 122.195 193.830 122.365 ;
        RECT 193.660 121.835 193.830 122.005 ;
        RECT 193.660 121.475 193.830 121.645 ;
        RECT 193.660 121.115 193.830 121.285 ;
        RECT 193.660 116.725 193.830 116.895 ;
        RECT 193.660 116.365 193.830 116.535 ;
        RECT 193.660 116.005 193.830 116.175 ;
        RECT 193.660 115.645 193.830 115.815 ;
        RECT 193.660 111.255 193.830 111.425 ;
        RECT 193.660 110.895 193.830 111.065 ;
        RECT 193.660 110.535 193.830 110.705 ;
        RECT 193.660 110.175 193.830 110.345 ;
        RECT 193.660 105.785 193.830 105.955 ;
        RECT 172.500 105.425 172.670 105.595 ;
        RECT 172.500 105.065 172.670 105.235 ;
        RECT 172.500 104.705 172.670 104.875 ;
        RECT 183.080 105.425 183.250 105.595 ;
        RECT 183.080 105.065 183.250 105.235 ;
        RECT 183.080 104.705 183.250 104.875 ;
        RECT 193.660 105.425 193.830 105.595 ;
        RECT 193.660 105.065 193.830 105.235 ;
        RECT 193.660 104.705 193.830 104.875 ;
        RECT 107.340 98.235 107.510 98.405 ;
        RECT 117.920 98.235 118.090 98.405 ;
        RECT 128.500 98.235 128.670 98.405 ;
        RECT 107.340 97.875 107.510 98.045 ;
        RECT 139.950 98.315 140.120 98.485 ;
        RECT 150.530 98.315 150.700 98.485 ;
        RECT 161.110 98.315 161.280 98.485 ;
        RECT 107.340 97.515 107.510 97.685 ;
        RECT 107.340 97.155 107.510 97.325 ;
        RECT 117.920 97.875 118.090 98.045 ;
        RECT 117.920 97.515 118.090 97.685 ;
        RECT 117.920 97.155 118.090 97.325 ;
        RECT 107.340 92.765 107.510 92.935 ;
        RECT 107.340 92.405 107.510 92.575 ;
        RECT 107.340 92.045 107.510 92.215 ;
        RECT 107.340 91.685 107.510 91.855 ;
        RECT 117.920 92.765 118.090 92.935 ;
        RECT 117.920 92.405 118.090 92.575 ;
        RECT 117.920 92.045 118.090 92.215 ;
        RECT 117.920 91.685 118.090 91.855 ;
        RECT 107.340 87.295 107.510 87.465 ;
        RECT 107.340 86.935 107.510 87.105 ;
        RECT 107.340 86.575 107.510 86.745 ;
        RECT 107.340 86.215 107.510 86.385 ;
        RECT 117.920 87.295 118.090 87.465 ;
        RECT 117.920 86.935 118.090 87.105 ;
        RECT 117.920 86.575 118.090 86.745 ;
        RECT 117.920 86.215 118.090 86.385 ;
        RECT 107.340 81.825 107.510 81.995 ;
        RECT 107.340 81.465 107.510 81.635 ;
        RECT 107.340 81.105 107.510 81.275 ;
        RECT 107.340 80.745 107.510 80.915 ;
        RECT 117.920 81.825 118.090 81.995 ;
        RECT 117.920 81.465 118.090 81.635 ;
        RECT 117.920 81.105 118.090 81.275 ;
        RECT 117.920 80.745 118.090 80.915 ;
        RECT 107.340 76.355 107.510 76.525 ;
        RECT 117.920 76.355 118.090 76.525 ;
        RECT 128.500 97.875 128.670 98.045 ;
        RECT 128.500 97.515 128.670 97.685 ;
        RECT 128.500 97.155 128.670 97.325 ;
        RECT 128.500 92.765 128.670 92.935 ;
        RECT 128.500 92.405 128.670 92.575 ;
        RECT 128.500 92.045 128.670 92.215 ;
        RECT 128.500 91.685 128.670 91.855 ;
        RECT 128.500 87.295 128.670 87.465 ;
        RECT 128.500 86.935 128.670 87.105 ;
        RECT 128.500 86.575 128.670 86.745 ;
        RECT 128.500 86.215 128.670 86.385 ;
        RECT 128.500 81.825 128.670 81.995 ;
        RECT 128.500 81.465 128.670 81.635 ;
        RECT 128.500 81.105 128.670 81.275 ;
        RECT 128.500 80.745 128.670 80.915 ;
        RECT 139.950 97.955 140.120 98.125 ;
        RECT 172.500 98.345 172.670 98.515 ;
        RECT 183.080 98.345 183.250 98.515 ;
        RECT 193.660 98.345 193.830 98.515 ;
        RECT 139.950 97.595 140.120 97.765 ;
        RECT 139.950 97.235 140.120 97.405 ;
        RECT 150.530 97.955 150.700 98.125 ;
        RECT 150.530 97.595 150.700 97.765 ;
        RECT 150.530 97.235 150.700 97.405 ;
        RECT 139.950 92.845 140.120 93.015 ;
        RECT 139.950 92.485 140.120 92.655 ;
        RECT 139.950 92.125 140.120 92.295 ;
        RECT 139.950 91.765 140.120 91.935 ;
        RECT 150.530 92.845 150.700 93.015 ;
        RECT 150.530 92.485 150.700 92.655 ;
        RECT 150.530 92.125 150.700 92.295 ;
        RECT 150.530 91.765 150.700 91.935 ;
        RECT 139.950 87.375 140.120 87.545 ;
        RECT 139.950 87.015 140.120 87.185 ;
        RECT 139.950 86.655 140.120 86.825 ;
        RECT 139.950 86.295 140.120 86.465 ;
        RECT 150.530 87.375 150.700 87.545 ;
        RECT 150.530 87.015 150.700 87.185 ;
        RECT 150.530 86.655 150.700 86.825 ;
        RECT 150.530 86.295 150.700 86.465 ;
        RECT 139.950 81.905 140.120 82.075 ;
        RECT 139.950 81.545 140.120 81.715 ;
        RECT 139.950 81.185 140.120 81.355 ;
        RECT 139.950 80.825 140.120 80.995 ;
        RECT 150.530 81.905 150.700 82.075 ;
        RECT 150.530 81.545 150.700 81.715 ;
        RECT 150.530 81.185 150.700 81.355 ;
        RECT 150.530 80.825 150.700 80.995 ;
        RECT 128.500 76.355 128.670 76.525 ;
        RECT 107.340 75.995 107.510 76.165 ;
        RECT 107.340 75.635 107.510 75.805 ;
        RECT 107.340 75.275 107.510 75.445 ;
        RECT 117.920 75.995 118.090 76.165 ;
        RECT 117.920 75.635 118.090 75.805 ;
        RECT 117.920 75.275 118.090 75.445 ;
        RECT 128.500 75.995 128.670 76.165 ;
        RECT 128.500 75.635 128.670 75.805 ;
        RECT 128.500 75.275 128.670 75.445 ;
        RECT 139.950 76.435 140.120 76.605 ;
        RECT 150.530 76.435 150.700 76.605 ;
        RECT 161.110 97.955 161.280 98.125 ;
        RECT 161.110 97.595 161.280 97.765 ;
        RECT 161.110 97.235 161.280 97.405 ;
        RECT 161.110 92.845 161.280 93.015 ;
        RECT 161.110 92.485 161.280 92.655 ;
        RECT 161.110 92.125 161.280 92.295 ;
        RECT 161.110 91.765 161.280 91.935 ;
        RECT 161.110 87.375 161.280 87.545 ;
        RECT 161.110 87.015 161.280 87.185 ;
        RECT 161.110 86.655 161.280 86.825 ;
        RECT 161.110 86.295 161.280 86.465 ;
        RECT 161.110 81.905 161.280 82.075 ;
        RECT 161.110 81.545 161.280 81.715 ;
        RECT 161.110 81.185 161.280 81.355 ;
        RECT 161.110 80.825 161.280 80.995 ;
        RECT 161.110 76.435 161.280 76.605 ;
        RECT 172.500 97.985 172.670 98.155 ;
        RECT 172.500 97.625 172.670 97.795 ;
        RECT 172.500 97.265 172.670 97.435 ;
        RECT 183.080 97.985 183.250 98.155 ;
        RECT 183.080 97.625 183.250 97.795 ;
        RECT 183.080 97.265 183.250 97.435 ;
        RECT 172.500 92.875 172.670 93.045 ;
        RECT 172.500 92.515 172.670 92.685 ;
        RECT 172.500 92.155 172.670 92.325 ;
        RECT 172.500 91.795 172.670 91.965 ;
        RECT 183.080 92.875 183.250 93.045 ;
        RECT 183.080 92.515 183.250 92.685 ;
        RECT 183.080 92.155 183.250 92.325 ;
        RECT 183.080 91.795 183.250 91.965 ;
        RECT 172.500 87.405 172.670 87.575 ;
        RECT 172.500 87.045 172.670 87.215 ;
        RECT 172.500 86.685 172.670 86.855 ;
        RECT 172.500 86.325 172.670 86.495 ;
        RECT 183.080 87.405 183.250 87.575 ;
        RECT 183.080 87.045 183.250 87.215 ;
        RECT 183.080 86.685 183.250 86.855 ;
        RECT 183.080 86.325 183.250 86.495 ;
        RECT 172.500 81.935 172.670 82.105 ;
        RECT 172.500 81.575 172.670 81.745 ;
        RECT 172.500 81.215 172.670 81.385 ;
        RECT 172.500 80.855 172.670 81.025 ;
        RECT 183.080 81.935 183.250 82.105 ;
        RECT 183.080 81.575 183.250 81.745 ;
        RECT 183.080 81.215 183.250 81.385 ;
        RECT 183.080 80.855 183.250 81.025 ;
        RECT 172.500 76.465 172.670 76.635 ;
        RECT 183.080 76.465 183.250 76.635 ;
        RECT 193.660 97.985 193.830 98.155 ;
        RECT 193.660 97.625 193.830 97.795 ;
        RECT 193.660 97.265 193.830 97.435 ;
        RECT 193.660 92.875 193.830 93.045 ;
        RECT 193.660 92.515 193.830 92.685 ;
        RECT 193.660 92.155 193.830 92.325 ;
        RECT 193.660 91.795 193.830 91.965 ;
        RECT 193.660 87.405 193.830 87.575 ;
        RECT 193.660 87.045 193.830 87.215 ;
        RECT 193.660 86.685 193.830 86.855 ;
        RECT 193.660 86.325 193.830 86.495 ;
        RECT 193.660 81.935 193.830 82.105 ;
        RECT 193.660 81.575 193.830 81.745 ;
        RECT 193.660 81.215 193.830 81.385 ;
        RECT 193.660 80.855 193.830 81.025 ;
        RECT 193.660 76.465 193.830 76.635 ;
        RECT 139.950 76.075 140.120 76.245 ;
        RECT 139.950 75.715 140.120 75.885 ;
        RECT 139.950 75.355 140.120 75.525 ;
        RECT 150.530 76.075 150.700 76.245 ;
        RECT 150.530 75.715 150.700 75.885 ;
        RECT 150.530 75.355 150.700 75.525 ;
        RECT 161.110 76.075 161.280 76.245 ;
        RECT 161.110 75.715 161.280 75.885 ;
        RECT 161.110 75.355 161.280 75.525 ;
        RECT 172.500 76.105 172.670 76.275 ;
        RECT 172.500 75.745 172.670 75.915 ;
        RECT 172.500 75.385 172.670 75.555 ;
        RECT 183.080 76.105 183.250 76.275 ;
        RECT 183.080 75.745 183.250 75.915 ;
        RECT 183.080 75.385 183.250 75.555 ;
        RECT 193.660 76.105 193.830 76.275 ;
        RECT 193.660 75.745 193.830 75.915 ;
        RECT 193.660 75.385 193.830 75.555 ;
        RECT 107.390 68.955 107.560 69.125 ;
        RECT 117.970 68.955 118.140 69.125 ;
        RECT 128.550 68.955 128.720 69.125 ;
        RECT 107.390 68.595 107.560 68.765 ;
        RECT 140.000 69.035 140.170 69.205 ;
        RECT 150.580 69.035 150.750 69.205 ;
        RECT 161.160 69.035 161.330 69.205 ;
        RECT 107.390 68.235 107.560 68.405 ;
        RECT 107.390 67.875 107.560 68.045 ;
        RECT 117.970 68.595 118.140 68.765 ;
        RECT 117.970 68.235 118.140 68.405 ;
        RECT 117.970 67.875 118.140 68.045 ;
        RECT 107.390 63.485 107.560 63.655 ;
        RECT 107.390 63.125 107.560 63.295 ;
        RECT 107.390 62.765 107.560 62.935 ;
        RECT 107.390 62.405 107.560 62.575 ;
        RECT 117.970 63.485 118.140 63.655 ;
        RECT 117.970 63.125 118.140 63.295 ;
        RECT 117.970 62.765 118.140 62.935 ;
        RECT 117.970 62.405 118.140 62.575 ;
        RECT 107.390 58.015 107.560 58.185 ;
        RECT 107.390 57.655 107.560 57.825 ;
        RECT 107.390 57.295 107.560 57.465 ;
        RECT 107.390 56.935 107.560 57.105 ;
        RECT 117.970 58.015 118.140 58.185 ;
        RECT 117.970 57.655 118.140 57.825 ;
        RECT 117.970 57.295 118.140 57.465 ;
        RECT 117.970 56.935 118.140 57.105 ;
        RECT 107.390 52.545 107.560 52.715 ;
        RECT 107.390 52.185 107.560 52.355 ;
        RECT 107.390 51.825 107.560 51.995 ;
        RECT 107.390 51.465 107.560 51.635 ;
        RECT 117.970 52.545 118.140 52.715 ;
        RECT 117.970 52.185 118.140 52.355 ;
        RECT 117.970 51.825 118.140 51.995 ;
        RECT 117.970 51.465 118.140 51.635 ;
        RECT 107.390 47.075 107.560 47.245 ;
        RECT 117.970 47.075 118.140 47.245 ;
        RECT 128.550 68.595 128.720 68.765 ;
        RECT 128.550 68.235 128.720 68.405 ;
        RECT 128.550 67.875 128.720 68.045 ;
        RECT 128.550 63.485 128.720 63.655 ;
        RECT 128.550 63.125 128.720 63.295 ;
        RECT 128.550 62.765 128.720 62.935 ;
        RECT 128.550 62.405 128.720 62.575 ;
        RECT 128.550 58.015 128.720 58.185 ;
        RECT 128.550 57.655 128.720 57.825 ;
        RECT 128.550 57.295 128.720 57.465 ;
        RECT 128.550 56.935 128.720 57.105 ;
        RECT 128.550 52.545 128.720 52.715 ;
        RECT 128.550 52.185 128.720 52.355 ;
        RECT 128.550 51.825 128.720 51.995 ;
        RECT 128.550 51.465 128.720 51.635 ;
        RECT 140.000 68.675 140.170 68.845 ;
        RECT 172.550 69.065 172.720 69.235 ;
        RECT 183.130 69.065 183.300 69.235 ;
        RECT 193.710 69.065 193.880 69.235 ;
        RECT 140.000 68.315 140.170 68.485 ;
        RECT 140.000 67.955 140.170 68.125 ;
        RECT 150.580 68.675 150.750 68.845 ;
        RECT 150.580 68.315 150.750 68.485 ;
        RECT 150.580 67.955 150.750 68.125 ;
        RECT 140.000 63.565 140.170 63.735 ;
        RECT 140.000 63.205 140.170 63.375 ;
        RECT 140.000 62.845 140.170 63.015 ;
        RECT 140.000 62.485 140.170 62.655 ;
        RECT 150.580 63.565 150.750 63.735 ;
        RECT 150.580 63.205 150.750 63.375 ;
        RECT 150.580 62.845 150.750 63.015 ;
        RECT 150.580 62.485 150.750 62.655 ;
        RECT 140.000 58.095 140.170 58.265 ;
        RECT 140.000 57.735 140.170 57.905 ;
        RECT 140.000 57.375 140.170 57.545 ;
        RECT 140.000 57.015 140.170 57.185 ;
        RECT 150.580 58.095 150.750 58.265 ;
        RECT 150.580 57.735 150.750 57.905 ;
        RECT 150.580 57.375 150.750 57.545 ;
        RECT 150.580 57.015 150.750 57.185 ;
        RECT 140.000 52.625 140.170 52.795 ;
        RECT 140.000 52.265 140.170 52.435 ;
        RECT 140.000 51.905 140.170 52.075 ;
        RECT 140.000 51.545 140.170 51.715 ;
        RECT 150.580 52.625 150.750 52.795 ;
        RECT 150.580 52.265 150.750 52.435 ;
        RECT 150.580 51.905 150.750 52.075 ;
        RECT 150.580 51.545 150.750 51.715 ;
        RECT 128.550 47.075 128.720 47.245 ;
        RECT 107.390 46.715 107.560 46.885 ;
        RECT 107.390 46.355 107.560 46.525 ;
        RECT 107.390 45.995 107.560 46.165 ;
        RECT 117.970 46.715 118.140 46.885 ;
        RECT 117.970 46.355 118.140 46.525 ;
        RECT 117.970 45.995 118.140 46.165 ;
        RECT 140.000 47.155 140.170 47.325 ;
        RECT 150.580 47.155 150.750 47.325 ;
        RECT 161.160 68.675 161.330 68.845 ;
        RECT 161.160 68.315 161.330 68.485 ;
        RECT 161.160 67.955 161.330 68.125 ;
        RECT 161.160 63.565 161.330 63.735 ;
        RECT 161.160 63.205 161.330 63.375 ;
        RECT 161.160 62.845 161.330 63.015 ;
        RECT 161.160 62.485 161.330 62.655 ;
        RECT 161.160 58.095 161.330 58.265 ;
        RECT 161.160 57.735 161.330 57.905 ;
        RECT 161.160 57.375 161.330 57.545 ;
        RECT 161.160 57.015 161.330 57.185 ;
        RECT 161.160 52.625 161.330 52.795 ;
        RECT 161.160 52.265 161.330 52.435 ;
        RECT 161.160 51.905 161.330 52.075 ;
        RECT 161.160 51.545 161.330 51.715 ;
        RECT 161.160 47.155 161.330 47.325 ;
        RECT 172.550 68.705 172.720 68.875 ;
        RECT 172.550 68.345 172.720 68.515 ;
        RECT 172.550 67.985 172.720 68.155 ;
        RECT 183.130 68.705 183.300 68.875 ;
        RECT 183.130 68.345 183.300 68.515 ;
        RECT 183.130 67.985 183.300 68.155 ;
        RECT 172.550 63.595 172.720 63.765 ;
        RECT 172.550 63.235 172.720 63.405 ;
        RECT 172.550 62.875 172.720 63.045 ;
        RECT 172.550 62.515 172.720 62.685 ;
        RECT 183.130 63.595 183.300 63.765 ;
        RECT 183.130 63.235 183.300 63.405 ;
        RECT 183.130 62.875 183.300 63.045 ;
        RECT 183.130 62.515 183.300 62.685 ;
        RECT 172.550 58.125 172.720 58.295 ;
        RECT 172.550 57.765 172.720 57.935 ;
        RECT 172.550 57.405 172.720 57.575 ;
        RECT 172.550 57.045 172.720 57.215 ;
        RECT 183.130 58.125 183.300 58.295 ;
        RECT 183.130 57.765 183.300 57.935 ;
        RECT 183.130 57.405 183.300 57.575 ;
        RECT 183.130 57.045 183.300 57.215 ;
        RECT 172.550 52.655 172.720 52.825 ;
        RECT 172.550 52.295 172.720 52.465 ;
        RECT 172.550 51.935 172.720 52.105 ;
        RECT 172.550 51.575 172.720 51.745 ;
        RECT 183.130 52.655 183.300 52.825 ;
        RECT 183.130 52.295 183.300 52.465 ;
        RECT 183.130 51.935 183.300 52.105 ;
        RECT 183.130 51.575 183.300 51.745 ;
        RECT 172.550 47.185 172.720 47.355 ;
        RECT 183.130 47.185 183.300 47.355 ;
        RECT 193.710 68.705 193.880 68.875 ;
        RECT 193.710 68.345 193.880 68.515 ;
        RECT 193.710 67.985 193.880 68.155 ;
        RECT 193.710 63.595 193.880 63.765 ;
        RECT 193.710 63.235 193.880 63.405 ;
        RECT 193.710 62.875 193.880 63.045 ;
        RECT 193.710 62.515 193.880 62.685 ;
        RECT 193.710 58.125 193.880 58.295 ;
        RECT 193.710 57.765 193.880 57.935 ;
        RECT 193.710 57.405 193.880 57.575 ;
        RECT 193.710 57.045 193.880 57.215 ;
        RECT 193.710 52.655 193.880 52.825 ;
        RECT 193.710 52.295 193.880 52.465 ;
        RECT 193.710 51.935 193.880 52.105 ;
        RECT 193.710 51.575 193.880 51.745 ;
        RECT 193.710 47.185 193.880 47.355 ;
        RECT 128.550 46.715 128.720 46.885 ;
        RECT 128.550 46.355 128.720 46.525 ;
        RECT 128.550 45.995 128.720 46.165 ;
        RECT 140.000 46.795 140.170 46.965 ;
        RECT 140.000 46.435 140.170 46.605 ;
        RECT 140.000 46.075 140.170 46.245 ;
        RECT 150.580 46.795 150.750 46.965 ;
        RECT 150.580 46.435 150.750 46.605 ;
        RECT 150.580 46.075 150.750 46.245 ;
        RECT 161.160 46.795 161.330 46.965 ;
        RECT 172.550 46.825 172.720 46.995 ;
        RECT 183.130 46.825 183.300 46.995 ;
        RECT 161.160 46.435 161.330 46.605 ;
        RECT 161.160 46.075 161.330 46.245 ;
        RECT 172.550 46.465 172.720 46.635 ;
        RECT 172.550 46.105 172.720 46.275 ;
        RECT 183.130 46.465 183.300 46.635 ;
        RECT 183.130 46.105 183.300 46.275 ;
        RECT 193.710 46.825 193.880 46.995 ;
        RECT 193.710 46.465 193.880 46.635 ;
        RECT 193.710 46.105 193.880 46.275 ;
        RECT 107.480 39.415 107.650 39.585 ;
        RECT 118.060 39.415 118.230 39.585 ;
        RECT 128.640 39.415 128.810 39.585 ;
        RECT 107.480 39.055 107.650 39.225 ;
        RECT 140.090 39.495 140.260 39.665 ;
        RECT 150.670 39.495 150.840 39.665 ;
        RECT 161.250 39.495 161.420 39.665 ;
        RECT 107.480 38.695 107.650 38.865 ;
        RECT 107.480 38.335 107.650 38.505 ;
        RECT 118.060 39.055 118.230 39.225 ;
        RECT 118.060 38.695 118.230 38.865 ;
        RECT 118.060 38.335 118.230 38.505 ;
        RECT 107.480 33.945 107.650 34.115 ;
        RECT 107.480 33.585 107.650 33.755 ;
        RECT 107.480 33.225 107.650 33.395 ;
        RECT 107.480 32.865 107.650 33.035 ;
        RECT 118.060 33.945 118.230 34.115 ;
        RECT 118.060 33.585 118.230 33.755 ;
        RECT 118.060 33.225 118.230 33.395 ;
        RECT 118.060 32.865 118.230 33.035 ;
        RECT 107.480 28.475 107.650 28.645 ;
        RECT 107.480 28.115 107.650 28.285 ;
        RECT 107.480 27.755 107.650 27.925 ;
        RECT 107.480 27.395 107.650 27.565 ;
        RECT 118.060 28.475 118.230 28.645 ;
        RECT 118.060 28.115 118.230 28.285 ;
        RECT 118.060 27.755 118.230 27.925 ;
        RECT 118.060 27.395 118.230 27.565 ;
        RECT 107.480 23.005 107.650 23.175 ;
        RECT 107.480 22.645 107.650 22.815 ;
        RECT 107.480 22.285 107.650 22.455 ;
        RECT 107.480 21.925 107.650 22.095 ;
        RECT 118.060 23.005 118.230 23.175 ;
        RECT 118.060 22.645 118.230 22.815 ;
        RECT 118.060 22.285 118.230 22.455 ;
        RECT 118.060 21.925 118.230 22.095 ;
        RECT 107.480 17.535 107.650 17.705 ;
        RECT 118.060 17.535 118.230 17.705 ;
        RECT 128.640 39.055 128.810 39.225 ;
        RECT 128.640 38.695 128.810 38.865 ;
        RECT 128.640 38.335 128.810 38.505 ;
        RECT 128.640 33.945 128.810 34.115 ;
        RECT 128.640 33.585 128.810 33.755 ;
        RECT 128.640 33.225 128.810 33.395 ;
        RECT 128.640 32.865 128.810 33.035 ;
        RECT 128.640 28.475 128.810 28.645 ;
        RECT 128.640 28.115 128.810 28.285 ;
        RECT 128.640 27.755 128.810 27.925 ;
        RECT 128.640 27.395 128.810 27.565 ;
        RECT 128.640 23.005 128.810 23.175 ;
        RECT 128.640 22.645 128.810 22.815 ;
        RECT 128.640 22.285 128.810 22.455 ;
        RECT 128.640 21.925 128.810 22.095 ;
        RECT 128.640 17.535 128.810 17.705 ;
        RECT 140.090 39.135 140.260 39.305 ;
        RECT 172.640 39.525 172.810 39.695 ;
        RECT 183.220 39.525 183.390 39.695 ;
        RECT 193.800 39.525 193.970 39.695 ;
        RECT 140.090 38.775 140.260 38.945 ;
        RECT 140.090 38.415 140.260 38.585 ;
        RECT 150.670 39.135 150.840 39.305 ;
        RECT 150.670 38.775 150.840 38.945 ;
        RECT 150.670 38.415 150.840 38.585 ;
        RECT 140.090 34.025 140.260 34.195 ;
        RECT 140.090 33.665 140.260 33.835 ;
        RECT 140.090 33.305 140.260 33.475 ;
        RECT 140.090 32.945 140.260 33.115 ;
        RECT 150.670 34.025 150.840 34.195 ;
        RECT 150.670 33.665 150.840 33.835 ;
        RECT 150.670 33.305 150.840 33.475 ;
        RECT 150.670 32.945 150.840 33.115 ;
        RECT 140.090 28.555 140.260 28.725 ;
        RECT 140.090 28.195 140.260 28.365 ;
        RECT 140.090 27.835 140.260 28.005 ;
        RECT 140.090 27.475 140.260 27.645 ;
        RECT 150.670 28.555 150.840 28.725 ;
        RECT 150.670 28.195 150.840 28.365 ;
        RECT 150.670 27.835 150.840 28.005 ;
        RECT 150.670 27.475 150.840 27.645 ;
        RECT 140.090 23.085 140.260 23.255 ;
        RECT 140.090 22.725 140.260 22.895 ;
        RECT 140.090 22.365 140.260 22.535 ;
        RECT 140.090 22.005 140.260 22.175 ;
        RECT 150.670 23.085 150.840 23.255 ;
        RECT 150.670 22.725 150.840 22.895 ;
        RECT 150.670 22.365 150.840 22.535 ;
        RECT 150.670 22.005 150.840 22.175 ;
        RECT 140.090 17.615 140.260 17.785 ;
        RECT 150.670 17.615 150.840 17.785 ;
        RECT 161.250 39.135 161.420 39.305 ;
        RECT 161.250 38.775 161.420 38.945 ;
        RECT 161.250 38.415 161.420 38.585 ;
        RECT 161.250 34.025 161.420 34.195 ;
        RECT 161.250 33.665 161.420 33.835 ;
        RECT 161.250 33.305 161.420 33.475 ;
        RECT 161.250 32.945 161.420 33.115 ;
        RECT 161.250 28.555 161.420 28.725 ;
        RECT 161.250 28.195 161.420 28.365 ;
        RECT 161.250 27.835 161.420 28.005 ;
        RECT 161.250 27.475 161.420 27.645 ;
        RECT 161.250 23.085 161.420 23.255 ;
        RECT 161.250 22.725 161.420 22.895 ;
        RECT 161.250 22.365 161.420 22.535 ;
        RECT 161.250 22.005 161.420 22.175 ;
        RECT 161.250 17.615 161.420 17.785 ;
        RECT 172.640 39.165 172.810 39.335 ;
        RECT 172.640 38.805 172.810 38.975 ;
        RECT 172.640 38.445 172.810 38.615 ;
        RECT 183.220 39.165 183.390 39.335 ;
        RECT 183.220 38.805 183.390 38.975 ;
        RECT 183.220 38.445 183.390 38.615 ;
        RECT 172.640 34.055 172.810 34.225 ;
        RECT 172.640 33.695 172.810 33.865 ;
        RECT 172.640 33.335 172.810 33.505 ;
        RECT 172.640 32.975 172.810 33.145 ;
        RECT 183.220 34.055 183.390 34.225 ;
        RECT 183.220 33.695 183.390 33.865 ;
        RECT 183.220 33.335 183.390 33.505 ;
        RECT 183.220 32.975 183.390 33.145 ;
        RECT 172.640 28.585 172.810 28.755 ;
        RECT 172.640 28.225 172.810 28.395 ;
        RECT 172.640 27.865 172.810 28.035 ;
        RECT 172.640 27.505 172.810 27.675 ;
        RECT 183.220 28.585 183.390 28.755 ;
        RECT 183.220 28.225 183.390 28.395 ;
        RECT 183.220 27.865 183.390 28.035 ;
        RECT 183.220 27.505 183.390 27.675 ;
        RECT 172.640 23.115 172.810 23.285 ;
        RECT 172.640 22.755 172.810 22.925 ;
        RECT 172.640 22.395 172.810 22.565 ;
        RECT 172.640 22.035 172.810 22.205 ;
        RECT 183.220 23.115 183.390 23.285 ;
        RECT 183.220 22.755 183.390 22.925 ;
        RECT 183.220 22.395 183.390 22.565 ;
        RECT 183.220 22.035 183.390 22.205 ;
        RECT 172.640 17.645 172.810 17.815 ;
        RECT 183.220 17.645 183.390 17.815 ;
        RECT 193.800 39.165 193.970 39.335 ;
        RECT 193.800 38.805 193.970 38.975 ;
        RECT 193.800 38.445 193.970 38.615 ;
        RECT 193.800 34.055 193.970 34.225 ;
        RECT 193.800 33.695 193.970 33.865 ;
        RECT 193.800 33.335 193.970 33.505 ;
        RECT 193.800 32.975 193.970 33.145 ;
        RECT 193.800 28.585 193.970 28.755 ;
        RECT 193.800 28.225 193.970 28.395 ;
        RECT 193.800 27.865 193.970 28.035 ;
        RECT 193.800 27.505 193.970 27.675 ;
        RECT 193.800 23.115 193.970 23.285 ;
        RECT 193.800 22.755 193.970 22.925 ;
        RECT 193.800 22.395 193.970 22.565 ;
        RECT 193.800 22.035 193.970 22.205 ;
        RECT 193.800 17.645 193.970 17.815 ;
        RECT 107.480 17.175 107.650 17.345 ;
        RECT 107.480 16.815 107.650 16.985 ;
        RECT 107.480 16.455 107.650 16.625 ;
        RECT 118.060 17.175 118.230 17.345 ;
        RECT 118.060 16.815 118.230 16.985 ;
        RECT 118.060 16.455 118.230 16.625 ;
        RECT 128.640 17.175 128.810 17.345 ;
        RECT 128.640 16.815 128.810 16.985 ;
        RECT 128.640 16.455 128.810 16.625 ;
        RECT 140.090 17.255 140.260 17.425 ;
        RECT 140.090 16.895 140.260 17.065 ;
        RECT 140.090 16.535 140.260 16.705 ;
        RECT 150.670 17.255 150.840 17.425 ;
        RECT 150.670 16.895 150.840 17.065 ;
        RECT 150.670 16.535 150.840 16.705 ;
        RECT 161.250 17.255 161.420 17.425 ;
        RECT 161.250 16.895 161.420 17.065 ;
        RECT 161.250 16.535 161.420 16.705 ;
        RECT 172.640 17.285 172.810 17.455 ;
        RECT 172.640 16.925 172.810 17.095 ;
        RECT 172.640 16.565 172.810 16.735 ;
        RECT 183.220 17.285 183.390 17.455 ;
        RECT 183.220 16.925 183.390 17.095 ;
        RECT 183.220 16.565 183.390 16.735 ;
        RECT 193.800 17.285 193.970 17.455 ;
        RECT 193.800 16.925 193.970 17.095 ;
        RECT 193.800 16.565 193.970 16.735 ;
      LAYER met1 ;
        RECT 103.290 273.140 104.120 273.360 ;
        RECT 106.770 273.140 108.040 273.190 ;
        RECT 116.390 273.140 117.070 273.900 ;
        RECT 103.290 272.520 117.070 273.140 ;
        RECT 103.290 271.960 104.120 272.520 ;
        RECT 106.770 246.590 108.040 272.520 ;
        RECT 116.390 271.830 117.070 272.520 ;
        RECT -75.965 235.590 -75.735 237.865 ;
        RECT -94.670 235.505 -73.930 235.590 ;
        RECT -96.595 235.205 -73.085 235.505 ;
        RECT -96.595 234.530 -96.385 235.205 ;
        RECT -94.670 235.030 -73.930 235.205 ;
        RECT -94.015 234.530 -93.805 235.030 ;
        RECT -91.445 234.530 -91.235 235.030 ;
        RECT -88.885 234.530 -88.675 235.030 ;
        RECT -86.245 234.530 -86.035 235.030 ;
        RECT -96.595 234.195 -96.360 234.530 ;
        RECT -94.015 234.235 -93.780 234.530 ;
        RECT -91.445 234.235 -91.200 234.530 ;
        RECT -96.590 232.950 -96.360 234.195 ;
        RECT -94.010 232.950 -93.780 234.235 ;
        RECT -91.430 232.950 -91.200 234.235 ;
        RECT -88.885 234.215 -88.620 234.530 ;
        RECT -88.850 232.950 -88.620 234.215 ;
        RECT -86.270 234.195 -86.035 234.530 ;
        RECT -83.705 234.530 -83.495 235.030 ;
        RECT -81.065 234.530 -80.855 235.030 ;
        RECT -78.515 234.530 -78.305 235.030 ;
        RECT -75.955 234.530 -75.745 235.030 ;
        RECT -73.335 234.530 -73.125 235.205 ;
        RECT -86.270 232.950 -86.040 234.195 ;
        RECT -83.705 234.165 -83.460 234.530 ;
        RECT -83.690 232.950 -83.460 234.165 ;
        RECT -81.110 234.065 -80.855 234.530 ;
        RECT -81.110 232.950 -80.880 234.065 ;
        RECT -78.530 232.950 -78.300 234.530 ;
        RECT -75.955 234.105 -75.720 234.530 ;
        RECT -75.950 232.950 -75.720 234.105 ;
        RECT -73.370 234.195 -73.125 234.530 ;
        RECT -73.370 232.950 -73.140 234.195 ;
        RECT -51.150 232.810 -50.920 234.135 ;
        RECT -51.155 231.740 -50.915 232.810 ;
        RECT -48.570 232.730 -48.340 234.135 ;
        RECT -45.990 232.750 -45.760 234.135 ;
        RECT -43.410 232.810 -43.180 234.135 ;
        RECT -48.595 232.555 -48.340 232.730 ;
        RECT -48.595 231.740 -48.355 232.555 ;
        RECT -45.995 231.790 -45.755 232.750 ;
        RECT -43.435 232.555 -43.180 232.810 ;
        RECT -40.830 232.770 -40.600 234.135 ;
        RECT -38.250 232.810 -38.020 234.135 ;
        RECT -40.855 232.555 -40.600 232.770 ;
        RECT -43.435 231.790 -43.195 232.555 ;
        RECT -40.855 231.790 -40.615 232.555 ;
        RECT -38.255 231.790 -38.015 232.810 ;
        RECT -35.670 232.790 -35.440 234.135 ;
        RECT -35.675 231.790 -35.435 232.790 ;
        RECT -33.090 232.730 -32.860 234.135 ;
        RECT -30.510 232.770 -30.280 234.135 ;
        RECT -33.095 231.790 -32.855 232.730 ;
        RECT -30.535 232.555 -30.280 232.770 ;
        RECT -27.930 232.750 -27.700 234.135 ;
        RECT 106.770 233.690 108.170 246.590 ;
        RECT -27.930 232.555 -27.645 232.750 ;
        RECT -30.535 231.790 -30.295 232.555 ;
        RECT -47.690 231.740 -29.860 231.790 ;
        RECT -27.885 231.740 -27.645 232.555 ;
        RECT -51.155 231.440 -27.645 231.740 ;
        RECT -47.690 231.320 -29.860 231.440 ;
        RECT -27.955 229.270 -27.645 231.440 ;
        RECT 105.020 229.710 110.200 233.690 ;
        RECT 106.920 214.730 108.200 229.710 ;
        RECT 107.310 213.740 107.540 214.730 ;
        RECT 117.890 213.740 118.120 215.320 ;
        RECT 128.470 213.740 128.700 215.320 ;
        RECT 139.920 213.820 140.150 215.400 ;
        RECT 150.500 213.820 150.730 215.400 ;
        RECT 161.080 213.820 161.310 215.400 ;
        RECT 172.470 213.850 172.700 215.430 ;
        RECT 183.050 213.850 183.280 215.430 ;
        RECT 193.630 213.850 193.860 215.430 ;
        RECT 107.310 208.270 107.540 209.850 ;
        RECT 117.890 208.270 118.120 209.850 ;
        RECT 128.470 208.270 128.700 209.850 ;
        RECT 139.920 208.350 140.150 209.930 ;
        RECT 150.500 208.350 150.730 209.930 ;
        RECT 161.080 208.350 161.310 209.930 ;
        RECT 172.470 208.380 172.700 209.960 ;
        RECT 183.050 208.380 183.280 209.960 ;
        RECT 193.630 208.380 193.860 209.960 ;
        RECT 107.310 202.800 107.540 204.380 ;
        RECT 117.890 202.800 118.120 204.380 ;
        RECT 128.470 202.800 128.700 204.380 ;
        RECT 139.920 202.880 140.150 204.460 ;
        RECT 150.500 202.880 150.730 204.460 ;
        RECT 161.080 202.880 161.310 204.460 ;
        RECT 172.470 202.910 172.700 204.490 ;
        RECT 183.050 202.910 183.280 204.490 ;
        RECT 193.630 202.910 193.860 204.490 ;
        RECT 107.310 197.330 107.540 198.910 ;
        RECT 117.890 197.330 118.120 198.910 ;
        RECT 128.470 197.330 128.700 198.910 ;
        RECT 139.920 197.410 140.150 198.990 ;
        RECT 150.500 197.410 150.730 198.990 ;
        RECT 161.080 197.410 161.310 198.990 ;
        RECT 172.470 197.440 172.700 199.020 ;
        RECT 183.050 197.440 183.280 199.020 ;
        RECT 193.630 197.440 193.860 199.020 ;
        RECT 107.310 191.860 107.540 193.440 ;
        RECT 117.890 191.860 118.120 193.440 ;
        RECT 128.470 191.860 128.700 193.440 ;
        RECT 139.920 191.940 140.150 193.520 ;
        RECT 150.500 191.940 150.730 193.520 ;
        RECT 161.080 191.940 161.310 193.520 ;
        RECT 172.470 191.970 172.700 193.550 ;
        RECT 183.050 191.970 183.280 193.550 ;
        RECT 193.630 191.970 193.860 193.550 ;
        RECT 107.310 184.660 107.540 186.240 ;
        RECT 117.890 184.660 118.120 186.240 ;
        RECT 128.470 184.660 128.700 186.240 ;
        RECT 139.920 184.740 140.150 186.320 ;
        RECT 150.500 184.740 150.730 186.320 ;
        RECT 161.080 184.740 161.310 186.320 ;
        RECT 172.470 184.770 172.700 186.350 ;
        RECT 183.050 184.770 183.280 186.350 ;
        RECT 193.630 184.770 193.860 186.350 ;
        RECT 107.310 179.190 107.540 180.770 ;
        RECT 117.890 179.190 118.120 180.770 ;
        RECT 128.470 179.190 128.700 180.770 ;
        RECT 139.920 179.270 140.150 180.850 ;
        RECT 150.500 179.270 150.730 180.850 ;
        RECT 161.080 179.270 161.310 180.850 ;
        RECT 172.470 179.300 172.700 180.880 ;
        RECT 183.050 179.300 183.280 180.880 ;
        RECT 193.630 179.300 193.860 180.880 ;
        RECT 107.310 173.720 107.540 175.300 ;
        RECT 117.890 173.720 118.120 175.300 ;
        RECT 128.470 173.720 128.700 175.300 ;
        RECT 139.920 173.800 140.150 175.380 ;
        RECT 150.500 173.800 150.730 175.380 ;
        RECT 161.080 173.800 161.310 175.380 ;
        RECT 172.470 173.830 172.700 175.410 ;
        RECT 183.050 173.830 183.280 175.410 ;
        RECT 193.630 173.830 193.860 175.410 ;
        RECT 107.310 168.250 107.540 169.830 ;
        RECT 117.890 168.250 118.120 169.830 ;
        RECT 128.470 168.250 128.700 169.830 ;
        RECT 139.920 168.330 140.150 169.910 ;
        RECT 150.500 168.330 150.730 169.910 ;
        RECT 161.080 168.330 161.310 169.910 ;
        RECT 172.470 168.360 172.700 169.940 ;
        RECT 183.050 168.360 183.280 169.940 ;
        RECT 193.630 168.360 193.860 169.940 ;
        RECT 107.310 162.780 107.540 164.360 ;
        RECT 117.890 162.780 118.120 164.360 ;
        RECT 128.470 162.780 128.700 164.360 ;
        RECT 139.920 162.860 140.150 164.440 ;
        RECT 150.500 162.860 150.730 164.440 ;
        RECT 161.080 162.860 161.310 164.440 ;
        RECT 172.470 162.890 172.700 164.470 ;
        RECT 183.050 162.890 183.280 164.470 ;
        RECT 193.630 162.890 193.860 164.470 ;
        RECT 107.310 155.490 107.540 157.070 ;
        RECT 117.890 155.490 118.120 157.070 ;
        RECT 128.470 155.490 128.700 157.070 ;
        RECT 139.920 155.570 140.150 157.150 ;
        RECT 150.500 155.570 150.730 157.150 ;
        RECT 161.080 155.570 161.310 157.150 ;
        RECT 172.470 155.600 172.700 157.180 ;
        RECT 183.050 155.600 183.280 157.180 ;
        RECT 193.630 155.600 193.860 157.180 ;
        RECT 107.310 150.020 107.540 151.600 ;
        RECT 117.890 150.020 118.120 151.600 ;
        RECT 128.470 150.020 128.700 151.600 ;
        RECT 139.920 150.100 140.150 151.680 ;
        RECT 150.500 150.100 150.730 151.680 ;
        RECT 161.080 150.100 161.310 151.680 ;
        RECT 172.470 150.130 172.700 151.710 ;
        RECT 183.050 150.130 183.280 151.710 ;
        RECT 193.630 150.130 193.860 151.710 ;
        RECT 107.310 144.550 107.540 146.130 ;
        RECT 117.890 144.550 118.120 146.130 ;
        RECT 128.470 144.550 128.700 146.130 ;
        RECT 139.920 144.630 140.150 146.210 ;
        RECT 150.500 144.630 150.730 146.210 ;
        RECT 161.080 144.630 161.310 146.210 ;
        RECT 172.470 144.660 172.700 146.240 ;
        RECT 183.050 144.660 183.280 146.240 ;
        RECT 193.630 144.660 193.860 146.240 ;
        RECT 107.310 139.080 107.540 140.660 ;
        RECT 117.890 139.080 118.120 140.660 ;
        RECT 128.470 139.080 128.700 140.660 ;
        RECT 139.920 139.160 140.150 140.740 ;
        RECT 150.500 139.160 150.730 140.740 ;
        RECT 161.080 139.160 161.310 140.740 ;
        RECT 172.470 139.190 172.700 140.770 ;
        RECT 183.050 139.190 183.280 140.770 ;
        RECT 193.630 139.190 193.860 140.770 ;
        RECT 107.310 133.610 107.540 135.190 ;
        RECT 117.890 133.610 118.120 135.190 ;
        RECT 128.470 133.610 128.700 135.190 ;
        RECT 139.920 133.690 140.150 135.270 ;
        RECT 150.500 133.690 150.730 135.270 ;
        RECT 161.080 133.690 161.310 135.270 ;
        RECT 172.470 133.720 172.700 135.300 ;
        RECT 183.050 133.720 183.280 135.300 ;
        RECT 193.630 133.720 193.860 135.300 ;
        RECT 107.310 126.310 107.540 127.890 ;
        RECT 117.890 126.310 118.120 127.890 ;
        RECT 128.470 126.310 128.700 127.890 ;
        RECT 139.920 126.390 140.150 127.970 ;
        RECT 150.500 126.390 150.730 127.970 ;
        RECT 161.080 126.390 161.310 127.970 ;
        RECT 172.470 126.420 172.700 128.000 ;
        RECT 183.050 126.420 183.280 128.000 ;
        RECT 193.630 126.420 193.860 128.000 ;
        RECT 107.310 120.840 107.540 122.420 ;
        RECT 117.890 120.840 118.120 122.420 ;
        RECT 128.470 120.840 128.700 122.420 ;
        RECT 139.920 120.920 140.150 122.500 ;
        RECT 150.500 120.920 150.730 122.500 ;
        RECT 161.080 120.920 161.310 122.500 ;
        RECT 172.470 120.950 172.700 122.530 ;
        RECT 183.050 120.950 183.280 122.530 ;
        RECT 193.630 120.950 193.860 122.530 ;
        RECT 107.310 115.370 107.540 116.950 ;
        RECT 117.890 115.370 118.120 116.950 ;
        RECT 128.470 115.370 128.700 116.950 ;
        RECT 139.920 115.450 140.150 117.030 ;
        RECT 150.500 115.450 150.730 117.030 ;
        RECT 161.080 115.450 161.310 117.030 ;
        RECT 172.470 115.480 172.700 117.060 ;
        RECT 183.050 115.480 183.280 117.060 ;
        RECT 193.630 115.480 193.860 117.060 ;
        RECT 107.310 109.900 107.540 111.480 ;
        RECT 117.890 109.900 118.120 111.480 ;
        RECT 128.470 109.900 128.700 111.480 ;
        RECT 139.920 109.980 140.150 111.560 ;
        RECT 150.500 109.980 150.730 111.560 ;
        RECT 161.080 109.980 161.310 111.560 ;
        RECT 172.470 110.010 172.700 111.590 ;
        RECT 183.050 110.010 183.280 111.590 ;
        RECT 193.630 110.010 193.860 111.590 ;
        RECT 107.310 104.430 107.540 106.010 ;
        RECT 117.890 104.430 118.120 106.010 ;
        RECT 128.470 104.430 128.700 106.010 ;
        RECT 139.920 104.510 140.150 106.090 ;
        RECT 150.500 104.510 150.730 106.090 ;
        RECT 161.080 104.510 161.310 106.090 ;
        RECT 172.470 104.540 172.700 106.120 ;
        RECT 183.050 104.540 183.280 106.120 ;
        RECT 193.630 104.540 193.860 106.120 ;
        RECT 107.310 96.990 107.540 98.570 ;
        RECT 117.890 96.990 118.120 98.570 ;
        RECT 128.470 96.990 128.700 98.570 ;
        RECT 139.920 97.070 140.150 98.650 ;
        RECT 150.500 97.070 150.730 98.650 ;
        RECT 161.080 97.070 161.310 98.650 ;
        RECT 172.470 97.100 172.700 98.680 ;
        RECT 183.050 97.100 183.280 98.680 ;
        RECT 193.630 97.100 193.860 98.680 ;
        RECT 107.310 91.520 107.540 93.100 ;
        RECT 117.890 91.520 118.120 93.100 ;
        RECT 128.470 91.520 128.700 93.100 ;
        RECT 139.920 91.600 140.150 93.180 ;
        RECT 150.500 91.600 150.730 93.180 ;
        RECT 161.080 91.600 161.310 93.180 ;
        RECT 172.470 91.630 172.700 93.210 ;
        RECT 183.050 91.630 183.280 93.210 ;
        RECT 193.630 91.630 193.860 93.210 ;
        RECT 107.310 86.050 107.540 87.630 ;
        RECT 117.890 86.050 118.120 87.630 ;
        RECT 128.470 86.050 128.700 87.630 ;
        RECT 139.920 86.130 140.150 87.710 ;
        RECT 150.500 86.130 150.730 87.710 ;
        RECT 161.080 86.130 161.310 87.710 ;
        RECT 172.470 86.160 172.700 87.740 ;
        RECT 183.050 86.160 183.280 87.740 ;
        RECT 193.630 86.160 193.860 87.740 ;
        RECT 107.310 80.580 107.540 82.160 ;
        RECT 117.890 80.580 118.120 82.160 ;
        RECT 128.470 80.580 128.700 82.160 ;
        RECT 139.920 80.660 140.150 82.240 ;
        RECT 150.500 80.660 150.730 82.240 ;
        RECT 161.080 80.660 161.310 82.240 ;
        RECT 172.470 80.690 172.700 82.270 ;
        RECT 183.050 80.690 183.280 82.270 ;
        RECT 193.630 80.690 193.860 82.270 ;
        RECT 107.310 75.110 107.540 76.690 ;
        RECT 117.890 75.110 118.120 76.690 ;
        RECT 128.470 75.110 128.700 76.690 ;
        RECT 139.920 75.190 140.150 76.770 ;
        RECT 150.500 75.190 150.730 76.770 ;
        RECT 161.080 75.190 161.310 76.770 ;
        RECT 172.470 75.220 172.700 76.800 ;
        RECT 183.050 75.220 183.280 76.800 ;
        RECT 193.630 75.220 193.860 76.800 ;
        RECT 107.360 67.710 107.590 69.290 ;
        RECT 117.940 67.710 118.170 69.290 ;
        RECT 128.520 67.710 128.750 69.290 ;
        RECT 139.970 67.790 140.200 69.370 ;
        RECT 150.550 67.790 150.780 69.370 ;
        RECT 161.130 67.790 161.360 69.370 ;
        RECT 172.520 67.820 172.750 69.400 ;
        RECT 183.100 67.820 183.330 69.400 ;
        RECT 193.680 67.820 193.910 69.400 ;
        RECT 107.360 62.240 107.590 63.820 ;
        RECT 117.940 62.240 118.170 63.820 ;
        RECT 128.520 62.240 128.750 63.820 ;
        RECT 139.970 62.320 140.200 63.900 ;
        RECT 150.550 62.320 150.780 63.900 ;
        RECT 161.130 62.320 161.360 63.900 ;
        RECT 172.520 62.350 172.750 63.930 ;
        RECT 183.100 62.350 183.330 63.930 ;
        RECT 193.680 62.350 193.910 63.930 ;
        RECT 107.360 56.770 107.590 58.350 ;
        RECT 117.940 56.770 118.170 58.350 ;
        RECT 128.520 56.770 128.750 58.350 ;
        RECT 139.970 56.850 140.200 58.430 ;
        RECT 150.550 56.850 150.780 58.430 ;
        RECT 161.130 56.850 161.360 58.430 ;
        RECT 172.520 56.880 172.750 58.460 ;
        RECT 183.100 56.880 183.330 58.460 ;
        RECT 193.680 56.880 193.910 58.460 ;
        RECT 107.360 51.300 107.590 52.880 ;
        RECT 117.940 51.300 118.170 52.880 ;
        RECT 128.520 51.300 128.750 52.880 ;
        RECT 139.970 51.380 140.200 52.960 ;
        RECT 150.550 51.380 150.780 52.960 ;
        RECT 161.130 51.380 161.360 52.960 ;
        RECT 172.520 51.410 172.750 52.990 ;
        RECT 183.100 51.410 183.330 52.990 ;
        RECT 193.680 51.410 193.910 52.990 ;
        RECT 107.360 45.830 107.590 47.410 ;
        RECT 117.940 45.830 118.170 47.410 ;
        RECT 128.520 45.830 128.750 47.410 ;
        RECT 139.970 45.910 140.200 47.490 ;
        RECT 150.550 45.910 150.780 47.490 ;
        RECT 161.130 45.910 161.360 47.490 ;
        RECT 172.520 45.940 172.750 47.520 ;
        RECT 183.100 45.940 183.330 47.520 ;
        RECT 193.680 45.940 193.910 47.520 ;
        RECT 107.450 38.170 107.680 39.750 ;
        RECT 118.030 38.170 118.260 39.750 ;
        RECT 128.610 38.170 128.840 39.750 ;
        RECT 140.060 38.250 140.290 39.830 ;
        RECT 150.640 38.250 150.870 39.830 ;
        RECT 161.220 38.250 161.450 39.830 ;
        RECT 172.610 38.280 172.840 39.860 ;
        RECT 183.190 38.280 183.420 39.860 ;
        RECT 193.770 38.280 194.000 39.860 ;
        RECT 107.450 32.700 107.680 34.280 ;
        RECT 118.030 32.700 118.260 34.280 ;
        RECT 128.610 32.700 128.840 34.280 ;
        RECT 140.060 32.780 140.290 34.360 ;
        RECT 150.640 32.780 150.870 34.360 ;
        RECT 161.220 32.780 161.450 34.360 ;
        RECT 172.610 32.810 172.840 34.390 ;
        RECT 183.190 32.810 183.420 34.390 ;
        RECT 193.770 32.810 194.000 34.390 ;
        RECT 107.450 27.230 107.680 28.810 ;
        RECT 118.030 27.230 118.260 28.810 ;
        RECT 128.610 27.230 128.840 28.810 ;
        RECT 140.060 27.310 140.290 28.890 ;
        RECT 150.640 27.310 150.870 28.890 ;
        RECT 161.220 27.310 161.450 28.890 ;
        RECT 172.610 27.340 172.840 28.920 ;
        RECT 183.190 27.340 183.420 28.920 ;
        RECT 193.770 27.340 194.000 28.920 ;
        RECT 107.450 21.760 107.680 23.340 ;
        RECT 118.030 21.760 118.260 23.340 ;
        RECT 128.610 21.760 128.840 23.340 ;
        RECT 140.060 21.840 140.290 23.420 ;
        RECT 150.640 21.840 150.870 23.420 ;
        RECT 161.220 21.840 161.450 23.420 ;
        RECT 172.610 21.870 172.840 23.450 ;
        RECT 183.190 21.870 183.420 23.450 ;
        RECT 193.770 21.870 194.000 23.450 ;
        RECT 107.450 16.290 107.680 17.870 ;
        RECT 118.030 16.290 118.260 17.870 ;
        RECT 128.610 16.290 128.840 17.870 ;
        RECT 140.060 16.370 140.290 17.950 ;
        RECT 150.640 16.370 150.870 17.950 ;
        RECT 161.220 16.370 161.450 17.950 ;
        RECT 172.610 16.400 172.840 17.980 ;
        RECT 183.190 16.400 183.420 17.980 ;
        RECT 193.770 16.400 194.000 17.980 ;
      LAYER via ;
        RECT -94.510 235.180 -94.250 235.440 ;
        RECT -94.190 235.180 -93.930 235.440 ;
        RECT -93.870 235.180 -93.610 235.440 ;
        RECT -93.550 235.180 -93.290 235.440 ;
        RECT -93.230 235.180 -92.970 235.440 ;
        RECT -92.910 235.180 -92.650 235.440 ;
        RECT -92.590 235.180 -92.330 235.440 ;
        RECT -92.270 235.180 -92.010 235.440 ;
        RECT -91.950 235.180 -91.690 235.440 ;
        RECT -91.630 235.180 -91.370 235.440 ;
        RECT -91.310 235.180 -91.050 235.440 ;
        RECT -90.990 235.180 -90.730 235.440 ;
        RECT -90.670 235.180 -90.410 235.440 ;
        RECT -90.350 235.180 -90.090 235.440 ;
        RECT -90.030 235.180 -89.770 235.440 ;
        RECT -89.710 235.180 -89.450 235.440 ;
        RECT -89.390 235.180 -89.130 235.440 ;
        RECT -89.070 235.180 -88.810 235.440 ;
        RECT -88.750 235.180 -88.490 235.440 ;
        RECT -88.430 235.180 -88.170 235.440 ;
        RECT -88.110 235.180 -87.850 235.440 ;
        RECT -87.790 235.180 -87.530 235.440 ;
        RECT -87.470 235.180 -87.210 235.440 ;
        RECT -87.150 235.180 -86.890 235.440 ;
        RECT -86.830 235.180 -86.570 235.440 ;
        RECT -86.510 235.180 -86.250 235.440 ;
        RECT -86.190 235.180 -85.930 235.440 ;
        RECT -85.870 235.180 -85.610 235.440 ;
        RECT -85.550 235.180 -85.290 235.440 ;
        RECT -85.230 235.180 -84.970 235.440 ;
        RECT -84.910 235.180 -84.650 235.440 ;
        RECT -84.590 235.180 -84.330 235.440 ;
        RECT -84.270 235.180 -84.010 235.440 ;
        RECT -83.950 235.180 -83.690 235.440 ;
        RECT -83.630 235.180 -83.370 235.440 ;
        RECT -83.310 235.180 -83.050 235.440 ;
        RECT -82.990 235.180 -82.730 235.440 ;
        RECT -82.670 235.180 -82.410 235.440 ;
        RECT -82.350 235.180 -82.090 235.440 ;
        RECT -82.030 235.180 -81.770 235.440 ;
        RECT -81.710 235.180 -81.450 235.440 ;
        RECT -81.390 235.180 -81.130 235.440 ;
        RECT -81.070 235.180 -80.810 235.440 ;
        RECT -80.750 235.180 -80.490 235.440 ;
        RECT -80.430 235.180 -80.170 235.440 ;
        RECT -80.110 235.180 -79.850 235.440 ;
        RECT -79.790 235.180 -79.530 235.440 ;
        RECT -79.470 235.180 -79.210 235.440 ;
        RECT -79.150 235.180 -78.890 235.440 ;
        RECT -78.830 235.180 -78.570 235.440 ;
        RECT -78.510 235.180 -78.250 235.440 ;
        RECT -78.190 235.180 -77.930 235.440 ;
        RECT -77.870 235.180 -77.610 235.440 ;
        RECT -77.550 235.180 -77.290 235.440 ;
        RECT -77.230 235.180 -76.970 235.440 ;
        RECT -76.910 235.180 -76.650 235.440 ;
        RECT -76.590 235.180 -76.330 235.440 ;
        RECT -76.270 235.180 -76.010 235.440 ;
        RECT -75.950 235.180 -75.690 235.440 ;
        RECT -75.630 235.180 -75.370 235.440 ;
        RECT -75.310 235.180 -75.050 235.440 ;
        RECT -74.990 235.180 -74.730 235.440 ;
        RECT -74.670 235.180 -74.410 235.440 ;
        RECT -74.350 235.180 -74.090 235.440 ;
        RECT -47.545 231.425 -47.285 231.685 ;
        RECT -47.225 231.425 -46.965 231.685 ;
        RECT -46.905 231.425 -46.645 231.685 ;
        RECT -46.585 231.425 -46.325 231.685 ;
        RECT -46.265 231.425 -46.005 231.685 ;
        RECT -45.945 231.425 -45.685 231.685 ;
        RECT -45.625 231.425 -45.365 231.685 ;
        RECT -45.305 231.425 -45.045 231.685 ;
        RECT -44.985 231.425 -44.725 231.685 ;
        RECT -44.665 231.425 -44.405 231.685 ;
        RECT -44.345 231.425 -44.085 231.685 ;
        RECT -44.025 231.425 -43.765 231.685 ;
        RECT -43.705 231.425 -43.445 231.685 ;
        RECT -43.385 231.425 -43.125 231.685 ;
        RECT -43.065 231.425 -42.805 231.685 ;
        RECT -42.745 231.425 -42.485 231.685 ;
        RECT -42.425 231.425 -42.165 231.685 ;
        RECT -42.105 231.425 -41.845 231.685 ;
        RECT -41.785 231.425 -41.525 231.685 ;
        RECT -41.465 231.425 -41.205 231.685 ;
        RECT -41.145 231.425 -40.885 231.685 ;
        RECT -40.825 231.425 -40.565 231.685 ;
        RECT -40.505 231.425 -40.245 231.685 ;
        RECT -40.185 231.425 -39.925 231.685 ;
        RECT -39.865 231.425 -39.605 231.685 ;
        RECT -39.545 231.425 -39.285 231.685 ;
        RECT -39.225 231.425 -38.965 231.685 ;
        RECT -38.905 231.425 -38.645 231.685 ;
        RECT -38.585 231.425 -38.325 231.685 ;
        RECT -38.265 231.425 -38.005 231.685 ;
        RECT -37.945 231.425 -37.685 231.685 ;
        RECT -37.625 231.425 -37.365 231.685 ;
        RECT -37.305 231.425 -37.045 231.685 ;
        RECT -36.985 231.425 -36.725 231.685 ;
        RECT -36.665 231.425 -36.405 231.685 ;
        RECT -36.345 231.425 -36.085 231.685 ;
        RECT -36.025 231.425 -35.765 231.685 ;
        RECT -35.705 231.425 -35.445 231.685 ;
        RECT -35.385 231.425 -35.125 231.685 ;
        RECT -35.065 231.425 -34.805 231.685 ;
        RECT -34.745 231.425 -34.485 231.685 ;
        RECT -34.425 231.425 -34.165 231.685 ;
        RECT -34.105 231.425 -33.845 231.685 ;
        RECT -33.785 231.425 -33.525 231.685 ;
        RECT -33.465 231.425 -33.205 231.685 ;
        RECT -33.145 231.425 -32.885 231.685 ;
        RECT -32.825 231.425 -32.565 231.685 ;
        RECT -32.505 231.425 -32.245 231.685 ;
        RECT -32.185 231.425 -31.925 231.685 ;
        RECT -31.865 231.425 -31.605 231.685 ;
        RECT -31.545 231.425 -31.285 231.685 ;
        RECT -31.225 231.425 -30.965 231.685 ;
        RECT -30.905 231.425 -30.645 231.685 ;
        RECT -30.585 231.425 -30.325 231.685 ;
        RECT -30.265 231.425 -30.005 231.685 ;
        RECT 105.080 229.810 110.140 233.590 ;
      LAYER met2 ;
        RECT -94.620 235.640 -92.530 235.710 ;
        RECT -60.330 235.700 -57.090 235.890 ;
        RECT -74.950 235.640 -57.090 235.700 ;
        RECT -94.620 235.020 -57.090 235.640 ;
        RECT -94.620 234.980 -73.980 235.020 ;
        RECT -94.620 234.910 -92.530 234.980 ;
        RECT -60.330 234.960 -57.090 235.020 ;
        RECT -57.840 231.960 -57.210 234.960 ;
        RECT 105.070 232.470 110.150 233.740 ;
        RECT -57.840 231.840 -42.260 231.960 ;
        RECT -10.930 231.870 110.150 232.470 ;
        RECT -30.820 231.840 110.150 231.870 ;
        RECT -57.840 231.290 110.150 231.840 ;
        RECT -57.840 231.280 -29.910 231.290 ;
        RECT -47.640 231.270 -29.910 231.280 ;
        RECT -10.930 230.930 110.150 231.290 ;
        RECT 105.070 229.660 110.150 230.930 ;
      LAYER via2 ;
        RECT -94.515 234.970 -92.635 235.650 ;
      LAYER met3 ;
        RECT -130.110 235.685 -93.600 236.100 ;
        RECT -130.110 234.935 -92.480 235.685 ;
        RECT -130.110 233.840 -93.600 234.935 ;
    END
  END vout
  PIN va
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13125.000000 ;
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER li1 ;
        RECT -95.870 220.830 -95.700 222.450 ;
        RECT -93.290 220.830 -93.120 222.450 ;
        RECT -90.710 220.830 -90.540 222.450 ;
        RECT -88.130 220.830 -87.960 222.450 ;
        RECT -85.550 220.830 -85.380 222.450 ;
        RECT -82.970 220.830 -82.800 222.450 ;
        RECT -80.390 220.830 -80.220 222.450 ;
        RECT -77.810 220.830 -77.640 222.450 ;
        RECT -75.230 220.830 -75.060 222.450 ;
        RECT -72.650 220.830 -72.480 222.450 ;
        RECT -51.010 220.385 -50.840 222.005 ;
        RECT -48.430 220.385 -48.260 222.005 ;
        RECT -45.850 220.385 -45.680 222.005 ;
        RECT -43.270 220.385 -43.100 222.005 ;
        RECT -40.690 220.385 -40.520 222.005 ;
        RECT -38.110 220.385 -37.940 222.005 ;
        RECT -35.530 220.385 -35.360 222.005 ;
        RECT -32.950 220.385 -32.780 222.005 ;
        RECT -30.370 220.385 -30.200 222.005 ;
        RECT -27.790 220.385 -27.620 222.005 ;
        RECT 99.540 220.030 101.480 220.170 ;
        RECT 105.350 220.030 120.110 220.040 ;
        RECT 99.540 219.750 120.110 220.030 ;
        RECT 99.540 219.080 122.550 219.750 ;
        RECT 99.540 219.070 114.550 219.080 ;
        RECT 99.540 218.390 101.480 219.070 ;
        RECT 119.600 217.820 122.550 219.080 ;
      LAYER mcon ;
        RECT -95.870 222.095 -95.700 222.265 ;
        RECT -95.870 221.735 -95.700 221.905 ;
        RECT -95.870 221.375 -95.700 221.545 ;
        RECT -95.870 221.015 -95.700 221.185 ;
        RECT -93.290 222.095 -93.120 222.265 ;
        RECT -93.290 221.735 -93.120 221.905 ;
        RECT -93.290 221.375 -93.120 221.545 ;
        RECT -93.290 221.015 -93.120 221.185 ;
        RECT -90.710 222.095 -90.540 222.265 ;
        RECT -90.710 221.735 -90.540 221.905 ;
        RECT -90.710 221.375 -90.540 221.545 ;
        RECT -90.710 221.015 -90.540 221.185 ;
        RECT -88.130 222.095 -87.960 222.265 ;
        RECT -88.130 221.735 -87.960 221.905 ;
        RECT -88.130 221.375 -87.960 221.545 ;
        RECT -88.130 221.015 -87.960 221.185 ;
        RECT -85.550 222.095 -85.380 222.265 ;
        RECT -85.550 221.735 -85.380 221.905 ;
        RECT -85.550 221.375 -85.380 221.545 ;
        RECT -85.550 221.015 -85.380 221.185 ;
        RECT -82.970 222.095 -82.800 222.265 ;
        RECT -82.970 221.735 -82.800 221.905 ;
        RECT -82.970 221.375 -82.800 221.545 ;
        RECT -82.970 221.015 -82.800 221.185 ;
        RECT -80.390 222.095 -80.220 222.265 ;
        RECT -80.390 221.735 -80.220 221.905 ;
        RECT -80.390 221.375 -80.220 221.545 ;
        RECT -80.390 221.015 -80.220 221.185 ;
        RECT -77.810 222.095 -77.640 222.265 ;
        RECT -77.810 221.735 -77.640 221.905 ;
        RECT -77.810 221.375 -77.640 221.545 ;
        RECT -77.810 221.015 -77.640 221.185 ;
        RECT -75.230 222.095 -75.060 222.265 ;
        RECT -75.230 221.735 -75.060 221.905 ;
        RECT -75.230 221.375 -75.060 221.545 ;
        RECT -75.230 221.015 -75.060 221.185 ;
        RECT -72.650 222.095 -72.480 222.265 ;
        RECT -72.650 221.735 -72.480 221.905 ;
        RECT -72.650 221.375 -72.480 221.545 ;
        RECT -72.650 221.015 -72.480 221.185 ;
        RECT -51.010 221.650 -50.840 221.820 ;
        RECT -51.010 221.290 -50.840 221.460 ;
        RECT -51.010 220.930 -50.840 221.100 ;
        RECT -51.010 220.570 -50.840 220.740 ;
        RECT -48.430 221.650 -48.260 221.820 ;
        RECT -48.430 221.290 -48.260 221.460 ;
        RECT -48.430 220.930 -48.260 221.100 ;
        RECT -48.430 220.570 -48.260 220.740 ;
        RECT -45.850 221.650 -45.680 221.820 ;
        RECT -45.850 221.290 -45.680 221.460 ;
        RECT -45.850 220.930 -45.680 221.100 ;
        RECT -45.850 220.570 -45.680 220.740 ;
        RECT -43.270 221.650 -43.100 221.820 ;
        RECT -43.270 221.290 -43.100 221.460 ;
        RECT -43.270 220.930 -43.100 221.100 ;
        RECT -43.270 220.570 -43.100 220.740 ;
        RECT -40.690 221.650 -40.520 221.820 ;
        RECT -40.690 221.290 -40.520 221.460 ;
        RECT -40.690 220.930 -40.520 221.100 ;
        RECT -40.690 220.570 -40.520 220.740 ;
        RECT -38.110 221.650 -37.940 221.820 ;
        RECT -38.110 221.290 -37.940 221.460 ;
        RECT -38.110 220.930 -37.940 221.100 ;
        RECT -38.110 220.570 -37.940 220.740 ;
        RECT -35.530 221.650 -35.360 221.820 ;
        RECT -35.530 221.290 -35.360 221.460 ;
        RECT -35.530 220.930 -35.360 221.100 ;
        RECT -35.530 220.570 -35.360 220.740 ;
        RECT -32.950 221.650 -32.780 221.820 ;
        RECT -32.950 221.290 -32.780 221.460 ;
        RECT -32.950 220.930 -32.780 221.100 ;
        RECT -32.950 220.570 -32.780 220.740 ;
        RECT -30.370 221.650 -30.200 221.820 ;
        RECT -30.370 221.290 -30.200 221.460 ;
        RECT -30.370 220.930 -30.200 221.100 ;
        RECT -30.370 220.570 -30.200 220.740 ;
        RECT -27.790 221.650 -27.620 221.820 ;
        RECT -27.790 221.290 -27.620 221.460 ;
        RECT -27.790 220.930 -27.620 221.100 ;
        RECT -27.790 220.570 -27.620 220.740 ;
        RECT 99.705 218.475 101.315 220.085 ;
        RECT 119.960 217.975 121.930 219.585 ;
      LAYER met1 ;
        RECT -75.275 223.530 -75.045 225.765 ;
        RECT -96.030 223.020 -72.230 223.530 ;
        RECT -95.905 222.430 -95.695 223.020 ;
        RECT -93.325 222.430 -93.115 223.020 ;
        RECT -90.755 222.430 -90.545 223.020 ;
        RECT -88.195 222.430 -87.985 223.020 ;
        RECT -85.555 222.430 -85.345 223.020 ;
        RECT -95.905 222.095 -95.670 222.430 ;
        RECT -93.325 222.135 -93.090 222.430 ;
        RECT -90.755 222.135 -90.510 222.430 ;
        RECT -95.900 220.850 -95.670 222.095 ;
        RECT -93.320 220.850 -93.090 222.135 ;
        RECT -90.740 220.850 -90.510 222.135 ;
        RECT -88.195 222.115 -87.930 222.430 ;
        RECT -88.160 220.850 -87.930 222.115 ;
        RECT -85.580 222.095 -85.345 222.430 ;
        RECT -83.015 222.430 -82.805 223.020 ;
        RECT -80.375 222.430 -80.165 223.020 ;
        RECT -77.825 222.430 -77.615 223.020 ;
        RECT -75.275 222.985 -75.045 223.020 ;
        RECT -75.265 222.430 -75.055 222.985 ;
        RECT -72.645 222.430 -72.435 223.020 ;
        RECT -85.580 220.850 -85.350 222.095 ;
        RECT -83.015 222.065 -82.770 222.430 ;
        RECT -83.000 220.850 -82.770 222.065 ;
        RECT -80.420 221.965 -80.165 222.430 ;
        RECT -80.420 220.850 -80.190 221.965 ;
        RECT -77.840 220.850 -77.610 222.430 ;
        RECT -75.265 222.005 -75.030 222.430 ;
        RECT -75.260 220.850 -75.030 222.005 ;
        RECT -72.680 222.095 -72.435 222.430 ;
        RECT -72.680 220.850 -72.450 222.095 ;
        RECT -51.040 220.660 -50.810 221.985 ;
        RECT -51.045 219.590 -50.805 220.660 ;
        RECT -48.460 220.580 -48.230 221.985 ;
        RECT -45.880 220.600 -45.650 221.985 ;
        RECT -43.300 220.660 -43.070 221.985 ;
        RECT -48.485 220.405 -48.230 220.580 ;
        RECT -48.485 219.630 -48.245 220.405 ;
        RECT -45.885 219.630 -45.645 220.600 ;
        RECT -43.325 220.405 -43.070 220.660 ;
        RECT -40.720 220.620 -40.490 221.985 ;
        RECT -38.140 220.660 -37.910 221.985 ;
        RECT -40.745 220.405 -40.490 220.620 ;
        RECT -43.325 219.630 -43.085 220.405 ;
        RECT -40.745 219.630 -40.505 220.405 ;
        RECT -38.145 219.630 -37.905 220.660 ;
        RECT -35.560 220.640 -35.330 221.985 ;
        RECT -35.565 219.630 -35.325 220.640 ;
        RECT -32.980 220.580 -32.750 221.985 ;
        RECT -30.400 220.620 -30.170 221.985 ;
        RECT -32.985 219.630 -32.745 220.580 ;
        RECT -30.425 220.405 -30.170 220.620 ;
        RECT -27.820 220.600 -27.590 221.985 ;
        RECT -27.820 220.405 -27.535 220.600 ;
        RECT -30.425 219.630 -30.185 220.405 ;
        RECT -27.775 219.630 -27.535 220.405 ;
        RECT -49.970 219.590 -27.160 219.630 ;
        RECT -51.045 219.290 -27.160 219.590 ;
        RECT -49.970 219.070 -27.160 219.290 ;
        RECT -27.845 217.120 -27.535 219.070 ;
        RECT 99.480 218.360 101.540 220.200 ;
        RECT 119.600 217.820 122.550 219.750 ;
      LAYER via ;
        RECT -95.940 223.145 -95.680 223.405 ;
        RECT -95.620 223.145 -95.360 223.405 ;
        RECT -95.300 223.145 -95.040 223.405 ;
        RECT -94.980 223.145 -94.720 223.405 ;
        RECT -94.660 223.145 -94.400 223.405 ;
        RECT -94.340 223.145 -94.080 223.405 ;
        RECT -94.020 223.145 -93.760 223.405 ;
        RECT -93.700 223.145 -93.440 223.405 ;
        RECT -93.380 223.145 -93.120 223.405 ;
        RECT -93.060 223.145 -92.800 223.405 ;
        RECT -92.740 223.145 -92.480 223.405 ;
        RECT -92.420 223.145 -92.160 223.405 ;
        RECT -92.100 223.145 -91.840 223.405 ;
        RECT -91.780 223.145 -91.520 223.405 ;
        RECT -91.460 223.145 -91.200 223.405 ;
        RECT -91.140 223.145 -90.880 223.405 ;
        RECT -90.820 223.145 -90.560 223.405 ;
        RECT -90.500 223.145 -90.240 223.405 ;
        RECT -90.180 223.145 -89.920 223.405 ;
        RECT -89.860 223.145 -89.600 223.405 ;
        RECT -89.540 223.145 -89.280 223.405 ;
        RECT -89.220 223.145 -88.960 223.405 ;
        RECT -88.900 223.145 -88.640 223.405 ;
        RECT -88.580 223.145 -88.320 223.405 ;
        RECT -88.260 223.145 -88.000 223.405 ;
        RECT -87.940 223.145 -87.680 223.405 ;
        RECT -87.620 223.145 -87.360 223.405 ;
        RECT -87.300 223.145 -87.040 223.405 ;
        RECT -86.980 223.145 -86.720 223.405 ;
        RECT -86.660 223.145 -86.400 223.405 ;
        RECT -86.340 223.145 -86.080 223.405 ;
        RECT -86.020 223.145 -85.760 223.405 ;
        RECT -85.700 223.145 -85.440 223.405 ;
        RECT -85.380 223.145 -85.120 223.405 ;
        RECT -85.060 223.145 -84.800 223.405 ;
        RECT -84.740 223.145 -84.480 223.405 ;
        RECT -84.420 223.145 -84.160 223.405 ;
        RECT -84.100 223.145 -83.840 223.405 ;
        RECT -83.780 223.145 -83.520 223.405 ;
        RECT -83.460 223.145 -83.200 223.405 ;
        RECT -83.140 223.145 -82.880 223.405 ;
        RECT -82.820 223.145 -82.560 223.405 ;
        RECT -82.500 223.145 -82.240 223.405 ;
        RECT -82.180 223.145 -81.920 223.405 ;
        RECT -81.860 223.145 -81.600 223.405 ;
        RECT -81.540 223.145 -81.280 223.405 ;
        RECT -81.220 223.145 -80.960 223.405 ;
        RECT -80.900 223.145 -80.640 223.405 ;
        RECT -80.580 223.145 -80.320 223.405 ;
        RECT -80.260 223.145 -80.000 223.405 ;
        RECT -79.940 223.145 -79.680 223.405 ;
        RECT -79.620 223.145 -79.360 223.405 ;
        RECT -79.300 223.145 -79.040 223.405 ;
        RECT -78.980 223.145 -78.720 223.405 ;
        RECT -78.660 223.145 -78.400 223.405 ;
        RECT -78.340 223.145 -78.080 223.405 ;
        RECT -78.020 223.145 -77.760 223.405 ;
        RECT -77.700 223.145 -77.440 223.405 ;
        RECT -77.380 223.145 -77.120 223.405 ;
        RECT -77.060 223.145 -76.800 223.405 ;
        RECT -76.740 223.145 -76.480 223.405 ;
        RECT -76.420 223.145 -76.160 223.405 ;
        RECT -76.100 223.145 -75.840 223.405 ;
        RECT -75.780 223.145 -75.520 223.405 ;
        RECT -75.460 223.145 -75.200 223.405 ;
        RECT -75.140 223.145 -74.880 223.405 ;
        RECT -74.820 223.145 -74.560 223.405 ;
        RECT -74.500 223.145 -74.240 223.405 ;
        RECT -74.180 223.145 -73.920 223.405 ;
        RECT -73.860 223.145 -73.600 223.405 ;
        RECT -73.540 223.145 -73.280 223.405 ;
        RECT -73.220 223.145 -72.960 223.405 ;
        RECT -72.900 223.145 -72.640 223.405 ;
        RECT -72.580 223.145 -72.320 223.405 ;
        RECT -49.895 219.220 -49.635 219.480 ;
        RECT -49.575 219.220 -49.315 219.480 ;
        RECT -49.255 219.220 -48.995 219.480 ;
        RECT -48.935 219.220 -48.675 219.480 ;
        RECT -48.615 219.220 -48.355 219.480 ;
        RECT -48.295 219.220 -48.035 219.480 ;
        RECT -47.975 219.220 -47.715 219.480 ;
        RECT -47.655 219.220 -47.395 219.480 ;
        RECT -47.335 219.220 -47.075 219.480 ;
        RECT -47.015 219.220 -46.755 219.480 ;
        RECT -46.695 219.220 -46.435 219.480 ;
        RECT -46.375 219.220 -46.115 219.480 ;
        RECT -46.055 219.220 -45.795 219.480 ;
        RECT -45.735 219.220 -45.475 219.480 ;
        RECT -45.415 219.220 -45.155 219.480 ;
        RECT -45.095 219.220 -44.835 219.480 ;
        RECT -44.775 219.220 -44.515 219.480 ;
        RECT -44.455 219.220 -44.195 219.480 ;
        RECT -44.135 219.220 -43.875 219.480 ;
        RECT -43.815 219.220 -43.555 219.480 ;
        RECT -43.495 219.220 -43.235 219.480 ;
        RECT -43.175 219.220 -42.915 219.480 ;
        RECT -42.855 219.220 -42.595 219.480 ;
        RECT -42.535 219.220 -42.275 219.480 ;
        RECT -42.215 219.220 -41.955 219.480 ;
        RECT -41.895 219.220 -41.635 219.480 ;
        RECT -41.575 219.220 -41.315 219.480 ;
        RECT -41.255 219.220 -40.995 219.480 ;
        RECT -40.935 219.220 -40.675 219.480 ;
        RECT -40.615 219.220 -40.355 219.480 ;
        RECT -40.295 219.220 -40.035 219.480 ;
        RECT -39.975 219.220 -39.715 219.480 ;
        RECT -39.655 219.220 -39.395 219.480 ;
        RECT -39.335 219.220 -39.075 219.480 ;
        RECT -39.015 219.220 -38.755 219.480 ;
        RECT -38.695 219.220 -38.435 219.480 ;
        RECT -38.375 219.220 -38.115 219.480 ;
        RECT -38.055 219.220 -37.795 219.480 ;
        RECT -37.735 219.220 -37.475 219.480 ;
        RECT -37.415 219.220 -37.155 219.480 ;
        RECT -37.095 219.220 -36.835 219.480 ;
        RECT -36.775 219.220 -36.515 219.480 ;
        RECT -36.455 219.220 -36.195 219.480 ;
        RECT -36.135 219.220 -35.875 219.480 ;
        RECT -35.815 219.220 -35.555 219.480 ;
        RECT -35.495 219.220 -35.235 219.480 ;
        RECT -35.175 219.220 -34.915 219.480 ;
        RECT -34.855 219.220 -34.595 219.480 ;
        RECT -34.535 219.220 -34.275 219.480 ;
        RECT -34.215 219.220 -33.955 219.480 ;
        RECT -33.895 219.220 -33.635 219.480 ;
        RECT -33.575 219.220 -33.315 219.480 ;
        RECT -33.255 219.220 -32.995 219.480 ;
        RECT -32.935 219.220 -32.675 219.480 ;
        RECT -32.615 219.220 -32.355 219.480 ;
        RECT -32.295 219.220 -32.035 219.480 ;
        RECT -31.975 219.220 -31.715 219.480 ;
        RECT -31.655 219.220 -31.395 219.480 ;
        RECT -31.335 219.220 -31.075 219.480 ;
        RECT -31.015 219.220 -30.755 219.480 ;
        RECT -30.695 219.220 -30.435 219.480 ;
        RECT -30.375 219.220 -30.115 219.480 ;
        RECT -30.055 219.220 -29.795 219.480 ;
        RECT -29.735 219.220 -29.475 219.480 ;
        RECT -29.415 219.220 -29.155 219.480 ;
        RECT -29.095 219.220 -28.835 219.480 ;
        RECT -28.775 219.220 -28.515 219.480 ;
        RECT -28.455 219.220 -28.195 219.480 ;
        RECT -28.135 219.220 -27.875 219.480 ;
        RECT -27.815 219.220 -27.555 219.480 ;
        RECT -27.495 219.220 -27.235 219.480 ;
        RECT 99.580 218.510 101.440 220.050 ;
      LAYER met2 ;
        RECT -97.340 223.580 -95.490 223.660 ;
        RECT -97.340 223.500 -72.280 223.580 ;
        RECT -57.720 223.500 -57.050 223.520 ;
        RECT -97.340 223.000 -57.050 223.500 ;
        RECT -97.340 222.970 -72.280 223.000 ;
        RECT -97.340 222.730 -95.490 222.970 ;
        RECT -57.720 219.660 -57.050 223.000 ;
        RECT -49.920 219.660 -27.210 219.680 ;
        RECT 99.540 219.670 101.480 220.220 ;
        RECT -57.720 219.630 -27.210 219.660 ;
        RECT -10.630 219.630 101.480 219.670 ;
        RECT -57.720 219.070 101.480 219.630 ;
        RECT -57.720 219.020 -27.210 219.070 ;
        RECT -10.630 218.470 101.480 219.070 ;
        RECT 99.540 218.340 101.480 218.470 ;
      LAYER via2 ;
        RECT -97.155 222.855 -95.675 223.535 ;
      LAYER met3 ;
        RECT -129.840 223.635 -96.190 224.220 ;
        RECT -129.840 222.755 -95.440 223.635 ;
        RECT -129.840 222.090 -96.190 222.755 ;
    END
  END va
  PIN vb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5000.000000 ;
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER li1 ;
        RECT -96.270 133.080 -96.100 134.700 ;
        RECT -93.690 133.080 -93.520 134.700 ;
        RECT -91.110 133.080 -90.940 134.700 ;
        RECT -88.530 133.080 -88.360 134.700 ;
        RECT -85.950 133.080 -85.780 134.700 ;
        RECT -83.370 133.080 -83.200 134.700 ;
        RECT -80.790 133.080 -80.620 134.700 ;
        RECT -78.210 133.080 -78.040 134.700 ;
        RECT -75.630 133.080 -75.460 134.700 ;
        RECT -73.050 133.080 -72.880 134.700 ;
        RECT -51.050 132.735 -50.880 134.355 ;
        RECT -48.470 132.735 -48.300 134.355 ;
        RECT -45.890 132.735 -45.720 134.355 ;
        RECT -43.310 132.735 -43.140 134.355 ;
        RECT -40.730 132.735 -40.560 134.355 ;
        RECT -38.150 132.735 -37.980 134.355 ;
        RECT -35.570 132.735 -35.400 134.355 ;
        RECT -32.990 132.735 -32.820 134.355 ;
        RECT -30.410 132.735 -30.240 134.355 ;
        RECT -27.830 132.735 -27.660 134.355 ;
        RECT 389.910 132.690 391.580 133.450 ;
        RECT 401.690 132.690 405.410 133.130 ;
        RECT 389.910 132.060 405.410 132.690 ;
        RECT 389.910 131.560 391.580 132.060 ;
        RECT 401.690 131.380 405.410 132.060 ;
      LAYER mcon ;
        RECT -96.270 134.345 -96.100 134.515 ;
        RECT -96.270 133.985 -96.100 134.155 ;
        RECT -96.270 133.625 -96.100 133.795 ;
        RECT -96.270 133.265 -96.100 133.435 ;
        RECT -93.690 134.345 -93.520 134.515 ;
        RECT -93.690 133.985 -93.520 134.155 ;
        RECT -93.690 133.625 -93.520 133.795 ;
        RECT -93.690 133.265 -93.520 133.435 ;
        RECT -91.110 134.345 -90.940 134.515 ;
        RECT -91.110 133.985 -90.940 134.155 ;
        RECT -91.110 133.625 -90.940 133.795 ;
        RECT -91.110 133.265 -90.940 133.435 ;
        RECT -88.530 134.345 -88.360 134.515 ;
        RECT -88.530 133.985 -88.360 134.155 ;
        RECT -88.530 133.625 -88.360 133.795 ;
        RECT -88.530 133.265 -88.360 133.435 ;
        RECT -85.950 134.345 -85.780 134.515 ;
        RECT -85.950 133.985 -85.780 134.155 ;
        RECT -85.950 133.625 -85.780 133.795 ;
        RECT -85.950 133.265 -85.780 133.435 ;
        RECT -83.370 134.345 -83.200 134.515 ;
        RECT -83.370 133.985 -83.200 134.155 ;
        RECT -83.370 133.625 -83.200 133.795 ;
        RECT -83.370 133.265 -83.200 133.435 ;
        RECT -80.790 134.345 -80.620 134.515 ;
        RECT -80.790 133.985 -80.620 134.155 ;
        RECT -80.790 133.625 -80.620 133.795 ;
        RECT -80.790 133.265 -80.620 133.435 ;
        RECT -78.210 134.345 -78.040 134.515 ;
        RECT -78.210 133.985 -78.040 134.155 ;
        RECT -78.210 133.625 -78.040 133.795 ;
        RECT -78.210 133.265 -78.040 133.435 ;
        RECT -75.630 134.345 -75.460 134.515 ;
        RECT -75.630 133.985 -75.460 134.155 ;
        RECT -75.630 133.625 -75.460 133.795 ;
        RECT -75.630 133.265 -75.460 133.435 ;
        RECT -73.050 134.345 -72.880 134.515 ;
        RECT -73.050 133.985 -72.880 134.155 ;
        RECT -73.050 133.625 -72.880 133.795 ;
        RECT -73.050 133.265 -72.880 133.435 ;
        RECT -51.050 134.000 -50.880 134.170 ;
        RECT -51.050 133.640 -50.880 133.810 ;
        RECT -51.050 133.280 -50.880 133.450 ;
        RECT -51.050 132.920 -50.880 133.090 ;
        RECT -48.470 134.000 -48.300 134.170 ;
        RECT -48.470 133.640 -48.300 133.810 ;
        RECT -48.470 133.280 -48.300 133.450 ;
        RECT -48.470 132.920 -48.300 133.090 ;
        RECT -45.890 134.000 -45.720 134.170 ;
        RECT -45.890 133.640 -45.720 133.810 ;
        RECT -45.890 133.280 -45.720 133.450 ;
        RECT -45.890 132.920 -45.720 133.090 ;
        RECT -43.310 134.000 -43.140 134.170 ;
        RECT -43.310 133.640 -43.140 133.810 ;
        RECT -43.310 133.280 -43.140 133.450 ;
        RECT -43.310 132.920 -43.140 133.090 ;
        RECT -40.730 134.000 -40.560 134.170 ;
        RECT -40.730 133.640 -40.560 133.810 ;
        RECT -40.730 133.280 -40.560 133.450 ;
        RECT -40.730 132.920 -40.560 133.090 ;
        RECT -38.150 134.000 -37.980 134.170 ;
        RECT -38.150 133.640 -37.980 133.810 ;
        RECT -38.150 133.280 -37.980 133.450 ;
        RECT -38.150 132.920 -37.980 133.090 ;
        RECT -35.570 134.000 -35.400 134.170 ;
        RECT -35.570 133.640 -35.400 133.810 ;
        RECT -35.570 133.280 -35.400 133.450 ;
        RECT -35.570 132.920 -35.400 133.090 ;
        RECT -32.990 134.000 -32.820 134.170 ;
        RECT -32.990 133.640 -32.820 133.810 ;
        RECT -32.990 133.280 -32.820 133.450 ;
        RECT -32.990 132.920 -32.820 133.090 ;
        RECT -30.410 134.000 -30.240 134.170 ;
        RECT -30.410 133.640 -30.240 133.810 ;
        RECT -30.410 133.280 -30.240 133.450 ;
        RECT -30.410 132.920 -30.240 133.090 ;
        RECT -27.830 134.000 -27.660 134.170 ;
        RECT -27.830 133.640 -27.660 133.810 ;
        RECT -27.830 133.280 -27.660 133.450 ;
        RECT -27.830 132.920 -27.660 133.090 ;
        RECT 389.940 131.700 391.550 133.310 ;
        RECT 402.115 131.815 404.805 132.705 ;
      LAYER met1 ;
        RECT -75.675 135.880 -75.445 138.015 ;
        RECT -96.580 135.200 -72.410 135.880 ;
        RECT -96.305 134.680 -96.095 135.200 ;
        RECT -93.725 134.680 -93.515 135.200 ;
        RECT -91.155 134.680 -90.945 135.200 ;
        RECT -88.595 134.680 -88.385 135.200 ;
        RECT -85.955 134.680 -85.745 135.200 ;
        RECT -96.305 134.345 -96.070 134.680 ;
        RECT -93.725 134.385 -93.490 134.680 ;
        RECT -91.155 134.385 -90.910 134.680 ;
        RECT -96.300 133.100 -96.070 134.345 ;
        RECT -93.720 133.100 -93.490 134.385 ;
        RECT -91.140 133.100 -90.910 134.385 ;
        RECT -88.595 134.365 -88.330 134.680 ;
        RECT -88.560 133.100 -88.330 134.365 ;
        RECT -85.980 134.345 -85.745 134.680 ;
        RECT -83.415 134.680 -83.205 135.200 ;
        RECT -80.775 134.680 -80.565 135.200 ;
        RECT -78.225 134.680 -78.015 135.200 ;
        RECT -75.665 134.680 -75.455 135.200 ;
        RECT -73.045 134.680 -72.835 135.200 ;
        RECT -85.980 133.100 -85.750 134.345 ;
        RECT -83.415 134.315 -83.170 134.680 ;
        RECT -83.400 133.100 -83.170 134.315 ;
        RECT -80.820 134.215 -80.565 134.680 ;
        RECT -80.820 133.100 -80.590 134.215 ;
        RECT -78.240 133.100 -78.010 134.680 ;
        RECT -75.665 134.255 -75.430 134.680 ;
        RECT -75.660 133.100 -75.430 134.255 ;
        RECT -73.080 134.345 -72.835 134.680 ;
        RECT -73.080 133.100 -72.850 134.345 ;
        RECT -51.080 133.010 -50.850 134.335 ;
        RECT -51.085 132.140 -50.845 133.010 ;
        RECT -48.500 132.930 -48.270 134.335 ;
        RECT -45.920 132.950 -45.690 134.335 ;
        RECT -43.340 133.010 -43.110 134.335 ;
        RECT -48.525 132.755 -48.270 132.930 ;
        RECT -48.525 132.140 -48.285 132.755 ;
        RECT -45.925 132.140 -45.685 132.950 ;
        RECT -43.365 132.755 -43.110 133.010 ;
        RECT -40.760 132.970 -40.530 134.335 ;
        RECT -38.180 133.010 -37.950 134.335 ;
        RECT -40.785 132.755 -40.530 132.970 ;
        RECT -43.365 132.140 -43.125 132.755 ;
        RECT -40.785 132.140 -40.545 132.755 ;
        RECT -38.185 132.140 -37.945 133.010 ;
        RECT -35.600 132.990 -35.370 134.335 ;
        RECT -35.605 132.140 -35.365 132.990 ;
        RECT -33.020 132.930 -32.790 134.335 ;
        RECT -30.440 132.970 -30.210 134.335 ;
        RECT -33.025 132.140 -32.785 132.930 ;
        RECT -30.465 132.755 -30.210 132.970 ;
        RECT -27.860 132.950 -27.630 134.335 ;
        RECT 389.880 133.450 391.610 133.510 ;
        RECT -27.860 132.755 -27.575 132.950 ;
        RECT -30.465 132.140 -30.225 132.755 ;
        RECT -27.815 132.140 -27.575 132.755 ;
        RECT -51.450 131.630 -27.220 132.140 ;
        RECT -27.885 129.470 -27.575 131.630 ;
        RECT 389.860 131.560 391.630 133.450 ;
        RECT 389.880 131.500 391.610 131.560 ;
        RECT 401.690 131.380 405.410 133.130 ;
      LAYER via ;
        RECT -96.465 135.250 -72.525 135.830 ;
        RECT -51.305 131.755 -51.045 132.015 ;
        RECT -50.985 131.755 -50.725 132.015 ;
        RECT -50.665 131.755 -50.405 132.015 ;
        RECT -50.345 131.755 -50.085 132.015 ;
        RECT -50.025 131.755 -49.765 132.015 ;
        RECT -49.705 131.755 -49.445 132.015 ;
        RECT -49.385 131.755 -49.125 132.015 ;
        RECT -49.065 131.755 -48.805 132.015 ;
        RECT -48.745 131.755 -48.485 132.015 ;
        RECT -48.425 131.755 -48.165 132.015 ;
        RECT -48.105 131.755 -47.845 132.015 ;
        RECT -47.785 131.755 -47.525 132.015 ;
        RECT -47.465 131.755 -47.205 132.015 ;
        RECT -47.145 131.755 -46.885 132.015 ;
        RECT -46.825 131.755 -46.565 132.015 ;
        RECT -46.505 131.755 -46.245 132.015 ;
        RECT -46.185 131.755 -45.925 132.015 ;
        RECT -45.865 131.755 -45.605 132.015 ;
        RECT -45.545 131.755 -45.285 132.015 ;
        RECT -45.225 131.755 -44.965 132.015 ;
        RECT -44.905 131.755 -44.645 132.015 ;
        RECT -44.585 131.755 -44.325 132.015 ;
        RECT -44.265 131.755 -44.005 132.015 ;
        RECT -43.945 131.755 -43.685 132.015 ;
        RECT -43.625 131.755 -43.365 132.015 ;
        RECT -43.305 131.755 -43.045 132.015 ;
        RECT -42.985 131.755 -42.725 132.015 ;
        RECT -42.665 131.755 -42.405 132.015 ;
        RECT -42.345 131.755 -42.085 132.015 ;
        RECT -42.025 131.755 -41.765 132.015 ;
        RECT -41.705 131.755 -41.445 132.015 ;
        RECT -41.385 131.755 -41.125 132.015 ;
        RECT -41.065 131.755 -40.805 132.015 ;
        RECT -40.745 131.755 -40.485 132.015 ;
        RECT -40.425 131.755 -40.165 132.015 ;
        RECT -40.105 131.755 -39.845 132.015 ;
        RECT -39.785 131.755 -39.525 132.015 ;
        RECT -39.465 131.755 -39.205 132.015 ;
        RECT -39.145 131.755 -38.885 132.015 ;
        RECT -38.825 131.755 -38.565 132.015 ;
        RECT -38.505 131.755 -38.245 132.015 ;
        RECT -38.185 131.755 -37.925 132.015 ;
        RECT -37.865 131.755 -37.605 132.015 ;
        RECT -37.545 131.755 -37.285 132.015 ;
        RECT -37.225 131.755 -36.965 132.015 ;
        RECT -36.905 131.755 -36.645 132.015 ;
        RECT -36.585 131.755 -36.325 132.015 ;
        RECT -36.265 131.755 -36.005 132.015 ;
        RECT -35.945 131.755 -35.685 132.015 ;
        RECT -35.625 131.755 -35.365 132.015 ;
        RECT -35.305 131.755 -35.045 132.015 ;
        RECT -34.985 131.755 -34.725 132.015 ;
        RECT -34.665 131.755 -34.405 132.015 ;
        RECT -34.345 131.755 -34.085 132.015 ;
        RECT -34.025 131.755 -33.765 132.015 ;
        RECT -33.705 131.755 -33.445 132.015 ;
        RECT -33.385 131.755 -33.125 132.015 ;
        RECT -33.065 131.755 -32.805 132.015 ;
        RECT -32.745 131.755 -32.485 132.015 ;
        RECT -32.425 131.755 -32.165 132.015 ;
        RECT -32.105 131.755 -31.845 132.015 ;
        RECT -31.785 131.755 -31.525 132.015 ;
        RECT -31.465 131.755 -31.205 132.015 ;
        RECT -31.145 131.755 -30.885 132.015 ;
        RECT -30.825 131.755 -30.565 132.015 ;
        RECT -30.505 131.755 -30.245 132.015 ;
        RECT -30.185 131.755 -29.925 132.015 ;
        RECT -29.865 131.755 -29.605 132.015 ;
        RECT -29.545 131.755 -29.285 132.015 ;
        RECT -29.225 131.755 -28.965 132.015 ;
        RECT -28.905 131.755 -28.645 132.015 ;
        RECT -28.585 131.755 -28.325 132.015 ;
        RECT -28.265 131.755 -28.005 132.015 ;
        RECT -27.945 131.755 -27.685 132.015 ;
        RECT -27.625 131.755 -27.365 132.015 ;
        RECT 389.975 131.575 391.515 133.435 ;
      LAYER met2 ;
        RECT -97.670 135.930 -93.970 136.100 ;
        RECT -97.670 135.830 -72.460 135.930 ;
        RECT -97.670 135.150 -60.480 135.830 ;
        RECT -97.670 135.060 -93.970 135.150 ;
        RECT -61.480 132.250 -60.480 135.150 ;
        RECT -10.080 133.150 -4.840 133.160 ;
        RECT -10.080 133.090 195.640 133.150 ;
        RECT 389.910 133.090 391.580 133.500 ;
        RECT -61.480 132.190 -47.880 132.250 ;
        RECT -10.080 132.230 391.580 133.090 ;
        RECT -28.330 132.190 391.580 132.230 ;
        RECT -61.480 132.170 391.580 132.190 ;
        RECT -61.480 132.020 195.640 132.170 ;
        RECT -61.480 131.710 -4.840 132.020 ;
        RECT -61.480 131.670 -4.880 131.710 ;
        RECT -61.480 131.580 -27.270 131.670 ;
        RECT -61.480 131.570 -47.880 131.580 ;
        RECT 389.910 131.510 391.580 132.170 ;
      LAYER via2 ;
        RECT -97.560 135.240 -94.080 135.920 ;
      LAYER met3 ;
        RECT -129.910 136.075 -96.260 136.940 ;
        RECT -129.910 135.085 -93.920 136.075 ;
        RECT -129.910 134.810 -96.260 135.085 ;
    END
  END vb
  PIN vcap
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 659.750000 ;
    PORT
      LAYER li1 ;
        RECT 198.520 215.550 200.240 219.390 ;
        RECT 112.630 214.790 112.800 215.340 ;
        RECT 123.210 214.820 123.380 215.340 ;
        RECT 133.790 214.900 133.960 215.340 ;
        RECT 112.610 192.980 112.840 214.790 ;
        RECT 123.210 193.010 123.440 214.820 ;
        RECT 133.750 193.090 133.980 214.900 ;
        RECT 145.240 214.870 145.410 215.420 ;
        RECT 155.820 214.900 155.990 215.420 ;
        RECT 166.400 214.980 166.570 215.420 ;
        RECT 112.630 192.420 112.800 192.980 ;
        RECT 112.530 191.370 112.940 192.420 ;
        RECT 123.210 192.280 123.380 193.010 ;
        RECT 133.790 192.650 133.960 193.090 ;
        RECT 145.220 193.060 145.450 214.870 ;
        RECT 155.820 193.090 156.050 214.900 ;
        RECT 166.360 193.170 166.590 214.980 ;
        RECT 177.790 214.900 177.960 215.450 ;
        RECT 188.370 214.930 188.540 215.450 ;
        RECT 123.160 191.370 123.570 192.280 ;
        RECT 133.520 191.370 134.180 192.650 ;
        RECT 145.240 192.500 145.410 193.060 ;
        RECT 145.140 191.450 145.550 192.500 ;
        RECT 155.820 192.360 155.990 193.090 ;
        RECT 166.400 192.470 166.570 193.170 ;
        RECT 177.770 193.090 178.000 214.900 ;
        RECT 188.370 193.120 188.600 214.930 ;
        RECT 198.790 213.650 199.610 215.550 ;
        RECT 198.910 193.200 199.140 213.650 ;
        RECT 177.790 192.530 177.960 193.090 ;
        RECT 155.770 191.450 156.180 192.360 ;
        RECT 166.250 191.450 166.910 192.470 ;
        RECT 177.690 191.480 178.100 192.530 ;
        RECT 188.370 192.390 188.540 193.120 ;
        RECT 198.950 192.500 199.120 193.200 ;
        RECT 198.830 192.480 199.240 192.500 ;
        RECT 188.320 191.480 188.730 192.390 ;
        RECT 198.830 191.480 199.470 192.480 ;
        RECT 112.530 190.920 134.780 191.370 ;
        RECT 145.140 191.000 167.390 191.450 ;
        RECT 177.690 191.030 199.940 191.480 ;
        RECT 177.750 191.000 199.940 191.030 ;
        RECT 145.200 190.970 167.390 191.000 ;
        RECT 112.590 190.890 134.780 190.920 ;
        RECT 123.160 190.780 123.570 190.890 ;
        RECT 112.630 185.710 112.800 186.260 ;
        RECT 123.210 185.740 123.380 186.260 ;
        RECT 112.610 163.900 112.840 185.710 ;
        RECT 123.210 163.930 123.440 185.740 ;
        RECT 133.520 185.610 134.180 190.890 ;
        RECT 155.770 190.860 156.180 190.970 ;
        RECT 145.240 185.790 145.410 186.340 ;
        RECT 155.820 185.820 155.990 186.340 ;
        RECT 133.750 164.010 133.980 185.610 ;
        RECT 112.630 163.340 112.800 163.900 ;
        RECT 112.530 162.290 112.940 163.340 ;
        RECT 123.210 163.200 123.380 163.930 ;
        RECT 133.790 163.310 133.960 164.010 ;
        RECT 145.220 163.980 145.450 185.790 ;
        RECT 155.820 164.010 156.050 185.820 ;
        RECT 166.250 185.430 166.910 190.970 ;
        RECT 188.320 190.890 188.730 191.000 ;
        RECT 177.790 185.820 177.960 186.370 ;
        RECT 188.370 185.850 188.540 186.370 ;
        RECT 166.360 164.090 166.590 185.430 ;
        RECT 145.240 163.420 145.410 163.980 ;
        RECT 133.670 163.240 134.080 163.310 ;
        RECT 123.160 162.290 123.570 163.200 ;
        RECT 133.670 162.290 134.400 163.240 ;
        RECT 145.140 162.370 145.550 163.420 ;
        RECT 155.820 163.280 155.990 164.010 ;
        RECT 166.400 163.390 166.570 164.090 ;
        RECT 177.770 164.010 178.000 185.820 ;
        RECT 188.370 164.040 188.600 185.850 ;
        RECT 198.840 185.560 199.470 191.000 ;
        RECT 198.910 164.120 199.140 185.560 ;
        RECT 177.790 163.450 177.960 164.010 ;
        RECT 155.770 162.370 156.180 163.280 ;
        RECT 166.280 163.200 166.690 163.390 ;
        RECT 166.140 162.370 166.800 163.200 ;
        RECT 177.690 162.400 178.100 163.450 ;
        RECT 188.370 163.310 188.540 164.040 ;
        RECT 198.950 163.580 199.120 164.120 ;
        RECT 188.320 162.400 188.730 163.310 ;
        RECT 198.770 162.400 199.400 163.580 ;
        RECT 112.530 161.840 134.780 162.290 ;
        RECT 145.140 161.920 167.390 162.370 ;
        RECT 177.690 161.950 199.940 162.400 ;
        RECT 177.750 161.920 199.940 161.950 ;
        RECT 145.200 161.890 167.390 161.920 ;
        RECT 112.590 161.810 134.780 161.840 ;
        RECT 123.160 161.700 123.570 161.810 ;
        RECT 112.630 156.540 112.800 157.090 ;
        RECT 123.210 156.570 123.380 157.090 ;
        RECT 112.610 134.730 112.840 156.540 ;
        RECT 123.210 134.760 123.440 156.570 ;
        RECT 133.740 156.200 134.400 161.810 ;
        RECT 155.770 161.780 156.180 161.890 ;
        RECT 145.240 156.620 145.410 157.170 ;
        RECT 155.820 156.650 155.990 157.170 ;
        RECT 133.750 134.840 133.980 156.200 ;
        RECT 112.630 134.170 112.800 134.730 ;
        RECT 112.530 133.120 112.940 134.170 ;
        RECT 123.210 134.030 123.380 134.760 ;
        RECT 133.790 134.390 133.960 134.840 ;
        RECT 145.220 134.810 145.450 156.620 ;
        RECT 155.820 134.840 156.050 156.650 ;
        RECT 166.140 156.160 166.800 161.890 ;
        RECT 188.320 161.810 188.730 161.920 ;
        RECT 177.790 156.650 177.960 157.200 ;
        RECT 188.370 156.680 188.540 157.200 ;
        RECT 166.360 134.920 166.590 156.160 ;
        RECT 133.700 134.140 134.360 134.390 ;
        RECT 145.240 134.250 145.410 134.810 ;
        RECT 123.160 133.120 123.570 134.030 ;
        RECT 133.670 133.120 134.360 134.140 ;
        RECT 145.140 133.200 145.550 134.250 ;
        RECT 155.820 134.110 155.990 134.840 ;
        RECT 166.400 134.220 166.570 134.920 ;
        RECT 177.770 134.840 178.000 156.650 ;
        RECT 188.370 134.870 188.600 156.680 ;
        RECT 198.770 156.660 199.400 161.920 ;
        RECT 198.910 134.950 199.140 156.660 ;
        RECT 177.790 134.280 177.960 134.840 ;
        RECT 166.280 134.120 166.690 134.220 ;
        RECT 155.770 133.200 156.180 134.110 ;
        RECT 166.280 133.200 166.920 134.120 ;
        RECT 177.690 133.230 178.100 134.280 ;
        RECT 188.370 134.140 188.540 134.870 ;
        RECT 198.950 134.250 199.120 134.950 ;
        RECT 188.320 133.230 188.730 134.140 ;
        RECT 198.830 133.770 199.240 134.250 ;
        RECT 198.770 133.230 199.400 133.770 ;
        RECT 112.530 132.670 134.780 133.120 ;
        RECT 145.140 132.750 167.390 133.200 ;
        RECT 177.690 132.780 199.940 133.230 ;
        RECT 177.750 132.750 199.940 132.780 ;
        RECT 145.200 132.720 167.390 132.750 ;
        RECT 112.590 132.640 134.780 132.670 ;
        RECT 123.160 132.530 123.570 132.640 ;
        RECT 112.630 127.360 112.800 127.910 ;
        RECT 123.210 127.390 123.380 127.910 ;
        RECT 112.610 105.550 112.840 127.360 ;
        RECT 123.210 105.580 123.440 127.390 ;
        RECT 133.700 127.350 134.360 132.640 ;
        RECT 155.770 132.610 156.180 132.720 ;
        RECT 145.240 127.440 145.410 127.990 ;
        RECT 155.820 127.470 155.990 127.990 ;
        RECT 133.750 105.660 133.980 127.350 ;
        RECT 112.630 104.990 112.800 105.550 ;
        RECT 112.530 103.940 112.940 104.990 ;
        RECT 123.210 104.850 123.380 105.580 ;
        RECT 133.790 105.020 133.960 105.660 ;
        RECT 145.220 105.630 145.450 127.440 ;
        RECT 155.820 105.660 156.050 127.470 ;
        RECT 166.290 127.200 166.920 132.720 ;
        RECT 188.320 132.640 188.730 132.750 ;
        RECT 177.790 127.470 177.960 128.020 ;
        RECT 188.370 127.500 188.540 128.020 ;
        RECT 166.360 105.740 166.590 127.200 ;
        RECT 145.240 105.070 145.410 105.630 ;
        RECT 123.160 103.940 123.570 104.850 ;
        RECT 133.440 103.940 134.100 105.020 ;
        RECT 145.140 104.020 145.550 105.070 ;
        RECT 155.820 104.930 155.990 105.660 ;
        RECT 166.400 105.040 166.570 105.740 ;
        RECT 177.770 105.660 178.000 127.470 ;
        RECT 188.370 105.690 188.600 127.500 ;
        RECT 198.770 126.850 199.400 132.750 ;
        RECT 397.410 129.180 397.750 129.250 ;
        RECT 376.270 129.090 376.610 129.140 ;
        RECT 386.790 129.090 387.130 129.170 ;
        RECT 397.310 129.090 410.400 129.180 ;
        RECT 376.270 129.080 410.400 129.090 ;
        RECT 419.100 129.080 419.440 129.160 ;
        RECT 429.720 129.080 430.060 129.240 ;
        RECT 376.270 129.040 430.060 129.080 ;
        RECT 375.580 128.810 430.060 129.040 ;
        RECT 375.580 128.640 430.100 128.810 ;
        RECT 375.580 128.590 397.030 128.640 ;
        RECT 397.310 128.630 430.100 128.640 ;
        RECT 376.270 127.190 376.610 128.590 ;
        RECT 386.790 127.520 387.130 128.590 ;
        RECT 397.310 128.580 429.340 128.630 ;
        RECT 397.310 128.410 410.400 128.580 ;
        RECT 386.790 127.260 387.160 127.520 ;
        RECT 198.910 105.770 199.140 126.850 ;
        RECT 376.270 126.160 376.510 127.190 ;
        RECT 376.270 122.310 376.500 126.160 ;
        RECT 376.270 120.690 376.510 122.310 ;
        RECT 376.270 116.840 376.500 120.690 ;
        RECT 376.270 115.220 376.510 116.840 ;
        RECT 376.270 111.370 376.500 115.220 ;
        RECT 376.270 109.750 376.510 111.370 ;
        RECT 376.270 105.900 376.500 109.750 ;
        RECT 177.790 105.100 177.960 105.660 ;
        RECT 155.770 104.020 156.180 104.930 ;
        RECT 166.280 104.790 166.690 105.040 ;
        RECT 166.220 104.020 166.850 104.790 ;
        RECT 177.690 104.050 178.100 105.100 ;
        RECT 188.370 104.960 188.540 105.690 ;
        RECT 198.950 105.070 199.120 105.770 ;
        RECT 376.270 105.530 376.510 105.900 ;
        RECT 386.870 105.530 387.100 127.260 ;
        RECT 397.370 127.240 397.790 128.410 ;
        RECT 397.470 105.670 397.700 127.240 ;
        RECT 408.580 127.180 408.920 128.410 ;
        RECT 419.100 127.510 419.440 128.580 ;
        RECT 419.100 127.250 419.470 127.510 ;
        RECT 408.580 126.150 408.820 127.180 ;
        RECT 408.580 122.300 408.810 126.150 ;
        RECT 408.580 120.680 408.820 122.300 ;
        RECT 408.580 116.830 408.810 120.680 ;
        RECT 408.580 115.210 408.820 116.830 ;
        RECT 408.580 111.360 408.810 115.210 ;
        RECT 408.580 109.740 408.820 111.360 ;
        RECT 408.580 105.890 408.810 109.740 ;
        RECT 188.320 104.050 188.730 104.960 ;
        RECT 198.830 104.790 199.240 105.070 ;
        RECT 198.770 104.050 199.400 104.790 ;
        RECT 376.340 104.280 376.510 105.530 ;
        RECT 386.920 104.280 387.090 105.530 ;
        RECT 397.500 104.280 397.670 105.670 ;
        RECT 408.580 105.520 408.820 105.890 ;
        RECT 419.180 105.520 419.410 127.250 ;
        RECT 429.680 127.230 430.100 128.630 ;
        RECT 429.780 105.660 430.010 127.230 ;
        RECT 408.650 104.270 408.820 105.520 ;
        RECT 419.230 104.270 419.400 105.520 ;
        RECT 429.810 104.270 429.980 105.660 ;
        RECT 112.530 103.490 134.780 103.940 ;
        RECT 145.140 103.570 167.390 104.020 ;
        RECT 177.690 103.600 199.940 104.050 ;
        RECT 177.750 103.570 199.940 103.600 ;
        RECT 145.200 103.540 167.390 103.570 ;
        RECT 112.590 103.460 134.780 103.490 ;
        RECT 123.160 103.350 123.570 103.460 ;
        RECT 112.630 98.040 112.800 98.590 ;
        RECT 123.210 98.070 123.380 98.590 ;
        RECT 112.610 76.230 112.840 98.040 ;
        RECT 123.210 76.260 123.440 98.070 ;
        RECT 133.440 97.980 134.100 103.460 ;
        RECT 155.770 103.430 156.180 103.540 ;
        RECT 145.240 98.120 145.410 98.670 ;
        RECT 155.820 98.150 155.990 98.670 ;
        RECT 133.750 76.340 133.980 97.980 ;
        RECT 112.630 75.670 112.800 76.230 ;
        RECT 112.530 74.620 112.940 75.670 ;
        RECT 123.210 75.530 123.380 76.260 ;
        RECT 133.790 75.800 133.960 76.340 ;
        RECT 145.220 76.310 145.450 98.120 ;
        RECT 155.820 76.340 156.050 98.150 ;
        RECT 166.220 97.870 166.850 103.540 ;
        RECT 188.320 103.460 188.730 103.570 ;
        RECT 177.790 98.150 177.960 98.700 ;
        RECT 188.370 98.180 188.540 98.700 ;
        RECT 166.360 76.420 166.590 97.870 ;
        RECT 133.740 75.640 134.400 75.800 ;
        RECT 145.240 75.750 145.410 76.310 ;
        RECT 123.160 74.620 123.570 75.530 ;
        RECT 133.670 74.620 134.400 75.640 ;
        RECT 145.140 74.700 145.550 75.750 ;
        RECT 155.820 75.610 155.990 76.340 ;
        RECT 166.400 75.720 166.570 76.420 ;
        RECT 177.770 76.340 178.000 98.150 ;
        RECT 188.370 76.370 188.600 98.180 ;
        RECT 198.770 97.870 199.400 103.570 ;
        RECT 376.300 99.900 376.640 99.950 ;
        RECT 386.820 99.900 387.160 99.980 ;
        RECT 397.440 99.900 397.780 100.060 ;
        RECT 408.620 99.960 408.960 100.010 ;
        RECT 419.140 99.960 419.480 100.040 ;
        RECT 429.760 99.960 430.100 100.120 ;
        RECT 408.620 99.910 430.100 99.960 ;
        RECT 376.300 99.850 397.780 99.900 ;
        RECT 375.610 99.630 397.780 99.850 ;
        RECT 407.930 99.690 430.100 99.910 ;
        RECT 375.610 99.450 397.820 99.630 ;
        RECT 407.930 99.510 430.140 99.690 ;
        RECT 407.930 99.460 429.380 99.510 ;
        RECT 375.610 99.400 397.060 99.450 ;
        RECT 376.300 98.000 376.640 99.400 ;
        RECT 386.820 98.330 387.160 99.400 ;
        RECT 386.820 98.070 387.190 98.330 ;
        RECT 198.910 76.450 199.140 97.870 ;
        RECT 376.300 96.970 376.540 98.000 ;
        RECT 376.300 93.120 376.530 96.970 ;
        RECT 376.300 91.500 376.540 93.120 ;
        RECT 376.300 87.650 376.530 91.500 ;
        RECT 376.300 86.030 376.540 87.650 ;
        RECT 376.300 82.180 376.530 86.030 ;
        RECT 376.300 80.560 376.540 82.180 ;
        RECT 376.300 76.710 376.530 80.560 ;
        RECT 177.790 75.780 177.960 76.340 ;
        RECT 155.770 74.700 156.180 75.610 ;
        RECT 166.280 75.190 166.690 75.720 ;
        RECT 166.220 74.700 166.850 75.190 ;
        RECT 177.690 74.730 178.100 75.780 ;
        RECT 188.370 75.640 188.540 76.370 ;
        RECT 198.950 75.750 199.120 76.450 ;
        RECT 376.300 76.340 376.540 76.710 ;
        RECT 386.900 76.340 387.130 98.070 ;
        RECT 397.400 98.050 397.820 99.450 ;
        RECT 408.620 98.060 408.960 99.460 ;
        RECT 419.140 98.390 419.480 99.460 ;
        RECT 419.140 98.130 419.510 98.390 ;
        RECT 397.500 76.480 397.730 98.050 ;
        RECT 408.620 97.030 408.860 98.060 ;
        RECT 408.620 93.180 408.850 97.030 ;
        RECT 408.620 91.560 408.860 93.180 ;
        RECT 408.620 87.710 408.850 91.560 ;
        RECT 408.620 86.090 408.860 87.710 ;
        RECT 408.620 82.240 408.850 86.090 ;
        RECT 408.620 80.620 408.860 82.240 ;
        RECT 408.620 76.770 408.850 80.620 ;
        RECT 188.320 74.730 188.730 75.640 ;
        RECT 198.830 75.400 199.240 75.750 ;
        RECT 198.830 74.730 199.470 75.400 ;
        RECT 376.370 75.090 376.540 76.340 ;
        RECT 386.950 75.090 387.120 76.340 ;
        RECT 397.530 75.090 397.700 76.480 ;
        RECT 408.620 76.400 408.860 76.770 ;
        RECT 419.220 76.400 419.450 98.130 ;
        RECT 429.720 98.110 430.140 99.510 ;
        RECT 429.820 76.540 430.050 98.110 ;
        RECT 408.690 75.150 408.860 76.400 ;
        RECT 419.270 75.150 419.440 76.400 ;
        RECT 429.850 75.150 430.020 76.540 ;
        RECT 112.530 74.170 134.780 74.620 ;
        RECT 145.140 74.250 167.390 74.700 ;
        RECT 177.690 74.280 199.940 74.730 ;
        RECT 177.750 74.250 199.940 74.280 ;
        RECT 145.200 74.220 167.390 74.250 ;
        RECT 112.590 74.140 134.780 74.170 ;
        RECT 123.160 74.030 123.570 74.140 ;
        RECT 112.680 68.760 112.850 69.310 ;
        RECT 123.260 68.790 123.430 69.310 ;
        RECT 112.660 46.950 112.890 68.760 ;
        RECT 123.260 46.980 123.490 68.790 ;
        RECT 133.740 68.760 134.400 74.140 ;
        RECT 155.770 74.110 156.180 74.220 ;
        RECT 145.290 68.840 145.460 69.390 ;
        RECT 155.870 68.870 156.040 69.390 ;
        RECT 133.800 47.060 134.030 68.760 ;
        RECT 112.680 46.390 112.850 46.950 ;
        RECT 112.580 45.340 112.990 46.390 ;
        RECT 123.260 46.250 123.430 46.980 ;
        RECT 133.840 46.360 134.010 47.060 ;
        RECT 145.270 47.030 145.500 68.840 ;
        RECT 155.870 47.060 156.100 68.870 ;
        RECT 166.220 68.270 166.850 74.220 ;
        RECT 188.320 74.140 188.730 74.250 ;
        RECT 177.840 68.870 178.010 69.420 ;
        RECT 188.420 68.900 188.590 69.420 ;
        RECT 166.410 47.140 166.640 68.270 ;
        RECT 145.290 46.470 145.460 47.030 ;
        RECT 123.210 45.340 123.620 46.250 ;
        RECT 133.720 46.090 134.130 46.360 ;
        RECT 133.550 45.340 134.210 46.090 ;
        RECT 145.190 45.420 145.600 46.470 ;
        RECT 155.870 46.330 156.040 47.060 ;
        RECT 166.450 46.440 166.620 47.140 ;
        RECT 177.820 47.060 178.050 68.870 ;
        RECT 188.420 47.090 188.650 68.900 ;
        RECT 198.840 68.480 199.470 74.250 ;
        RECT 376.300 70.610 376.640 70.660 ;
        RECT 386.820 70.610 387.160 70.690 ;
        RECT 397.440 70.610 397.780 70.770 ;
        RECT 376.300 70.560 397.780 70.610 ;
        RECT 375.610 70.340 397.780 70.560 ;
        RECT 408.640 70.600 408.980 70.650 ;
        RECT 419.160 70.600 419.500 70.680 ;
        RECT 429.780 70.600 430.120 70.760 ;
        RECT 408.640 70.550 430.120 70.600 ;
        RECT 375.610 70.160 397.820 70.340 ;
        RECT 375.610 70.110 397.060 70.160 ;
        RECT 376.300 68.710 376.640 70.110 ;
        RECT 386.820 69.040 387.160 70.110 ;
        RECT 386.820 68.780 387.190 69.040 ;
        RECT 198.960 47.170 199.190 68.480 ;
        RECT 376.300 67.680 376.540 68.710 ;
        RECT 376.300 63.830 376.530 67.680 ;
        RECT 376.300 62.210 376.540 63.830 ;
        RECT 376.300 58.360 376.530 62.210 ;
        RECT 376.300 56.740 376.540 58.360 ;
        RECT 376.300 52.890 376.530 56.740 ;
        RECT 376.300 51.270 376.540 52.890 ;
        RECT 376.300 47.420 376.530 51.270 ;
        RECT 177.840 46.500 178.010 47.060 ;
        RECT 155.820 45.420 156.230 46.330 ;
        RECT 166.330 46.010 166.740 46.440 ;
        RECT 166.290 45.420 166.920 46.010 ;
        RECT 177.740 45.450 178.150 46.500 ;
        RECT 188.420 46.360 188.590 47.090 ;
        RECT 199.000 46.470 199.170 47.170 ;
        RECT 376.300 47.050 376.540 47.420 ;
        RECT 386.900 47.050 387.130 68.780 ;
        RECT 397.400 68.760 397.820 70.160 ;
        RECT 407.950 70.330 430.120 70.550 ;
        RECT 407.950 70.150 430.160 70.330 ;
        RECT 407.950 70.100 429.400 70.150 ;
        RECT 397.500 47.190 397.730 68.760 ;
        RECT 408.640 68.700 408.980 70.100 ;
        RECT 419.160 69.030 419.500 70.100 ;
        RECT 419.160 68.770 419.530 69.030 ;
        RECT 408.640 67.670 408.880 68.700 ;
        RECT 408.640 63.820 408.870 67.670 ;
        RECT 408.640 62.200 408.880 63.820 ;
        RECT 408.640 58.350 408.870 62.200 ;
        RECT 408.640 56.730 408.880 58.350 ;
        RECT 408.640 52.880 408.870 56.730 ;
        RECT 408.640 51.260 408.880 52.880 ;
        RECT 408.640 47.410 408.870 51.260 ;
        RECT 188.370 45.450 188.780 46.360 ;
        RECT 198.880 46.290 199.290 46.470 ;
        RECT 198.880 45.450 199.540 46.290 ;
        RECT 376.370 45.800 376.540 47.050 ;
        RECT 386.950 45.800 387.120 47.050 ;
        RECT 397.530 45.800 397.700 47.190 ;
        RECT 408.640 47.040 408.880 47.410 ;
        RECT 419.240 47.040 419.470 68.770 ;
        RECT 429.740 68.750 430.160 70.150 ;
        RECT 429.840 47.180 430.070 68.750 ;
        RECT 408.710 45.790 408.880 47.040 ;
        RECT 419.290 45.790 419.460 47.040 ;
        RECT 429.870 45.790 430.040 47.180 ;
        RECT 112.580 44.890 134.830 45.340 ;
        RECT 145.190 44.970 167.440 45.420 ;
        RECT 177.740 45.000 199.990 45.450 ;
        RECT 177.800 44.970 199.990 45.000 ;
        RECT 145.250 44.940 167.440 44.970 ;
        RECT 112.640 44.860 134.830 44.890 ;
        RECT 123.210 44.750 123.620 44.860 ;
        RECT 112.770 39.220 112.940 39.770 ;
        RECT 123.350 39.250 123.520 39.770 ;
        RECT 112.750 17.410 112.980 39.220 ;
        RECT 123.350 17.440 123.580 39.250 ;
        RECT 133.550 39.050 134.210 44.860 ;
        RECT 155.820 44.830 156.230 44.940 ;
        RECT 145.380 39.300 145.550 39.850 ;
        RECT 155.960 39.330 156.130 39.850 ;
        RECT 133.890 17.520 134.120 39.050 ;
        RECT 112.770 16.850 112.940 17.410 ;
        RECT 112.670 15.800 113.080 16.850 ;
        RECT 123.350 16.710 123.520 17.440 ;
        RECT 133.930 16.820 134.100 17.520 ;
        RECT 145.360 17.490 145.590 39.300 ;
        RECT 155.960 17.520 156.190 39.330 ;
        RECT 166.290 39.090 166.920 44.940 ;
        RECT 188.370 44.860 188.780 44.970 ;
        RECT 177.930 39.330 178.100 39.880 ;
        RECT 188.510 39.360 188.680 39.880 ;
        RECT 198.910 39.370 199.540 44.970 ;
        RECT 376.300 41.320 376.640 41.370 ;
        RECT 386.820 41.320 387.160 41.400 ;
        RECT 397.440 41.320 397.780 41.480 ;
        RECT 376.300 41.270 397.780 41.320 ;
        RECT 375.610 41.050 397.780 41.270 ;
        RECT 408.660 41.310 409.000 41.360 ;
        RECT 419.180 41.310 419.520 41.390 ;
        RECT 429.800 41.310 430.140 41.470 ;
        RECT 408.660 41.260 430.140 41.310 ;
        RECT 375.610 40.870 397.820 41.050 ;
        RECT 375.610 40.820 397.060 40.870 ;
        RECT 376.300 39.420 376.640 40.820 ;
        RECT 386.820 39.750 387.160 40.820 ;
        RECT 386.820 39.490 387.190 39.750 ;
        RECT 166.500 17.600 166.730 39.090 ;
        RECT 145.380 16.930 145.550 17.490 ;
        RECT 123.300 15.800 123.710 16.710 ;
        RECT 133.810 15.820 134.220 16.820 ;
        RECT 145.280 15.880 145.690 16.930 ;
        RECT 155.960 16.790 156.130 17.520 ;
        RECT 166.540 16.900 166.710 17.600 ;
        RECT 177.910 17.520 178.140 39.330 ;
        RECT 188.510 17.550 188.740 39.360 ;
        RECT 199.050 17.630 199.280 39.370 ;
        RECT 376.300 38.390 376.540 39.420 ;
        RECT 376.300 34.540 376.530 38.390 ;
        RECT 376.300 32.920 376.540 34.540 ;
        RECT 376.300 29.070 376.530 32.920 ;
        RECT 376.300 27.450 376.540 29.070 ;
        RECT 376.300 23.600 376.530 27.450 ;
        RECT 376.300 21.980 376.540 23.600 ;
        RECT 376.300 18.130 376.530 21.980 ;
        RECT 376.300 17.760 376.540 18.130 ;
        RECT 386.900 17.760 387.130 39.490 ;
        RECT 397.400 39.470 397.820 40.870 ;
        RECT 407.970 41.040 430.140 41.260 ;
        RECT 407.970 40.860 430.180 41.040 ;
        RECT 407.970 40.810 429.420 40.860 ;
        RECT 397.500 17.900 397.730 39.470 ;
        RECT 408.660 39.410 409.000 40.810 ;
        RECT 419.180 39.740 419.520 40.810 ;
        RECT 419.180 39.480 419.550 39.740 ;
        RECT 408.660 38.380 408.900 39.410 ;
        RECT 408.660 34.530 408.890 38.380 ;
        RECT 408.660 32.910 408.900 34.530 ;
        RECT 408.660 29.060 408.890 32.910 ;
        RECT 408.660 27.440 408.900 29.060 ;
        RECT 408.660 23.590 408.890 27.440 ;
        RECT 408.660 21.970 408.900 23.590 ;
        RECT 408.660 18.120 408.890 21.970 ;
        RECT 177.930 16.960 178.100 17.520 ;
        RECT 155.910 15.880 156.320 16.790 ;
        RECT 166.420 16.140 166.830 16.900 ;
        RECT 177.830 16.140 178.240 16.960 ;
        RECT 188.510 16.820 188.680 17.550 ;
        RECT 199.090 16.930 199.260 17.630 ;
        RECT 165.130 15.910 180.110 16.140 ;
        RECT 188.460 15.910 188.870 16.820 ;
        RECT 198.970 15.910 199.380 16.930 ;
        RECT 376.370 16.510 376.540 17.760 ;
        RECT 386.950 16.510 387.120 17.760 ;
        RECT 397.530 16.510 397.700 17.900 ;
        RECT 408.660 17.750 408.900 18.120 ;
        RECT 419.260 17.750 419.490 39.480 ;
        RECT 429.760 39.460 430.180 40.860 ;
        RECT 429.860 17.890 430.090 39.460 ;
        RECT 408.730 16.500 408.900 17.750 ;
        RECT 419.310 16.500 419.480 17.750 ;
        RECT 429.890 16.500 430.060 17.890 ;
        RECT 165.130 15.880 200.080 15.910 ;
        RECT 145.280 15.820 200.080 15.880 ;
        RECT 132.510 15.800 200.080 15.820 ;
        RECT 112.670 15.430 200.080 15.800 ;
        RECT 112.670 15.400 180.110 15.430 ;
        RECT -95.840 13.750 -95.670 15.370 ;
        RECT -93.260 13.750 -93.090 15.370 ;
        RECT -90.680 13.750 -90.510 15.370 ;
        RECT -88.100 13.750 -87.930 15.370 ;
        RECT -85.520 13.750 -85.350 15.370 ;
        RECT -82.940 13.750 -82.770 15.370 ;
        RECT -80.360 13.750 -80.190 15.370 ;
        RECT -77.780 13.750 -77.610 15.370 ;
        RECT -75.200 13.750 -75.030 15.370 ;
        RECT -72.620 13.750 -72.450 15.370 ;
        RECT 112.670 15.350 147.620 15.400 ;
        RECT 112.730 15.320 147.620 15.350 ;
        RECT 123.300 15.210 123.710 15.320 ;
        RECT -50.930 13.295 -50.760 14.915 ;
        RECT -48.350 13.295 -48.180 14.915 ;
        RECT -45.770 13.295 -45.600 14.915 ;
        RECT -43.190 13.295 -43.020 14.915 ;
        RECT -40.610 13.295 -40.440 14.915 ;
        RECT -38.030 13.295 -37.860 14.915 ;
        RECT -35.450 13.295 -35.280 14.915 ;
        RECT -32.870 13.295 -32.700 14.915 ;
        RECT -30.290 13.295 -30.120 14.915 ;
        RECT -27.710 13.295 -27.540 14.915 ;
        RECT 132.510 14.800 147.620 15.320 ;
        RECT 155.910 15.290 156.320 15.400 ;
        RECT 165.130 14.850 180.110 15.400 ;
        RECT 188.460 15.320 188.870 15.430 ;
      LAYER mcon ;
        RECT 112.630 214.985 112.800 215.155 ;
        RECT 112.630 214.625 112.800 214.795 ;
        RECT 123.210 214.985 123.380 215.155 ;
        RECT 133.790 214.985 133.960 215.155 ;
        RECT 145.240 215.065 145.410 215.235 ;
        RECT 112.630 214.265 112.800 214.435 ;
        RECT 112.630 213.905 112.800 214.075 ;
        RECT 112.630 209.515 112.800 209.685 ;
        RECT 112.630 209.155 112.800 209.325 ;
        RECT 112.630 208.795 112.800 208.965 ;
        RECT 112.630 208.435 112.800 208.605 ;
        RECT 112.630 204.045 112.800 204.215 ;
        RECT 112.630 203.685 112.800 203.855 ;
        RECT 112.630 203.325 112.800 203.495 ;
        RECT 112.630 202.965 112.800 203.135 ;
        RECT 112.630 198.575 112.800 198.745 ;
        RECT 112.630 198.215 112.800 198.385 ;
        RECT 112.630 197.855 112.800 198.025 ;
        RECT 112.630 197.495 112.800 197.665 ;
        RECT 112.630 193.105 112.800 193.275 ;
        RECT 123.210 214.625 123.380 214.795 ;
        RECT 123.210 214.265 123.380 214.435 ;
        RECT 123.210 213.905 123.380 214.075 ;
        RECT 123.210 209.515 123.380 209.685 ;
        RECT 123.210 209.155 123.380 209.325 ;
        RECT 123.210 208.795 123.380 208.965 ;
        RECT 123.210 208.435 123.380 208.605 ;
        RECT 123.210 204.045 123.380 204.215 ;
        RECT 123.210 203.685 123.380 203.855 ;
        RECT 123.210 203.325 123.380 203.495 ;
        RECT 123.210 202.965 123.380 203.135 ;
        RECT 123.210 198.575 123.380 198.745 ;
        RECT 123.210 198.215 123.380 198.385 ;
        RECT 123.210 197.855 123.380 198.025 ;
        RECT 123.210 197.495 123.380 197.665 ;
        RECT 123.210 193.105 123.380 193.275 ;
        RECT 133.790 214.625 133.960 214.795 ;
        RECT 133.790 214.265 133.960 214.435 ;
        RECT 133.790 213.905 133.960 214.075 ;
        RECT 133.790 209.515 133.960 209.685 ;
        RECT 133.790 209.155 133.960 209.325 ;
        RECT 133.790 208.795 133.960 208.965 ;
        RECT 133.790 208.435 133.960 208.605 ;
        RECT 133.790 204.045 133.960 204.215 ;
        RECT 133.790 203.685 133.960 203.855 ;
        RECT 133.790 203.325 133.960 203.495 ;
        RECT 133.790 202.965 133.960 203.135 ;
        RECT 133.790 198.575 133.960 198.745 ;
        RECT 133.790 198.215 133.960 198.385 ;
        RECT 133.790 197.855 133.960 198.025 ;
        RECT 133.790 197.495 133.960 197.665 ;
        RECT 133.790 193.105 133.960 193.275 ;
        RECT 145.240 214.705 145.410 214.875 ;
        RECT 155.820 215.065 155.990 215.235 ;
        RECT 166.400 215.065 166.570 215.235 ;
        RECT 177.790 215.095 177.960 215.265 ;
        RECT 145.240 214.345 145.410 214.515 ;
        RECT 145.240 213.985 145.410 214.155 ;
        RECT 145.240 209.595 145.410 209.765 ;
        RECT 145.240 209.235 145.410 209.405 ;
        RECT 145.240 208.875 145.410 209.045 ;
        RECT 145.240 208.515 145.410 208.685 ;
        RECT 145.240 204.125 145.410 204.295 ;
        RECT 145.240 203.765 145.410 203.935 ;
        RECT 145.240 203.405 145.410 203.575 ;
        RECT 145.240 203.045 145.410 203.215 ;
        RECT 145.240 198.655 145.410 198.825 ;
        RECT 145.240 198.295 145.410 198.465 ;
        RECT 145.240 197.935 145.410 198.105 ;
        RECT 145.240 197.575 145.410 197.745 ;
        RECT 145.240 193.185 145.410 193.355 ;
        RECT 112.630 192.745 112.800 192.915 ;
        RECT 112.630 192.385 112.800 192.555 ;
        RECT 123.210 192.745 123.380 192.915 ;
        RECT 155.820 214.705 155.990 214.875 ;
        RECT 155.820 214.345 155.990 214.515 ;
        RECT 155.820 213.985 155.990 214.155 ;
        RECT 155.820 209.595 155.990 209.765 ;
        RECT 155.820 209.235 155.990 209.405 ;
        RECT 155.820 208.875 155.990 209.045 ;
        RECT 155.820 208.515 155.990 208.685 ;
        RECT 155.820 204.125 155.990 204.295 ;
        RECT 155.820 203.765 155.990 203.935 ;
        RECT 155.820 203.405 155.990 203.575 ;
        RECT 155.820 203.045 155.990 203.215 ;
        RECT 155.820 198.655 155.990 198.825 ;
        RECT 155.820 198.295 155.990 198.465 ;
        RECT 155.820 197.935 155.990 198.105 ;
        RECT 155.820 197.575 155.990 197.745 ;
        RECT 155.820 193.185 155.990 193.355 ;
        RECT 166.400 214.705 166.570 214.875 ;
        RECT 166.400 214.345 166.570 214.515 ;
        RECT 166.400 213.985 166.570 214.155 ;
        RECT 166.400 209.595 166.570 209.765 ;
        RECT 166.400 209.235 166.570 209.405 ;
        RECT 166.400 208.875 166.570 209.045 ;
        RECT 166.400 208.515 166.570 208.685 ;
        RECT 166.400 204.125 166.570 204.295 ;
        RECT 166.400 203.765 166.570 203.935 ;
        RECT 166.400 203.405 166.570 203.575 ;
        RECT 166.400 203.045 166.570 203.215 ;
        RECT 166.400 198.655 166.570 198.825 ;
        RECT 166.400 198.295 166.570 198.465 ;
        RECT 166.400 197.935 166.570 198.105 ;
        RECT 166.400 197.575 166.570 197.745 ;
        RECT 166.400 193.185 166.570 193.355 ;
        RECT 177.790 214.735 177.960 214.905 ;
        RECT 188.370 215.095 188.540 215.265 ;
        RECT 198.950 215.095 199.120 215.265 ;
        RECT 177.790 214.375 177.960 214.545 ;
        RECT 177.790 214.015 177.960 214.185 ;
        RECT 177.790 209.625 177.960 209.795 ;
        RECT 177.790 209.265 177.960 209.435 ;
        RECT 177.790 208.905 177.960 209.075 ;
        RECT 177.790 208.545 177.960 208.715 ;
        RECT 177.790 204.155 177.960 204.325 ;
        RECT 177.790 203.795 177.960 203.965 ;
        RECT 177.790 203.435 177.960 203.605 ;
        RECT 177.790 203.075 177.960 203.245 ;
        RECT 177.790 198.685 177.960 198.855 ;
        RECT 177.790 198.325 177.960 198.495 ;
        RECT 177.790 197.965 177.960 198.135 ;
        RECT 177.790 197.605 177.960 197.775 ;
        RECT 177.790 193.215 177.960 193.385 ;
        RECT 133.790 192.745 133.960 192.915 ;
        RECT 145.240 192.825 145.410 192.995 ;
        RECT 123.210 192.385 123.380 192.555 ;
        RECT 133.790 192.385 133.960 192.555 ;
        RECT 112.630 192.025 112.800 192.195 ;
        RECT 123.210 192.025 123.380 192.195 ;
        RECT 133.790 192.025 133.960 192.195 ;
        RECT 145.240 192.465 145.410 192.635 ;
        RECT 155.820 192.825 155.990 192.995 ;
        RECT 155.820 192.465 155.990 192.635 ;
        RECT 188.370 214.735 188.540 214.905 ;
        RECT 188.370 214.375 188.540 214.545 ;
        RECT 188.370 214.015 188.540 214.185 ;
        RECT 198.950 214.735 199.120 214.905 ;
        RECT 198.950 214.375 199.120 214.545 ;
        RECT 198.950 214.015 199.120 214.185 ;
        RECT 188.370 209.625 188.540 209.795 ;
        RECT 188.370 209.265 188.540 209.435 ;
        RECT 188.370 208.905 188.540 209.075 ;
        RECT 188.370 208.545 188.540 208.715 ;
        RECT 188.370 204.155 188.540 204.325 ;
        RECT 188.370 203.795 188.540 203.965 ;
        RECT 188.370 203.435 188.540 203.605 ;
        RECT 188.370 203.075 188.540 203.245 ;
        RECT 188.370 198.685 188.540 198.855 ;
        RECT 188.370 198.325 188.540 198.495 ;
        RECT 188.370 197.965 188.540 198.135 ;
        RECT 188.370 197.605 188.540 197.775 ;
        RECT 188.370 193.215 188.540 193.385 ;
        RECT 198.950 209.625 199.120 209.795 ;
        RECT 198.950 209.265 199.120 209.435 ;
        RECT 198.950 208.905 199.120 209.075 ;
        RECT 198.950 208.545 199.120 208.715 ;
        RECT 198.950 204.155 199.120 204.325 ;
        RECT 198.950 203.795 199.120 203.965 ;
        RECT 198.950 203.435 199.120 203.605 ;
        RECT 198.950 203.075 199.120 203.245 ;
        RECT 198.950 198.685 199.120 198.855 ;
        RECT 198.950 198.325 199.120 198.495 ;
        RECT 198.950 197.965 199.120 198.135 ;
        RECT 198.950 197.605 199.120 197.775 ;
        RECT 198.950 193.215 199.120 193.385 ;
        RECT 166.400 192.825 166.570 192.995 ;
        RECT 166.400 192.465 166.570 192.635 ;
        RECT 177.790 192.855 177.960 193.025 ;
        RECT 177.790 192.495 177.960 192.665 ;
        RECT 188.370 192.855 188.540 193.025 ;
        RECT 145.240 192.105 145.410 192.275 ;
        RECT 155.820 192.105 155.990 192.275 ;
        RECT 166.400 192.105 166.570 192.275 ;
        RECT 188.370 192.495 188.540 192.665 ;
        RECT 198.950 192.855 199.120 193.025 ;
        RECT 198.950 192.495 199.120 192.665 ;
        RECT 177.790 192.135 177.960 192.305 ;
        RECT 188.370 192.135 188.540 192.305 ;
        RECT 198.950 192.135 199.120 192.305 ;
        RECT 112.630 185.905 112.800 186.075 ;
        RECT 112.630 185.545 112.800 185.715 ;
        RECT 123.210 185.905 123.380 186.075 ;
        RECT 133.790 185.905 133.960 186.075 ;
        RECT 112.630 185.185 112.800 185.355 ;
        RECT 112.630 184.825 112.800 184.995 ;
        RECT 112.630 180.435 112.800 180.605 ;
        RECT 112.630 180.075 112.800 180.245 ;
        RECT 112.630 179.715 112.800 179.885 ;
        RECT 112.630 179.355 112.800 179.525 ;
        RECT 112.630 174.965 112.800 175.135 ;
        RECT 112.630 174.605 112.800 174.775 ;
        RECT 112.630 174.245 112.800 174.415 ;
        RECT 112.630 173.885 112.800 174.055 ;
        RECT 112.630 169.495 112.800 169.665 ;
        RECT 112.630 169.135 112.800 169.305 ;
        RECT 112.630 168.775 112.800 168.945 ;
        RECT 112.630 168.415 112.800 168.585 ;
        RECT 112.630 164.025 112.800 164.195 ;
        RECT 123.210 185.545 123.380 185.715 ;
        RECT 145.240 185.985 145.410 186.155 ;
        RECT 123.210 185.185 123.380 185.355 ;
        RECT 123.210 184.825 123.380 184.995 ;
        RECT 123.210 180.435 123.380 180.605 ;
        RECT 123.210 180.075 123.380 180.245 ;
        RECT 123.210 179.715 123.380 179.885 ;
        RECT 123.210 179.355 123.380 179.525 ;
        RECT 123.210 174.965 123.380 175.135 ;
        RECT 123.210 174.605 123.380 174.775 ;
        RECT 123.210 174.245 123.380 174.415 ;
        RECT 123.210 173.885 123.380 174.055 ;
        RECT 123.210 169.495 123.380 169.665 ;
        RECT 123.210 169.135 123.380 169.305 ;
        RECT 123.210 168.775 123.380 168.945 ;
        RECT 123.210 168.415 123.380 168.585 ;
        RECT 123.210 164.025 123.380 164.195 ;
        RECT 133.790 185.545 133.960 185.715 ;
        RECT 145.240 185.625 145.410 185.795 ;
        RECT 155.820 185.985 155.990 186.155 ;
        RECT 166.400 185.985 166.570 186.155 ;
        RECT 133.790 185.185 133.960 185.355 ;
        RECT 133.790 184.825 133.960 184.995 ;
        RECT 133.790 180.435 133.960 180.605 ;
        RECT 133.790 180.075 133.960 180.245 ;
        RECT 133.790 179.715 133.960 179.885 ;
        RECT 133.790 179.355 133.960 179.525 ;
        RECT 133.790 174.965 133.960 175.135 ;
        RECT 133.790 174.605 133.960 174.775 ;
        RECT 133.790 174.245 133.960 174.415 ;
        RECT 133.790 173.885 133.960 174.055 ;
        RECT 133.790 169.495 133.960 169.665 ;
        RECT 133.790 169.135 133.960 169.305 ;
        RECT 133.790 168.775 133.960 168.945 ;
        RECT 133.790 168.415 133.960 168.585 ;
        RECT 133.790 164.025 133.960 164.195 ;
        RECT 145.240 185.265 145.410 185.435 ;
        RECT 145.240 184.905 145.410 185.075 ;
        RECT 145.240 180.515 145.410 180.685 ;
        RECT 145.240 180.155 145.410 180.325 ;
        RECT 145.240 179.795 145.410 179.965 ;
        RECT 145.240 179.435 145.410 179.605 ;
        RECT 145.240 175.045 145.410 175.215 ;
        RECT 145.240 174.685 145.410 174.855 ;
        RECT 145.240 174.325 145.410 174.495 ;
        RECT 145.240 173.965 145.410 174.135 ;
        RECT 145.240 169.575 145.410 169.745 ;
        RECT 145.240 169.215 145.410 169.385 ;
        RECT 145.240 168.855 145.410 169.025 ;
        RECT 145.240 168.495 145.410 168.665 ;
        RECT 145.240 164.105 145.410 164.275 ;
        RECT 112.630 163.665 112.800 163.835 ;
        RECT 112.630 163.305 112.800 163.475 ;
        RECT 123.210 163.665 123.380 163.835 ;
        RECT 123.210 163.305 123.380 163.475 ;
        RECT 155.820 185.625 155.990 185.795 ;
        RECT 155.820 185.265 155.990 185.435 ;
        RECT 177.790 186.015 177.960 186.185 ;
        RECT 166.400 185.625 166.570 185.795 ;
        RECT 155.820 184.905 155.990 185.075 ;
        RECT 155.820 180.515 155.990 180.685 ;
        RECT 155.820 180.155 155.990 180.325 ;
        RECT 155.820 179.795 155.990 179.965 ;
        RECT 155.820 179.435 155.990 179.605 ;
        RECT 155.820 175.045 155.990 175.215 ;
        RECT 155.820 174.685 155.990 174.855 ;
        RECT 155.820 174.325 155.990 174.495 ;
        RECT 155.820 173.965 155.990 174.135 ;
        RECT 155.820 169.575 155.990 169.745 ;
        RECT 155.820 169.215 155.990 169.385 ;
        RECT 155.820 168.855 155.990 169.025 ;
        RECT 155.820 168.495 155.990 168.665 ;
        RECT 155.820 164.105 155.990 164.275 ;
        RECT 166.400 185.265 166.570 185.435 ;
        RECT 177.790 185.655 177.960 185.825 ;
        RECT 188.370 186.015 188.540 186.185 ;
        RECT 198.950 186.015 199.120 186.185 ;
        RECT 166.400 184.905 166.570 185.075 ;
        RECT 166.400 180.515 166.570 180.685 ;
        RECT 166.400 180.155 166.570 180.325 ;
        RECT 166.400 179.795 166.570 179.965 ;
        RECT 166.400 179.435 166.570 179.605 ;
        RECT 166.400 175.045 166.570 175.215 ;
        RECT 166.400 174.685 166.570 174.855 ;
        RECT 166.400 174.325 166.570 174.495 ;
        RECT 166.400 173.965 166.570 174.135 ;
        RECT 166.400 169.575 166.570 169.745 ;
        RECT 166.400 169.215 166.570 169.385 ;
        RECT 166.400 168.855 166.570 169.025 ;
        RECT 166.400 168.495 166.570 168.665 ;
        RECT 166.400 164.105 166.570 164.275 ;
        RECT 177.790 185.295 177.960 185.465 ;
        RECT 177.790 184.935 177.960 185.105 ;
        RECT 177.790 180.545 177.960 180.715 ;
        RECT 177.790 180.185 177.960 180.355 ;
        RECT 177.790 179.825 177.960 179.995 ;
        RECT 177.790 179.465 177.960 179.635 ;
        RECT 177.790 175.075 177.960 175.245 ;
        RECT 177.790 174.715 177.960 174.885 ;
        RECT 177.790 174.355 177.960 174.525 ;
        RECT 177.790 173.995 177.960 174.165 ;
        RECT 177.790 169.605 177.960 169.775 ;
        RECT 177.790 169.245 177.960 169.415 ;
        RECT 177.790 168.885 177.960 169.055 ;
        RECT 177.790 168.525 177.960 168.695 ;
        RECT 177.790 164.135 177.960 164.305 ;
        RECT 133.790 163.665 133.960 163.835 ;
        RECT 133.790 163.305 133.960 163.475 ;
        RECT 145.240 163.745 145.410 163.915 ;
        RECT 145.240 163.385 145.410 163.555 ;
        RECT 155.820 163.745 155.990 163.915 ;
        RECT 112.630 162.945 112.800 163.115 ;
        RECT 123.210 162.945 123.380 163.115 ;
        RECT 133.790 162.945 133.960 163.115 ;
        RECT 155.820 163.385 155.990 163.555 ;
        RECT 188.370 185.655 188.540 185.825 ;
        RECT 198.950 185.655 199.120 185.825 ;
        RECT 188.370 185.295 188.540 185.465 ;
        RECT 188.370 184.935 188.540 185.105 ;
        RECT 188.370 180.545 188.540 180.715 ;
        RECT 188.370 180.185 188.540 180.355 ;
        RECT 188.370 179.825 188.540 179.995 ;
        RECT 188.370 179.465 188.540 179.635 ;
        RECT 188.370 175.075 188.540 175.245 ;
        RECT 188.370 174.715 188.540 174.885 ;
        RECT 188.370 174.355 188.540 174.525 ;
        RECT 188.370 173.995 188.540 174.165 ;
        RECT 188.370 169.605 188.540 169.775 ;
        RECT 188.370 169.245 188.540 169.415 ;
        RECT 188.370 168.885 188.540 169.055 ;
        RECT 188.370 168.525 188.540 168.695 ;
        RECT 188.370 164.135 188.540 164.305 ;
        RECT 198.950 185.295 199.120 185.465 ;
        RECT 198.950 184.935 199.120 185.105 ;
        RECT 198.950 180.545 199.120 180.715 ;
        RECT 198.950 180.185 199.120 180.355 ;
        RECT 198.950 179.825 199.120 179.995 ;
        RECT 198.950 179.465 199.120 179.635 ;
        RECT 198.950 175.075 199.120 175.245 ;
        RECT 198.950 174.715 199.120 174.885 ;
        RECT 198.950 174.355 199.120 174.525 ;
        RECT 198.950 173.995 199.120 174.165 ;
        RECT 198.950 169.605 199.120 169.775 ;
        RECT 198.950 169.245 199.120 169.415 ;
        RECT 198.950 168.885 199.120 169.055 ;
        RECT 198.950 168.525 199.120 168.695 ;
        RECT 198.950 164.135 199.120 164.305 ;
        RECT 166.400 163.745 166.570 163.915 ;
        RECT 166.400 163.385 166.570 163.555 ;
        RECT 177.790 163.775 177.960 163.945 ;
        RECT 177.790 163.415 177.960 163.585 ;
        RECT 188.370 163.775 188.540 163.945 ;
        RECT 145.240 163.025 145.410 163.195 ;
        RECT 188.370 163.415 188.540 163.585 ;
        RECT 198.950 163.775 199.120 163.945 ;
        RECT 198.950 163.415 199.120 163.585 ;
        RECT 155.820 163.025 155.990 163.195 ;
        RECT 166.400 163.025 166.570 163.195 ;
        RECT 177.790 163.055 177.960 163.225 ;
        RECT 188.370 163.055 188.540 163.225 ;
        RECT 198.950 163.055 199.120 163.225 ;
        RECT 112.630 156.735 112.800 156.905 ;
        RECT 112.630 156.375 112.800 156.545 ;
        RECT 123.210 156.735 123.380 156.905 ;
        RECT 133.790 156.735 133.960 156.905 ;
        RECT 112.630 156.015 112.800 156.185 ;
        RECT 112.630 155.655 112.800 155.825 ;
        RECT 112.630 151.265 112.800 151.435 ;
        RECT 112.630 150.905 112.800 151.075 ;
        RECT 112.630 150.545 112.800 150.715 ;
        RECT 112.630 150.185 112.800 150.355 ;
        RECT 112.630 145.795 112.800 145.965 ;
        RECT 112.630 145.435 112.800 145.605 ;
        RECT 112.630 145.075 112.800 145.245 ;
        RECT 112.630 144.715 112.800 144.885 ;
        RECT 112.630 140.325 112.800 140.495 ;
        RECT 112.630 139.965 112.800 140.135 ;
        RECT 112.630 139.605 112.800 139.775 ;
        RECT 112.630 139.245 112.800 139.415 ;
        RECT 112.630 134.855 112.800 135.025 ;
        RECT 123.210 156.375 123.380 156.545 ;
        RECT 145.240 156.815 145.410 156.985 ;
        RECT 133.790 156.375 133.960 156.545 ;
        RECT 145.240 156.455 145.410 156.625 ;
        RECT 155.820 156.815 155.990 156.985 ;
        RECT 166.400 156.815 166.570 156.985 ;
        RECT 123.210 156.015 123.380 156.185 ;
        RECT 123.210 155.655 123.380 155.825 ;
        RECT 123.210 151.265 123.380 151.435 ;
        RECT 123.210 150.905 123.380 151.075 ;
        RECT 123.210 150.545 123.380 150.715 ;
        RECT 123.210 150.185 123.380 150.355 ;
        RECT 123.210 145.795 123.380 145.965 ;
        RECT 123.210 145.435 123.380 145.605 ;
        RECT 123.210 145.075 123.380 145.245 ;
        RECT 123.210 144.715 123.380 144.885 ;
        RECT 123.210 140.325 123.380 140.495 ;
        RECT 123.210 139.965 123.380 140.135 ;
        RECT 123.210 139.605 123.380 139.775 ;
        RECT 123.210 139.245 123.380 139.415 ;
        RECT 123.210 134.855 123.380 135.025 ;
        RECT 133.790 156.015 133.960 156.185 ;
        RECT 133.790 155.655 133.960 155.825 ;
        RECT 133.790 151.265 133.960 151.435 ;
        RECT 133.790 150.905 133.960 151.075 ;
        RECT 133.790 150.545 133.960 150.715 ;
        RECT 133.790 150.185 133.960 150.355 ;
        RECT 133.790 145.795 133.960 145.965 ;
        RECT 133.790 145.435 133.960 145.605 ;
        RECT 133.790 145.075 133.960 145.245 ;
        RECT 133.790 144.715 133.960 144.885 ;
        RECT 133.790 140.325 133.960 140.495 ;
        RECT 133.790 139.965 133.960 140.135 ;
        RECT 133.790 139.605 133.960 139.775 ;
        RECT 133.790 139.245 133.960 139.415 ;
        RECT 133.790 134.855 133.960 135.025 ;
        RECT 145.240 156.095 145.410 156.265 ;
        RECT 145.240 155.735 145.410 155.905 ;
        RECT 145.240 151.345 145.410 151.515 ;
        RECT 145.240 150.985 145.410 151.155 ;
        RECT 145.240 150.625 145.410 150.795 ;
        RECT 145.240 150.265 145.410 150.435 ;
        RECT 145.240 145.875 145.410 146.045 ;
        RECT 145.240 145.515 145.410 145.685 ;
        RECT 145.240 145.155 145.410 145.325 ;
        RECT 145.240 144.795 145.410 144.965 ;
        RECT 145.240 140.405 145.410 140.575 ;
        RECT 145.240 140.045 145.410 140.215 ;
        RECT 145.240 139.685 145.410 139.855 ;
        RECT 145.240 139.325 145.410 139.495 ;
        RECT 145.240 134.935 145.410 135.105 ;
        RECT 112.630 134.495 112.800 134.665 ;
        RECT 112.630 134.135 112.800 134.305 ;
        RECT 123.210 134.495 123.380 134.665 ;
        RECT 155.820 156.455 155.990 156.625 ;
        RECT 155.820 156.095 155.990 156.265 ;
        RECT 177.790 156.845 177.960 157.015 ;
        RECT 166.400 156.455 166.570 156.625 ;
        RECT 155.820 155.735 155.990 155.905 ;
        RECT 155.820 151.345 155.990 151.515 ;
        RECT 155.820 150.985 155.990 151.155 ;
        RECT 155.820 150.625 155.990 150.795 ;
        RECT 155.820 150.265 155.990 150.435 ;
        RECT 155.820 145.875 155.990 146.045 ;
        RECT 155.820 145.515 155.990 145.685 ;
        RECT 155.820 145.155 155.990 145.325 ;
        RECT 155.820 144.795 155.990 144.965 ;
        RECT 155.820 140.405 155.990 140.575 ;
        RECT 155.820 140.045 155.990 140.215 ;
        RECT 155.820 139.685 155.990 139.855 ;
        RECT 155.820 139.325 155.990 139.495 ;
        RECT 155.820 134.935 155.990 135.105 ;
        RECT 166.400 156.095 166.570 156.265 ;
        RECT 177.790 156.485 177.960 156.655 ;
        RECT 188.370 156.845 188.540 157.015 ;
        RECT 198.950 156.845 199.120 157.015 ;
        RECT 166.400 155.735 166.570 155.905 ;
        RECT 166.400 151.345 166.570 151.515 ;
        RECT 166.400 150.985 166.570 151.155 ;
        RECT 166.400 150.625 166.570 150.795 ;
        RECT 166.400 150.265 166.570 150.435 ;
        RECT 166.400 145.875 166.570 146.045 ;
        RECT 166.400 145.515 166.570 145.685 ;
        RECT 166.400 145.155 166.570 145.325 ;
        RECT 166.400 144.795 166.570 144.965 ;
        RECT 166.400 140.405 166.570 140.575 ;
        RECT 166.400 140.045 166.570 140.215 ;
        RECT 166.400 139.685 166.570 139.855 ;
        RECT 166.400 139.325 166.570 139.495 ;
        RECT 166.400 134.935 166.570 135.105 ;
        RECT 177.790 156.125 177.960 156.295 ;
        RECT 177.790 155.765 177.960 155.935 ;
        RECT 177.790 151.375 177.960 151.545 ;
        RECT 177.790 151.015 177.960 151.185 ;
        RECT 177.790 150.655 177.960 150.825 ;
        RECT 177.790 150.295 177.960 150.465 ;
        RECT 177.790 145.905 177.960 146.075 ;
        RECT 177.790 145.545 177.960 145.715 ;
        RECT 177.790 145.185 177.960 145.355 ;
        RECT 177.790 144.825 177.960 144.995 ;
        RECT 177.790 140.435 177.960 140.605 ;
        RECT 177.790 140.075 177.960 140.245 ;
        RECT 177.790 139.715 177.960 139.885 ;
        RECT 177.790 139.355 177.960 139.525 ;
        RECT 177.790 134.965 177.960 135.135 ;
        RECT 133.790 134.495 133.960 134.665 ;
        RECT 145.240 134.575 145.410 134.745 ;
        RECT 123.210 134.135 123.380 134.305 ;
        RECT 133.790 134.135 133.960 134.305 ;
        RECT 112.630 133.775 112.800 133.945 ;
        RECT 123.210 133.775 123.380 133.945 ;
        RECT 133.790 133.775 133.960 133.945 ;
        RECT 145.240 134.215 145.410 134.385 ;
        RECT 155.820 134.575 155.990 134.745 ;
        RECT 155.820 134.215 155.990 134.385 ;
        RECT 188.370 156.485 188.540 156.655 ;
        RECT 188.370 156.125 188.540 156.295 ;
        RECT 188.370 155.765 188.540 155.935 ;
        RECT 188.370 151.375 188.540 151.545 ;
        RECT 188.370 151.015 188.540 151.185 ;
        RECT 188.370 150.655 188.540 150.825 ;
        RECT 188.370 150.295 188.540 150.465 ;
        RECT 188.370 145.905 188.540 146.075 ;
        RECT 188.370 145.545 188.540 145.715 ;
        RECT 188.370 145.185 188.540 145.355 ;
        RECT 188.370 144.825 188.540 144.995 ;
        RECT 188.370 140.435 188.540 140.605 ;
        RECT 188.370 140.075 188.540 140.245 ;
        RECT 188.370 139.715 188.540 139.885 ;
        RECT 188.370 139.355 188.540 139.525 ;
        RECT 188.370 134.965 188.540 135.135 ;
        RECT 198.950 156.485 199.120 156.655 ;
        RECT 198.950 156.125 199.120 156.295 ;
        RECT 198.950 155.765 199.120 155.935 ;
        RECT 198.950 151.375 199.120 151.545 ;
        RECT 198.950 151.015 199.120 151.185 ;
        RECT 198.950 150.655 199.120 150.825 ;
        RECT 198.950 150.295 199.120 150.465 ;
        RECT 198.950 145.905 199.120 146.075 ;
        RECT 198.950 145.545 199.120 145.715 ;
        RECT 198.950 145.185 199.120 145.355 ;
        RECT 198.950 144.825 199.120 144.995 ;
        RECT 198.950 140.435 199.120 140.605 ;
        RECT 198.950 140.075 199.120 140.245 ;
        RECT 198.950 139.715 199.120 139.885 ;
        RECT 198.950 139.355 199.120 139.525 ;
        RECT 198.950 134.965 199.120 135.135 ;
        RECT 166.400 134.575 166.570 134.745 ;
        RECT 166.400 134.215 166.570 134.385 ;
        RECT 177.790 134.605 177.960 134.775 ;
        RECT 177.790 134.245 177.960 134.415 ;
        RECT 188.370 134.605 188.540 134.775 ;
        RECT 145.240 133.855 145.410 134.025 ;
        RECT 155.820 133.855 155.990 134.025 ;
        RECT 166.400 133.855 166.570 134.025 ;
        RECT 188.370 134.245 188.540 134.415 ;
        RECT 198.950 134.605 199.120 134.775 ;
        RECT 198.950 134.245 199.120 134.415 ;
        RECT 177.790 133.885 177.960 134.055 ;
        RECT 188.370 133.885 188.540 134.055 ;
        RECT 198.950 133.885 199.120 134.055 ;
        RECT 112.630 127.555 112.800 127.725 ;
        RECT 112.630 127.195 112.800 127.365 ;
        RECT 123.210 127.555 123.380 127.725 ;
        RECT 133.790 127.555 133.960 127.725 ;
        RECT 112.630 126.835 112.800 127.005 ;
        RECT 112.630 126.475 112.800 126.645 ;
        RECT 112.630 122.085 112.800 122.255 ;
        RECT 112.630 121.725 112.800 121.895 ;
        RECT 112.630 121.365 112.800 121.535 ;
        RECT 112.630 121.005 112.800 121.175 ;
        RECT 112.630 116.615 112.800 116.785 ;
        RECT 112.630 116.255 112.800 116.425 ;
        RECT 112.630 115.895 112.800 116.065 ;
        RECT 112.630 115.535 112.800 115.705 ;
        RECT 112.630 111.145 112.800 111.315 ;
        RECT 112.630 110.785 112.800 110.955 ;
        RECT 112.630 110.425 112.800 110.595 ;
        RECT 112.630 110.065 112.800 110.235 ;
        RECT 112.630 105.675 112.800 105.845 ;
        RECT 123.210 127.195 123.380 127.365 ;
        RECT 145.240 127.635 145.410 127.805 ;
        RECT 123.210 126.835 123.380 127.005 ;
        RECT 123.210 126.475 123.380 126.645 ;
        RECT 123.210 122.085 123.380 122.255 ;
        RECT 123.210 121.725 123.380 121.895 ;
        RECT 123.210 121.365 123.380 121.535 ;
        RECT 123.210 121.005 123.380 121.175 ;
        RECT 123.210 116.615 123.380 116.785 ;
        RECT 123.210 116.255 123.380 116.425 ;
        RECT 123.210 115.895 123.380 116.065 ;
        RECT 123.210 115.535 123.380 115.705 ;
        RECT 123.210 111.145 123.380 111.315 ;
        RECT 123.210 110.785 123.380 110.955 ;
        RECT 123.210 110.425 123.380 110.595 ;
        RECT 123.210 110.065 123.380 110.235 ;
        RECT 123.210 105.675 123.380 105.845 ;
        RECT 133.790 127.195 133.960 127.365 ;
        RECT 133.790 126.835 133.960 127.005 ;
        RECT 133.790 126.475 133.960 126.645 ;
        RECT 133.790 122.085 133.960 122.255 ;
        RECT 133.790 121.725 133.960 121.895 ;
        RECT 133.790 121.365 133.960 121.535 ;
        RECT 133.790 121.005 133.960 121.175 ;
        RECT 133.790 116.615 133.960 116.785 ;
        RECT 133.790 116.255 133.960 116.425 ;
        RECT 133.790 115.895 133.960 116.065 ;
        RECT 133.790 115.535 133.960 115.705 ;
        RECT 133.790 111.145 133.960 111.315 ;
        RECT 133.790 110.785 133.960 110.955 ;
        RECT 133.790 110.425 133.960 110.595 ;
        RECT 133.790 110.065 133.960 110.235 ;
        RECT 133.790 105.675 133.960 105.845 ;
        RECT 145.240 127.275 145.410 127.445 ;
        RECT 155.820 127.635 155.990 127.805 ;
        RECT 166.400 127.635 166.570 127.805 ;
        RECT 145.240 126.915 145.410 127.085 ;
        RECT 145.240 126.555 145.410 126.725 ;
        RECT 145.240 122.165 145.410 122.335 ;
        RECT 145.240 121.805 145.410 121.975 ;
        RECT 145.240 121.445 145.410 121.615 ;
        RECT 145.240 121.085 145.410 121.255 ;
        RECT 145.240 116.695 145.410 116.865 ;
        RECT 145.240 116.335 145.410 116.505 ;
        RECT 145.240 115.975 145.410 116.145 ;
        RECT 145.240 115.615 145.410 115.785 ;
        RECT 145.240 111.225 145.410 111.395 ;
        RECT 145.240 110.865 145.410 111.035 ;
        RECT 145.240 110.505 145.410 110.675 ;
        RECT 145.240 110.145 145.410 110.315 ;
        RECT 145.240 105.755 145.410 105.925 ;
        RECT 112.630 105.315 112.800 105.485 ;
        RECT 112.630 104.955 112.800 105.125 ;
        RECT 123.210 105.315 123.380 105.485 ;
        RECT 123.210 104.955 123.380 105.125 ;
        RECT 155.820 127.275 155.990 127.445 ;
        RECT 177.790 127.665 177.960 127.835 ;
        RECT 166.400 127.275 166.570 127.445 ;
        RECT 177.790 127.305 177.960 127.475 ;
        RECT 188.370 127.665 188.540 127.835 ;
        RECT 198.950 127.665 199.120 127.835 ;
        RECT 155.820 126.915 155.990 127.085 ;
        RECT 155.820 126.555 155.990 126.725 ;
        RECT 155.820 122.165 155.990 122.335 ;
        RECT 155.820 121.805 155.990 121.975 ;
        RECT 155.820 121.445 155.990 121.615 ;
        RECT 155.820 121.085 155.990 121.255 ;
        RECT 155.820 116.695 155.990 116.865 ;
        RECT 155.820 116.335 155.990 116.505 ;
        RECT 155.820 115.975 155.990 116.145 ;
        RECT 155.820 115.615 155.990 115.785 ;
        RECT 155.820 111.225 155.990 111.395 ;
        RECT 155.820 110.865 155.990 111.035 ;
        RECT 155.820 110.505 155.990 110.675 ;
        RECT 155.820 110.145 155.990 110.315 ;
        RECT 155.820 105.755 155.990 105.925 ;
        RECT 166.400 126.915 166.570 127.085 ;
        RECT 166.400 126.555 166.570 126.725 ;
        RECT 166.400 122.165 166.570 122.335 ;
        RECT 166.400 121.805 166.570 121.975 ;
        RECT 166.400 121.445 166.570 121.615 ;
        RECT 166.400 121.085 166.570 121.255 ;
        RECT 166.400 116.695 166.570 116.865 ;
        RECT 166.400 116.335 166.570 116.505 ;
        RECT 166.400 115.975 166.570 116.145 ;
        RECT 166.400 115.615 166.570 115.785 ;
        RECT 166.400 111.225 166.570 111.395 ;
        RECT 166.400 110.865 166.570 111.035 ;
        RECT 166.400 110.505 166.570 110.675 ;
        RECT 166.400 110.145 166.570 110.315 ;
        RECT 166.400 105.755 166.570 105.925 ;
        RECT 177.790 126.945 177.960 127.115 ;
        RECT 177.790 126.585 177.960 126.755 ;
        RECT 177.790 122.195 177.960 122.365 ;
        RECT 177.790 121.835 177.960 122.005 ;
        RECT 177.790 121.475 177.960 121.645 ;
        RECT 177.790 121.115 177.960 121.285 ;
        RECT 177.790 116.725 177.960 116.895 ;
        RECT 177.790 116.365 177.960 116.535 ;
        RECT 177.790 116.005 177.960 116.175 ;
        RECT 177.790 115.645 177.960 115.815 ;
        RECT 177.790 111.255 177.960 111.425 ;
        RECT 177.790 110.895 177.960 111.065 ;
        RECT 177.790 110.535 177.960 110.705 ;
        RECT 177.790 110.175 177.960 110.345 ;
        RECT 177.790 105.785 177.960 105.955 ;
        RECT 133.790 105.315 133.960 105.485 ;
        RECT 133.790 104.955 133.960 105.125 ;
        RECT 145.240 105.395 145.410 105.565 ;
        RECT 145.240 105.035 145.410 105.205 ;
        RECT 155.820 105.395 155.990 105.565 ;
        RECT 112.630 104.595 112.800 104.765 ;
        RECT 123.210 104.595 123.380 104.765 ;
        RECT 133.790 104.595 133.960 104.765 ;
        RECT 155.820 105.035 155.990 105.205 ;
        RECT 188.370 127.305 188.540 127.475 ;
        RECT 188.370 126.945 188.540 127.115 ;
        RECT 198.950 127.305 199.120 127.475 ;
        RECT 198.950 126.945 199.120 127.115 ;
        RECT 376.340 127.425 376.510 127.595 ;
        RECT 386.920 127.425 387.090 127.595 ;
        RECT 397.500 127.425 397.670 127.595 ;
        RECT 376.340 127.065 376.510 127.235 ;
        RECT 408.650 127.415 408.820 127.585 ;
        RECT 188.370 126.585 188.540 126.755 ;
        RECT 188.370 122.195 188.540 122.365 ;
        RECT 188.370 121.835 188.540 122.005 ;
        RECT 188.370 121.475 188.540 121.645 ;
        RECT 188.370 121.115 188.540 121.285 ;
        RECT 188.370 116.725 188.540 116.895 ;
        RECT 188.370 116.365 188.540 116.535 ;
        RECT 188.370 116.005 188.540 116.175 ;
        RECT 188.370 115.645 188.540 115.815 ;
        RECT 188.370 111.255 188.540 111.425 ;
        RECT 188.370 110.895 188.540 111.065 ;
        RECT 188.370 110.535 188.540 110.705 ;
        RECT 188.370 110.175 188.540 110.345 ;
        RECT 188.370 105.785 188.540 105.955 ;
        RECT 198.950 126.585 199.120 126.755 ;
        RECT 198.950 122.195 199.120 122.365 ;
        RECT 198.950 121.835 199.120 122.005 ;
        RECT 198.950 121.475 199.120 121.645 ;
        RECT 198.950 121.115 199.120 121.285 ;
        RECT 198.950 116.725 199.120 116.895 ;
        RECT 198.950 116.365 199.120 116.535 ;
        RECT 198.950 116.005 199.120 116.175 ;
        RECT 198.950 115.645 199.120 115.815 ;
        RECT 198.950 111.255 199.120 111.425 ;
        RECT 198.950 110.895 199.120 111.065 ;
        RECT 198.950 110.535 199.120 110.705 ;
        RECT 198.950 110.175 199.120 110.345 ;
        RECT 198.950 105.785 199.120 105.955 ;
        RECT 376.340 126.705 376.510 126.875 ;
        RECT 376.340 126.345 376.510 126.515 ;
        RECT 386.920 127.065 387.090 127.235 ;
        RECT 386.920 126.705 387.090 126.875 ;
        RECT 386.920 126.345 387.090 126.515 ;
        RECT 376.340 121.955 376.510 122.125 ;
        RECT 376.340 121.595 376.510 121.765 ;
        RECT 376.340 121.235 376.510 121.405 ;
        RECT 376.340 120.875 376.510 121.045 ;
        RECT 386.920 121.955 387.090 122.125 ;
        RECT 386.920 121.595 387.090 121.765 ;
        RECT 386.920 121.235 387.090 121.405 ;
        RECT 386.920 120.875 387.090 121.045 ;
        RECT 376.340 116.485 376.510 116.655 ;
        RECT 376.340 116.125 376.510 116.295 ;
        RECT 376.340 115.765 376.510 115.935 ;
        RECT 376.340 115.405 376.510 115.575 ;
        RECT 386.920 116.485 387.090 116.655 ;
        RECT 386.920 116.125 387.090 116.295 ;
        RECT 386.920 115.765 387.090 115.935 ;
        RECT 386.920 115.405 387.090 115.575 ;
        RECT 376.340 111.015 376.510 111.185 ;
        RECT 376.340 110.655 376.510 110.825 ;
        RECT 376.340 110.295 376.510 110.465 ;
        RECT 376.340 109.935 376.510 110.105 ;
        RECT 386.920 111.015 387.090 111.185 ;
        RECT 386.920 110.655 387.090 110.825 ;
        RECT 386.920 110.295 387.090 110.465 ;
        RECT 386.920 109.935 387.090 110.105 ;
        RECT 166.400 105.395 166.570 105.565 ;
        RECT 166.400 105.035 166.570 105.205 ;
        RECT 177.790 105.425 177.960 105.595 ;
        RECT 177.790 105.065 177.960 105.235 ;
        RECT 188.370 105.425 188.540 105.595 ;
        RECT 145.240 104.675 145.410 104.845 ;
        RECT 155.820 104.675 155.990 104.845 ;
        RECT 166.400 104.675 166.570 104.845 ;
        RECT 188.370 105.065 188.540 105.235 ;
        RECT 198.950 105.425 199.120 105.595 ;
        RECT 376.340 105.545 376.510 105.715 ;
        RECT 386.920 105.545 387.090 105.715 ;
        RECT 397.500 127.065 397.670 127.235 ;
        RECT 397.500 126.705 397.670 126.875 ;
        RECT 397.500 126.345 397.670 126.515 ;
        RECT 397.500 121.955 397.670 122.125 ;
        RECT 397.500 121.595 397.670 121.765 ;
        RECT 397.500 121.235 397.670 121.405 ;
        RECT 397.500 120.875 397.670 121.045 ;
        RECT 397.500 116.485 397.670 116.655 ;
        RECT 397.500 116.125 397.670 116.295 ;
        RECT 397.500 115.765 397.670 115.935 ;
        RECT 397.500 115.405 397.670 115.575 ;
        RECT 397.500 111.015 397.670 111.185 ;
        RECT 397.500 110.655 397.670 110.825 ;
        RECT 397.500 110.295 397.670 110.465 ;
        RECT 397.500 109.935 397.670 110.105 ;
        RECT 397.500 105.545 397.670 105.715 ;
        RECT 419.230 127.415 419.400 127.585 ;
        RECT 429.810 127.415 429.980 127.585 ;
        RECT 408.650 127.055 408.820 127.225 ;
        RECT 408.650 126.695 408.820 126.865 ;
        RECT 408.650 126.335 408.820 126.505 ;
        RECT 419.230 127.055 419.400 127.225 ;
        RECT 419.230 126.695 419.400 126.865 ;
        RECT 419.230 126.335 419.400 126.505 ;
        RECT 408.650 121.945 408.820 122.115 ;
        RECT 408.650 121.585 408.820 121.755 ;
        RECT 408.650 121.225 408.820 121.395 ;
        RECT 408.650 120.865 408.820 121.035 ;
        RECT 419.230 121.945 419.400 122.115 ;
        RECT 419.230 121.585 419.400 121.755 ;
        RECT 419.230 121.225 419.400 121.395 ;
        RECT 419.230 120.865 419.400 121.035 ;
        RECT 408.650 116.475 408.820 116.645 ;
        RECT 408.650 116.115 408.820 116.285 ;
        RECT 408.650 115.755 408.820 115.925 ;
        RECT 408.650 115.395 408.820 115.565 ;
        RECT 419.230 116.475 419.400 116.645 ;
        RECT 419.230 116.115 419.400 116.285 ;
        RECT 419.230 115.755 419.400 115.925 ;
        RECT 419.230 115.395 419.400 115.565 ;
        RECT 408.650 111.005 408.820 111.175 ;
        RECT 408.650 110.645 408.820 110.815 ;
        RECT 408.650 110.285 408.820 110.455 ;
        RECT 408.650 109.925 408.820 110.095 ;
        RECT 419.230 111.005 419.400 111.175 ;
        RECT 419.230 110.645 419.400 110.815 ;
        RECT 419.230 110.285 419.400 110.455 ;
        RECT 419.230 109.925 419.400 110.095 ;
        RECT 198.950 105.065 199.120 105.235 ;
        RECT 376.340 105.185 376.510 105.355 ;
        RECT 177.790 104.705 177.960 104.875 ;
        RECT 188.370 104.705 188.540 104.875 ;
        RECT 198.950 104.705 199.120 104.875 ;
        RECT 376.340 104.825 376.510 104.995 ;
        RECT 376.340 104.465 376.510 104.635 ;
        RECT 386.920 105.185 387.090 105.355 ;
        RECT 386.920 104.825 387.090 104.995 ;
        RECT 386.920 104.465 387.090 104.635 ;
        RECT 408.650 105.535 408.820 105.705 ;
        RECT 419.230 105.535 419.400 105.705 ;
        RECT 429.810 127.055 429.980 127.225 ;
        RECT 429.810 126.695 429.980 126.865 ;
        RECT 429.810 126.335 429.980 126.505 ;
        RECT 429.810 121.945 429.980 122.115 ;
        RECT 429.810 121.585 429.980 121.755 ;
        RECT 429.810 121.225 429.980 121.395 ;
        RECT 429.810 120.865 429.980 121.035 ;
        RECT 429.810 116.475 429.980 116.645 ;
        RECT 429.810 116.115 429.980 116.285 ;
        RECT 429.810 115.755 429.980 115.925 ;
        RECT 429.810 115.395 429.980 115.565 ;
        RECT 429.810 111.005 429.980 111.175 ;
        RECT 429.810 110.645 429.980 110.815 ;
        RECT 429.810 110.285 429.980 110.455 ;
        RECT 429.810 109.925 429.980 110.095 ;
        RECT 429.810 105.535 429.980 105.705 ;
        RECT 397.500 105.185 397.670 105.355 ;
        RECT 397.500 104.825 397.670 104.995 ;
        RECT 397.500 104.465 397.670 104.635 ;
        RECT 408.650 105.175 408.820 105.345 ;
        RECT 408.650 104.815 408.820 104.985 ;
        RECT 408.650 104.455 408.820 104.625 ;
        RECT 419.230 105.175 419.400 105.345 ;
        RECT 419.230 104.815 419.400 104.985 ;
        RECT 419.230 104.455 419.400 104.625 ;
        RECT 429.810 105.175 429.980 105.345 ;
        RECT 429.810 104.815 429.980 104.985 ;
        RECT 429.810 104.455 429.980 104.625 ;
        RECT 112.630 98.235 112.800 98.405 ;
        RECT 112.630 97.875 112.800 98.045 ;
        RECT 123.210 98.235 123.380 98.405 ;
        RECT 133.790 98.235 133.960 98.405 ;
        RECT 112.630 97.515 112.800 97.685 ;
        RECT 112.630 97.155 112.800 97.325 ;
        RECT 112.630 92.765 112.800 92.935 ;
        RECT 112.630 92.405 112.800 92.575 ;
        RECT 112.630 92.045 112.800 92.215 ;
        RECT 112.630 91.685 112.800 91.855 ;
        RECT 112.630 87.295 112.800 87.465 ;
        RECT 112.630 86.935 112.800 87.105 ;
        RECT 112.630 86.575 112.800 86.745 ;
        RECT 112.630 86.215 112.800 86.385 ;
        RECT 112.630 81.825 112.800 81.995 ;
        RECT 112.630 81.465 112.800 81.635 ;
        RECT 112.630 81.105 112.800 81.275 ;
        RECT 112.630 80.745 112.800 80.915 ;
        RECT 112.630 76.355 112.800 76.525 ;
        RECT 123.210 97.875 123.380 98.045 ;
        RECT 145.240 98.315 145.410 98.485 ;
        RECT 123.210 97.515 123.380 97.685 ;
        RECT 123.210 97.155 123.380 97.325 ;
        RECT 123.210 92.765 123.380 92.935 ;
        RECT 123.210 92.405 123.380 92.575 ;
        RECT 123.210 92.045 123.380 92.215 ;
        RECT 123.210 91.685 123.380 91.855 ;
        RECT 123.210 87.295 123.380 87.465 ;
        RECT 123.210 86.935 123.380 87.105 ;
        RECT 123.210 86.575 123.380 86.745 ;
        RECT 123.210 86.215 123.380 86.385 ;
        RECT 123.210 81.825 123.380 81.995 ;
        RECT 123.210 81.465 123.380 81.635 ;
        RECT 123.210 81.105 123.380 81.275 ;
        RECT 123.210 80.745 123.380 80.915 ;
        RECT 123.210 76.355 123.380 76.525 ;
        RECT 133.790 97.875 133.960 98.045 ;
        RECT 133.790 97.515 133.960 97.685 ;
        RECT 133.790 97.155 133.960 97.325 ;
        RECT 133.790 92.765 133.960 92.935 ;
        RECT 133.790 92.405 133.960 92.575 ;
        RECT 133.790 92.045 133.960 92.215 ;
        RECT 133.790 91.685 133.960 91.855 ;
        RECT 133.790 87.295 133.960 87.465 ;
        RECT 133.790 86.935 133.960 87.105 ;
        RECT 133.790 86.575 133.960 86.745 ;
        RECT 133.790 86.215 133.960 86.385 ;
        RECT 133.790 81.825 133.960 81.995 ;
        RECT 133.790 81.465 133.960 81.635 ;
        RECT 133.790 81.105 133.960 81.275 ;
        RECT 133.790 80.745 133.960 80.915 ;
        RECT 133.790 76.355 133.960 76.525 ;
        RECT 145.240 97.955 145.410 98.125 ;
        RECT 155.820 98.315 155.990 98.485 ;
        RECT 166.400 98.315 166.570 98.485 ;
        RECT 145.240 97.595 145.410 97.765 ;
        RECT 145.240 97.235 145.410 97.405 ;
        RECT 145.240 92.845 145.410 93.015 ;
        RECT 145.240 92.485 145.410 92.655 ;
        RECT 145.240 92.125 145.410 92.295 ;
        RECT 145.240 91.765 145.410 91.935 ;
        RECT 145.240 87.375 145.410 87.545 ;
        RECT 145.240 87.015 145.410 87.185 ;
        RECT 145.240 86.655 145.410 86.825 ;
        RECT 145.240 86.295 145.410 86.465 ;
        RECT 145.240 81.905 145.410 82.075 ;
        RECT 145.240 81.545 145.410 81.715 ;
        RECT 145.240 81.185 145.410 81.355 ;
        RECT 145.240 80.825 145.410 80.995 ;
        RECT 145.240 76.435 145.410 76.605 ;
        RECT 112.630 75.995 112.800 76.165 ;
        RECT 112.630 75.635 112.800 75.805 ;
        RECT 123.210 75.995 123.380 76.165 ;
        RECT 123.210 75.635 123.380 75.805 ;
        RECT 155.820 97.955 155.990 98.125 ;
        RECT 177.790 98.345 177.960 98.515 ;
        RECT 166.400 97.955 166.570 98.125 ;
        RECT 177.790 97.985 177.960 98.155 ;
        RECT 188.370 98.345 188.540 98.515 ;
        RECT 198.950 98.345 199.120 98.515 ;
        RECT 155.820 97.595 155.990 97.765 ;
        RECT 155.820 97.235 155.990 97.405 ;
        RECT 155.820 92.845 155.990 93.015 ;
        RECT 155.820 92.485 155.990 92.655 ;
        RECT 155.820 92.125 155.990 92.295 ;
        RECT 155.820 91.765 155.990 91.935 ;
        RECT 155.820 87.375 155.990 87.545 ;
        RECT 155.820 87.015 155.990 87.185 ;
        RECT 155.820 86.655 155.990 86.825 ;
        RECT 155.820 86.295 155.990 86.465 ;
        RECT 155.820 81.905 155.990 82.075 ;
        RECT 155.820 81.545 155.990 81.715 ;
        RECT 155.820 81.185 155.990 81.355 ;
        RECT 155.820 80.825 155.990 80.995 ;
        RECT 155.820 76.435 155.990 76.605 ;
        RECT 166.400 97.595 166.570 97.765 ;
        RECT 166.400 97.235 166.570 97.405 ;
        RECT 166.400 92.845 166.570 93.015 ;
        RECT 166.400 92.485 166.570 92.655 ;
        RECT 166.400 92.125 166.570 92.295 ;
        RECT 166.400 91.765 166.570 91.935 ;
        RECT 166.400 87.375 166.570 87.545 ;
        RECT 166.400 87.015 166.570 87.185 ;
        RECT 166.400 86.655 166.570 86.825 ;
        RECT 166.400 86.295 166.570 86.465 ;
        RECT 166.400 81.905 166.570 82.075 ;
        RECT 166.400 81.545 166.570 81.715 ;
        RECT 166.400 81.185 166.570 81.355 ;
        RECT 166.400 80.825 166.570 80.995 ;
        RECT 166.400 76.435 166.570 76.605 ;
        RECT 177.790 97.625 177.960 97.795 ;
        RECT 177.790 97.265 177.960 97.435 ;
        RECT 177.790 92.875 177.960 93.045 ;
        RECT 177.790 92.515 177.960 92.685 ;
        RECT 177.790 92.155 177.960 92.325 ;
        RECT 177.790 91.795 177.960 91.965 ;
        RECT 177.790 87.405 177.960 87.575 ;
        RECT 177.790 87.045 177.960 87.215 ;
        RECT 177.790 86.685 177.960 86.855 ;
        RECT 177.790 86.325 177.960 86.495 ;
        RECT 177.790 81.935 177.960 82.105 ;
        RECT 177.790 81.575 177.960 81.745 ;
        RECT 177.790 81.215 177.960 81.385 ;
        RECT 177.790 80.855 177.960 81.025 ;
        RECT 177.790 76.465 177.960 76.635 ;
        RECT 133.790 75.995 133.960 76.165 ;
        RECT 133.790 75.635 133.960 75.805 ;
        RECT 145.240 76.075 145.410 76.245 ;
        RECT 112.630 75.275 112.800 75.445 ;
        RECT 123.210 75.275 123.380 75.445 ;
        RECT 133.790 75.275 133.960 75.445 ;
        RECT 145.240 75.715 145.410 75.885 ;
        RECT 155.820 76.075 155.990 76.245 ;
        RECT 155.820 75.715 155.990 75.885 ;
        RECT 188.370 97.985 188.540 98.155 ;
        RECT 198.950 97.985 199.120 98.155 ;
        RECT 376.370 98.235 376.540 98.405 ;
        RECT 386.950 98.235 387.120 98.405 ;
        RECT 397.530 98.235 397.700 98.405 ;
        RECT 376.370 97.875 376.540 98.045 ;
        RECT 408.690 98.295 408.860 98.465 ;
        RECT 419.270 98.295 419.440 98.465 ;
        RECT 429.850 98.295 430.020 98.465 ;
        RECT 188.370 97.625 188.540 97.795 ;
        RECT 188.370 97.265 188.540 97.435 ;
        RECT 188.370 92.875 188.540 93.045 ;
        RECT 188.370 92.515 188.540 92.685 ;
        RECT 188.370 92.155 188.540 92.325 ;
        RECT 188.370 91.795 188.540 91.965 ;
        RECT 188.370 87.405 188.540 87.575 ;
        RECT 188.370 87.045 188.540 87.215 ;
        RECT 188.370 86.685 188.540 86.855 ;
        RECT 188.370 86.325 188.540 86.495 ;
        RECT 188.370 81.935 188.540 82.105 ;
        RECT 188.370 81.575 188.540 81.745 ;
        RECT 188.370 81.215 188.540 81.385 ;
        RECT 188.370 80.855 188.540 81.025 ;
        RECT 188.370 76.465 188.540 76.635 ;
        RECT 198.950 97.625 199.120 97.795 ;
        RECT 198.950 97.265 199.120 97.435 ;
        RECT 198.950 92.875 199.120 93.045 ;
        RECT 198.950 92.515 199.120 92.685 ;
        RECT 198.950 92.155 199.120 92.325 ;
        RECT 198.950 91.795 199.120 91.965 ;
        RECT 198.950 87.405 199.120 87.575 ;
        RECT 198.950 87.045 199.120 87.215 ;
        RECT 198.950 86.685 199.120 86.855 ;
        RECT 198.950 86.325 199.120 86.495 ;
        RECT 198.950 81.935 199.120 82.105 ;
        RECT 198.950 81.575 199.120 81.745 ;
        RECT 198.950 81.215 199.120 81.385 ;
        RECT 198.950 80.855 199.120 81.025 ;
        RECT 198.950 76.465 199.120 76.635 ;
        RECT 376.370 97.515 376.540 97.685 ;
        RECT 376.370 97.155 376.540 97.325 ;
        RECT 386.950 97.875 387.120 98.045 ;
        RECT 386.950 97.515 387.120 97.685 ;
        RECT 386.950 97.155 387.120 97.325 ;
        RECT 376.370 92.765 376.540 92.935 ;
        RECT 376.370 92.405 376.540 92.575 ;
        RECT 376.370 92.045 376.540 92.215 ;
        RECT 376.370 91.685 376.540 91.855 ;
        RECT 386.950 92.765 387.120 92.935 ;
        RECT 386.950 92.405 387.120 92.575 ;
        RECT 386.950 92.045 387.120 92.215 ;
        RECT 386.950 91.685 387.120 91.855 ;
        RECT 376.370 87.295 376.540 87.465 ;
        RECT 376.370 86.935 376.540 87.105 ;
        RECT 376.370 86.575 376.540 86.745 ;
        RECT 376.370 86.215 376.540 86.385 ;
        RECT 386.950 87.295 387.120 87.465 ;
        RECT 386.950 86.935 387.120 87.105 ;
        RECT 386.950 86.575 387.120 86.745 ;
        RECT 386.950 86.215 387.120 86.385 ;
        RECT 376.370 81.825 376.540 81.995 ;
        RECT 376.370 81.465 376.540 81.635 ;
        RECT 376.370 81.105 376.540 81.275 ;
        RECT 376.370 80.745 376.540 80.915 ;
        RECT 386.950 81.825 387.120 81.995 ;
        RECT 386.950 81.465 387.120 81.635 ;
        RECT 386.950 81.105 387.120 81.275 ;
        RECT 386.950 80.745 387.120 80.915 ;
        RECT 166.400 76.075 166.570 76.245 ;
        RECT 166.400 75.715 166.570 75.885 ;
        RECT 177.790 76.105 177.960 76.275 ;
        RECT 177.790 75.745 177.960 75.915 ;
        RECT 188.370 76.105 188.540 76.275 ;
        RECT 145.240 75.355 145.410 75.525 ;
        RECT 155.820 75.355 155.990 75.525 ;
        RECT 166.400 75.355 166.570 75.525 ;
        RECT 188.370 75.745 188.540 75.915 ;
        RECT 376.370 76.355 376.540 76.525 ;
        RECT 386.950 76.355 387.120 76.525 ;
        RECT 397.530 97.875 397.700 98.045 ;
        RECT 397.530 97.515 397.700 97.685 ;
        RECT 397.530 97.155 397.700 97.325 ;
        RECT 397.530 92.765 397.700 92.935 ;
        RECT 397.530 92.405 397.700 92.575 ;
        RECT 397.530 92.045 397.700 92.215 ;
        RECT 397.530 91.685 397.700 91.855 ;
        RECT 397.530 87.295 397.700 87.465 ;
        RECT 397.530 86.935 397.700 87.105 ;
        RECT 397.530 86.575 397.700 86.745 ;
        RECT 397.530 86.215 397.700 86.385 ;
        RECT 397.530 81.825 397.700 81.995 ;
        RECT 397.530 81.465 397.700 81.635 ;
        RECT 397.530 81.105 397.700 81.275 ;
        RECT 397.530 80.745 397.700 80.915 ;
        RECT 397.530 76.355 397.700 76.525 ;
        RECT 408.690 97.935 408.860 98.105 ;
        RECT 408.690 97.575 408.860 97.745 ;
        RECT 408.690 97.215 408.860 97.385 ;
        RECT 419.270 97.935 419.440 98.105 ;
        RECT 419.270 97.575 419.440 97.745 ;
        RECT 419.270 97.215 419.440 97.385 ;
        RECT 408.690 92.825 408.860 92.995 ;
        RECT 408.690 92.465 408.860 92.635 ;
        RECT 408.690 92.105 408.860 92.275 ;
        RECT 408.690 91.745 408.860 91.915 ;
        RECT 419.270 92.825 419.440 92.995 ;
        RECT 419.270 92.465 419.440 92.635 ;
        RECT 419.270 92.105 419.440 92.275 ;
        RECT 419.270 91.745 419.440 91.915 ;
        RECT 408.690 87.355 408.860 87.525 ;
        RECT 408.690 86.995 408.860 87.165 ;
        RECT 408.690 86.635 408.860 86.805 ;
        RECT 408.690 86.275 408.860 86.445 ;
        RECT 419.270 87.355 419.440 87.525 ;
        RECT 419.270 86.995 419.440 87.165 ;
        RECT 419.270 86.635 419.440 86.805 ;
        RECT 419.270 86.275 419.440 86.445 ;
        RECT 408.690 81.885 408.860 82.055 ;
        RECT 408.690 81.525 408.860 81.695 ;
        RECT 408.690 81.165 408.860 81.335 ;
        RECT 408.690 80.805 408.860 80.975 ;
        RECT 419.270 81.885 419.440 82.055 ;
        RECT 419.270 81.525 419.440 81.695 ;
        RECT 419.270 81.165 419.440 81.335 ;
        RECT 419.270 80.805 419.440 80.975 ;
        RECT 408.690 76.415 408.860 76.585 ;
        RECT 419.270 76.415 419.440 76.585 ;
        RECT 429.850 97.935 430.020 98.105 ;
        RECT 429.850 97.575 430.020 97.745 ;
        RECT 429.850 97.215 430.020 97.385 ;
        RECT 429.850 92.825 430.020 92.995 ;
        RECT 429.850 92.465 430.020 92.635 ;
        RECT 429.850 92.105 430.020 92.275 ;
        RECT 429.850 91.745 430.020 91.915 ;
        RECT 429.850 87.355 430.020 87.525 ;
        RECT 429.850 86.995 430.020 87.165 ;
        RECT 429.850 86.635 430.020 86.805 ;
        RECT 429.850 86.275 430.020 86.445 ;
        RECT 429.850 81.885 430.020 82.055 ;
        RECT 429.850 81.525 430.020 81.695 ;
        RECT 429.850 81.165 430.020 81.335 ;
        RECT 429.850 80.805 430.020 80.975 ;
        RECT 429.850 76.415 430.020 76.585 ;
        RECT 198.950 76.105 199.120 76.275 ;
        RECT 198.950 75.745 199.120 75.915 ;
        RECT 376.370 75.995 376.540 76.165 ;
        RECT 177.790 75.385 177.960 75.555 ;
        RECT 188.370 75.385 188.540 75.555 ;
        RECT 198.950 75.385 199.120 75.555 ;
        RECT 376.370 75.635 376.540 75.805 ;
        RECT 376.370 75.275 376.540 75.445 ;
        RECT 386.950 75.995 387.120 76.165 ;
        RECT 386.950 75.635 387.120 75.805 ;
        RECT 386.950 75.275 387.120 75.445 ;
        RECT 397.530 75.995 397.700 76.165 ;
        RECT 397.530 75.635 397.700 75.805 ;
        RECT 397.530 75.275 397.700 75.445 ;
        RECT 408.690 76.055 408.860 76.225 ;
        RECT 408.690 75.695 408.860 75.865 ;
        RECT 408.690 75.335 408.860 75.505 ;
        RECT 419.270 76.055 419.440 76.225 ;
        RECT 419.270 75.695 419.440 75.865 ;
        RECT 419.270 75.335 419.440 75.505 ;
        RECT 429.850 76.055 430.020 76.225 ;
        RECT 429.850 75.695 430.020 75.865 ;
        RECT 429.850 75.335 430.020 75.505 ;
        RECT 112.680 68.955 112.850 69.125 ;
        RECT 112.680 68.595 112.850 68.765 ;
        RECT 123.260 68.955 123.430 69.125 ;
        RECT 133.840 68.955 134.010 69.125 ;
        RECT 112.680 68.235 112.850 68.405 ;
        RECT 112.680 67.875 112.850 68.045 ;
        RECT 112.680 63.485 112.850 63.655 ;
        RECT 112.680 63.125 112.850 63.295 ;
        RECT 112.680 62.765 112.850 62.935 ;
        RECT 112.680 62.405 112.850 62.575 ;
        RECT 112.680 58.015 112.850 58.185 ;
        RECT 112.680 57.655 112.850 57.825 ;
        RECT 112.680 57.295 112.850 57.465 ;
        RECT 112.680 56.935 112.850 57.105 ;
        RECT 112.680 52.545 112.850 52.715 ;
        RECT 112.680 52.185 112.850 52.355 ;
        RECT 112.680 51.825 112.850 51.995 ;
        RECT 112.680 51.465 112.850 51.635 ;
        RECT 112.680 47.075 112.850 47.245 ;
        RECT 123.260 68.595 123.430 68.765 ;
        RECT 145.290 69.035 145.460 69.205 ;
        RECT 123.260 68.235 123.430 68.405 ;
        RECT 123.260 67.875 123.430 68.045 ;
        RECT 123.260 63.485 123.430 63.655 ;
        RECT 123.260 63.125 123.430 63.295 ;
        RECT 123.260 62.765 123.430 62.935 ;
        RECT 123.260 62.405 123.430 62.575 ;
        RECT 123.260 58.015 123.430 58.185 ;
        RECT 123.260 57.655 123.430 57.825 ;
        RECT 123.260 57.295 123.430 57.465 ;
        RECT 123.260 56.935 123.430 57.105 ;
        RECT 123.260 52.545 123.430 52.715 ;
        RECT 123.260 52.185 123.430 52.355 ;
        RECT 123.260 51.825 123.430 51.995 ;
        RECT 123.260 51.465 123.430 51.635 ;
        RECT 123.260 47.075 123.430 47.245 ;
        RECT 133.840 68.595 134.010 68.765 ;
        RECT 133.840 68.235 134.010 68.405 ;
        RECT 133.840 67.875 134.010 68.045 ;
        RECT 133.840 63.485 134.010 63.655 ;
        RECT 133.840 63.125 134.010 63.295 ;
        RECT 133.840 62.765 134.010 62.935 ;
        RECT 133.840 62.405 134.010 62.575 ;
        RECT 133.840 58.015 134.010 58.185 ;
        RECT 133.840 57.655 134.010 57.825 ;
        RECT 133.840 57.295 134.010 57.465 ;
        RECT 133.840 56.935 134.010 57.105 ;
        RECT 133.840 52.545 134.010 52.715 ;
        RECT 133.840 52.185 134.010 52.355 ;
        RECT 133.840 51.825 134.010 51.995 ;
        RECT 133.840 51.465 134.010 51.635 ;
        RECT 133.840 47.075 134.010 47.245 ;
        RECT 145.290 68.675 145.460 68.845 ;
        RECT 155.870 69.035 156.040 69.205 ;
        RECT 166.450 69.035 166.620 69.205 ;
        RECT 145.290 68.315 145.460 68.485 ;
        RECT 145.290 67.955 145.460 68.125 ;
        RECT 145.290 63.565 145.460 63.735 ;
        RECT 145.290 63.205 145.460 63.375 ;
        RECT 145.290 62.845 145.460 63.015 ;
        RECT 145.290 62.485 145.460 62.655 ;
        RECT 145.290 58.095 145.460 58.265 ;
        RECT 145.290 57.735 145.460 57.905 ;
        RECT 145.290 57.375 145.460 57.545 ;
        RECT 145.290 57.015 145.460 57.185 ;
        RECT 145.290 52.625 145.460 52.795 ;
        RECT 145.290 52.265 145.460 52.435 ;
        RECT 145.290 51.905 145.460 52.075 ;
        RECT 145.290 51.545 145.460 51.715 ;
        RECT 145.290 47.155 145.460 47.325 ;
        RECT 112.680 46.715 112.850 46.885 ;
        RECT 112.680 46.355 112.850 46.525 ;
        RECT 123.260 46.715 123.430 46.885 ;
        RECT 123.260 46.355 123.430 46.525 ;
        RECT 155.870 68.675 156.040 68.845 ;
        RECT 155.870 68.315 156.040 68.485 ;
        RECT 177.840 69.065 178.010 69.235 ;
        RECT 166.450 68.675 166.620 68.845 ;
        RECT 166.450 68.315 166.620 68.485 ;
        RECT 177.840 68.705 178.010 68.875 ;
        RECT 188.420 69.065 188.590 69.235 ;
        RECT 199.000 69.065 199.170 69.235 ;
        RECT 177.840 68.345 178.010 68.515 ;
        RECT 155.870 67.955 156.040 68.125 ;
        RECT 155.870 63.565 156.040 63.735 ;
        RECT 155.870 63.205 156.040 63.375 ;
        RECT 155.870 62.845 156.040 63.015 ;
        RECT 155.870 62.485 156.040 62.655 ;
        RECT 155.870 58.095 156.040 58.265 ;
        RECT 155.870 57.735 156.040 57.905 ;
        RECT 155.870 57.375 156.040 57.545 ;
        RECT 155.870 57.015 156.040 57.185 ;
        RECT 155.870 52.625 156.040 52.795 ;
        RECT 155.870 52.265 156.040 52.435 ;
        RECT 155.870 51.905 156.040 52.075 ;
        RECT 155.870 51.545 156.040 51.715 ;
        RECT 155.870 47.155 156.040 47.325 ;
        RECT 166.450 67.955 166.620 68.125 ;
        RECT 166.450 63.565 166.620 63.735 ;
        RECT 166.450 63.205 166.620 63.375 ;
        RECT 166.450 62.845 166.620 63.015 ;
        RECT 166.450 62.485 166.620 62.655 ;
        RECT 166.450 58.095 166.620 58.265 ;
        RECT 166.450 57.735 166.620 57.905 ;
        RECT 166.450 57.375 166.620 57.545 ;
        RECT 166.450 57.015 166.620 57.185 ;
        RECT 166.450 52.625 166.620 52.795 ;
        RECT 166.450 52.265 166.620 52.435 ;
        RECT 166.450 51.905 166.620 52.075 ;
        RECT 166.450 51.545 166.620 51.715 ;
        RECT 166.450 47.155 166.620 47.325 ;
        RECT 177.840 67.985 178.010 68.155 ;
        RECT 177.840 63.595 178.010 63.765 ;
        RECT 177.840 63.235 178.010 63.405 ;
        RECT 177.840 62.875 178.010 63.045 ;
        RECT 177.840 62.515 178.010 62.685 ;
        RECT 177.840 58.125 178.010 58.295 ;
        RECT 177.840 57.765 178.010 57.935 ;
        RECT 177.840 57.405 178.010 57.575 ;
        RECT 177.840 57.045 178.010 57.215 ;
        RECT 177.840 52.655 178.010 52.825 ;
        RECT 177.840 52.295 178.010 52.465 ;
        RECT 177.840 51.935 178.010 52.105 ;
        RECT 177.840 51.575 178.010 51.745 ;
        RECT 177.840 47.185 178.010 47.355 ;
        RECT 133.840 46.715 134.010 46.885 ;
        RECT 133.840 46.355 134.010 46.525 ;
        RECT 145.290 46.795 145.460 46.965 ;
        RECT 145.290 46.435 145.460 46.605 ;
        RECT 155.870 46.795 156.040 46.965 ;
        RECT 112.680 45.995 112.850 46.165 ;
        RECT 123.260 45.995 123.430 46.165 ;
        RECT 133.840 45.995 134.010 46.165 ;
        RECT 155.870 46.435 156.040 46.605 ;
        RECT 188.420 68.705 188.590 68.875 ;
        RECT 188.420 68.345 188.590 68.515 ;
        RECT 199.000 68.705 199.170 68.875 ;
        RECT 188.420 67.985 188.590 68.155 ;
        RECT 188.420 63.595 188.590 63.765 ;
        RECT 188.420 63.235 188.590 63.405 ;
        RECT 188.420 62.875 188.590 63.045 ;
        RECT 188.420 62.515 188.590 62.685 ;
        RECT 188.420 58.125 188.590 58.295 ;
        RECT 188.420 57.765 188.590 57.935 ;
        RECT 188.420 57.405 188.590 57.575 ;
        RECT 188.420 57.045 188.590 57.215 ;
        RECT 188.420 52.655 188.590 52.825 ;
        RECT 188.420 52.295 188.590 52.465 ;
        RECT 188.420 51.935 188.590 52.105 ;
        RECT 188.420 51.575 188.590 51.745 ;
        RECT 188.420 47.185 188.590 47.355 ;
        RECT 199.000 68.345 199.170 68.515 ;
        RECT 376.370 68.945 376.540 69.115 ;
        RECT 386.950 68.945 387.120 69.115 ;
        RECT 397.530 68.945 397.700 69.115 ;
        RECT 376.370 68.585 376.540 68.755 ;
        RECT 408.710 68.935 408.880 69.105 ;
        RECT 199.000 67.985 199.170 68.155 ;
        RECT 199.000 63.595 199.170 63.765 ;
        RECT 199.000 63.235 199.170 63.405 ;
        RECT 199.000 62.875 199.170 63.045 ;
        RECT 199.000 62.515 199.170 62.685 ;
        RECT 199.000 58.125 199.170 58.295 ;
        RECT 199.000 57.765 199.170 57.935 ;
        RECT 199.000 57.405 199.170 57.575 ;
        RECT 199.000 57.045 199.170 57.215 ;
        RECT 199.000 52.655 199.170 52.825 ;
        RECT 199.000 52.295 199.170 52.465 ;
        RECT 199.000 51.935 199.170 52.105 ;
        RECT 199.000 51.575 199.170 51.745 ;
        RECT 199.000 47.185 199.170 47.355 ;
        RECT 376.370 68.225 376.540 68.395 ;
        RECT 376.370 67.865 376.540 68.035 ;
        RECT 386.950 68.585 387.120 68.755 ;
        RECT 386.950 68.225 387.120 68.395 ;
        RECT 386.950 67.865 387.120 68.035 ;
        RECT 376.370 63.475 376.540 63.645 ;
        RECT 376.370 63.115 376.540 63.285 ;
        RECT 376.370 62.755 376.540 62.925 ;
        RECT 376.370 62.395 376.540 62.565 ;
        RECT 386.950 63.475 387.120 63.645 ;
        RECT 386.950 63.115 387.120 63.285 ;
        RECT 386.950 62.755 387.120 62.925 ;
        RECT 386.950 62.395 387.120 62.565 ;
        RECT 376.370 58.005 376.540 58.175 ;
        RECT 376.370 57.645 376.540 57.815 ;
        RECT 376.370 57.285 376.540 57.455 ;
        RECT 376.370 56.925 376.540 57.095 ;
        RECT 386.950 58.005 387.120 58.175 ;
        RECT 386.950 57.645 387.120 57.815 ;
        RECT 386.950 57.285 387.120 57.455 ;
        RECT 386.950 56.925 387.120 57.095 ;
        RECT 376.370 52.535 376.540 52.705 ;
        RECT 376.370 52.175 376.540 52.345 ;
        RECT 376.370 51.815 376.540 51.985 ;
        RECT 376.370 51.455 376.540 51.625 ;
        RECT 386.950 52.535 387.120 52.705 ;
        RECT 386.950 52.175 387.120 52.345 ;
        RECT 386.950 51.815 387.120 51.985 ;
        RECT 386.950 51.455 387.120 51.625 ;
        RECT 166.450 46.795 166.620 46.965 ;
        RECT 166.450 46.435 166.620 46.605 ;
        RECT 177.840 46.825 178.010 46.995 ;
        RECT 177.840 46.465 178.010 46.635 ;
        RECT 188.420 46.825 188.590 46.995 ;
        RECT 145.290 46.075 145.460 46.245 ;
        RECT 155.870 46.075 156.040 46.245 ;
        RECT 166.450 46.075 166.620 46.245 ;
        RECT 188.420 46.465 188.590 46.635 ;
        RECT 376.370 47.065 376.540 47.235 ;
        RECT 386.950 47.065 387.120 47.235 ;
        RECT 397.530 68.585 397.700 68.755 ;
        RECT 397.530 68.225 397.700 68.395 ;
        RECT 397.530 67.865 397.700 68.035 ;
        RECT 397.530 63.475 397.700 63.645 ;
        RECT 397.530 63.115 397.700 63.285 ;
        RECT 397.530 62.755 397.700 62.925 ;
        RECT 397.530 62.395 397.700 62.565 ;
        RECT 397.530 58.005 397.700 58.175 ;
        RECT 397.530 57.645 397.700 57.815 ;
        RECT 397.530 57.285 397.700 57.455 ;
        RECT 397.530 56.925 397.700 57.095 ;
        RECT 397.530 52.535 397.700 52.705 ;
        RECT 397.530 52.175 397.700 52.345 ;
        RECT 397.530 51.815 397.700 51.985 ;
        RECT 397.530 51.455 397.700 51.625 ;
        RECT 397.530 47.065 397.700 47.235 ;
        RECT 419.290 68.935 419.460 69.105 ;
        RECT 429.870 68.935 430.040 69.105 ;
        RECT 408.710 68.575 408.880 68.745 ;
        RECT 408.710 68.215 408.880 68.385 ;
        RECT 408.710 67.855 408.880 68.025 ;
        RECT 419.290 68.575 419.460 68.745 ;
        RECT 419.290 68.215 419.460 68.385 ;
        RECT 419.290 67.855 419.460 68.025 ;
        RECT 408.710 63.465 408.880 63.635 ;
        RECT 408.710 63.105 408.880 63.275 ;
        RECT 408.710 62.745 408.880 62.915 ;
        RECT 408.710 62.385 408.880 62.555 ;
        RECT 419.290 63.465 419.460 63.635 ;
        RECT 419.290 63.105 419.460 63.275 ;
        RECT 419.290 62.745 419.460 62.915 ;
        RECT 419.290 62.385 419.460 62.555 ;
        RECT 408.710 57.995 408.880 58.165 ;
        RECT 408.710 57.635 408.880 57.805 ;
        RECT 408.710 57.275 408.880 57.445 ;
        RECT 408.710 56.915 408.880 57.085 ;
        RECT 419.290 57.995 419.460 58.165 ;
        RECT 419.290 57.635 419.460 57.805 ;
        RECT 419.290 57.275 419.460 57.445 ;
        RECT 419.290 56.915 419.460 57.085 ;
        RECT 408.710 52.525 408.880 52.695 ;
        RECT 408.710 52.165 408.880 52.335 ;
        RECT 408.710 51.805 408.880 51.975 ;
        RECT 408.710 51.445 408.880 51.615 ;
        RECT 419.290 52.525 419.460 52.695 ;
        RECT 419.290 52.165 419.460 52.335 ;
        RECT 419.290 51.805 419.460 51.975 ;
        RECT 419.290 51.445 419.460 51.615 ;
        RECT 199.000 46.825 199.170 46.995 ;
        RECT 199.000 46.465 199.170 46.635 ;
        RECT 376.370 46.705 376.540 46.875 ;
        RECT 177.840 46.105 178.010 46.275 ;
        RECT 188.420 46.105 188.590 46.275 ;
        RECT 376.370 46.345 376.540 46.515 ;
        RECT 199.000 46.105 199.170 46.275 ;
        RECT 376.370 45.985 376.540 46.155 ;
        RECT 386.950 46.705 387.120 46.875 ;
        RECT 386.950 46.345 387.120 46.515 ;
        RECT 386.950 45.985 387.120 46.155 ;
        RECT 408.710 47.055 408.880 47.225 ;
        RECT 419.290 47.055 419.460 47.225 ;
        RECT 429.870 68.575 430.040 68.745 ;
        RECT 429.870 68.215 430.040 68.385 ;
        RECT 429.870 67.855 430.040 68.025 ;
        RECT 429.870 63.465 430.040 63.635 ;
        RECT 429.870 63.105 430.040 63.275 ;
        RECT 429.870 62.745 430.040 62.915 ;
        RECT 429.870 62.385 430.040 62.555 ;
        RECT 429.870 57.995 430.040 58.165 ;
        RECT 429.870 57.635 430.040 57.805 ;
        RECT 429.870 57.275 430.040 57.445 ;
        RECT 429.870 56.915 430.040 57.085 ;
        RECT 429.870 52.525 430.040 52.695 ;
        RECT 429.870 52.165 430.040 52.335 ;
        RECT 429.870 51.805 430.040 51.975 ;
        RECT 429.870 51.445 430.040 51.615 ;
        RECT 429.870 47.055 430.040 47.225 ;
        RECT 397.530 46.705 397.700 46.875 ;
        RECT 397.530 46.345 397.700 46.515 ;
        RECT 397.530 45.985 397.700 46.155 ;
        RECT 408.710 46.695 408.880 46.865 ;
        RECT 408.710 46.335 408.880 46.505 ;
        RECT 408.710 45.975 408.880 46.145 ;
        RECT 419.290 46.695 419.460 46.865 ;
        RECT 419.290 46.335 419.460 46.505 ;
        RECT 419.290 45.975 419.460 46.145 ;
        RECT 429.870 46.695 430.040 46.865 ;
        RECT 429.870 46.335 430.040 46.505 ;
        RECT 429.870 45.975 430.040 46.145 ;
        RECT 112.770 39.415 112.940 39.585 ;
        RECT 112.770 39.055 112.940 39.225 ;
        RECT 123.350 39.415 123.520 39.585 ;
        RECT 133.930 39.415 134.100 39.585 ;
        RECT 112.770 38.695 112.940 38.865 ;
        RECT 112.770 38.335 112.940 38.505 ;
        RECT 112.770 33.945 112.940 34.115 ;
        RECT 112.770 33.585 112.940 33.755 ;
        RECT 112.770 33.225 112.940 33.395 ;
        RECT 112.770 32.865 112.940 33.035 ;
        RECT 112.770 28.475 112.940 28.645 ;
        RECT 112.770 28.115 112.940 28.285 ;
        RECT 112.770 27.755 112.940 27.925 ;
        RECT 112.770 27.395 112.940 27.565 ;
        RECT 112.770 23.005 112.940 23.175 ;
        RECT 112.770 22.645 112.940 22.815 ;
        RECT 112.770 22.285 112.940 22.455 ;
        RECT 112.770 21.925 112.940 22.095 ;
        RECT 112.770 17.535 112.940 17.705 ;
        RECT 123.350 39.055 123.520 39.225 ;
        RECT 145.380 39.495 145.550 39.665 ;
        RECT 133.930 39.055 134.100 39.225 ;
        RECT 145.380 39.135 145.550 39.305 ;
        RECT 155.960 39.495 156.130 39.665 ;
        RECT 166.540 39.495 166.710 39.665 ;
        RECT 123.350 38.695 123.520 38.865 ;
        RECT 123.350 38.335 123.520 38.505 ;
        RECT 123.350 33.945 123.520 34.115 ;
        RECT 123.350 33.585 123.520 33.755 ;
        RECT 123.350 33.225 123.520 33.395 ;
        RECT 123.350 32.865 123.520 33.035 ;
        RECT 123.350 28.475 123.520 28.645 ;
        RECT 123.350 28.115 123.520 28.285 ;
        RECT 123.350 27.755 123.520 27.925 ;
        RECT 123.350 27.395 123.520 27.565 ;
        RECT 123.350 23.005 123.520 23.175 ;
        RECT 123.350 22.645 123.520 22.815 ;
        RECT 123.350 22.285 123.520 22.455 ;
        RECT 123.350 21.925 123.520 22.095 ;
        RECT 123.350 17.535 123.520 17.705 ;
        RECT 133.930 38.695 134.100 38.865 ;
        RECT 133.930 38.335 134.100 38.505 ;
        RECT 133.930 33.945 134.100 34.115 ;
        RECT 133.930 33.585 134.100 33.755 ;
        RECT 133.930 33.225 134.100 33.395 ;
        RECT 133.930 32.865 134.100 33.035 ;
        RECT 133.930 28.475 134.100 28.645 ;
        RECT 133.930 28.115 134.100 28.285 ;
        RECT 133.930 27.755 134.100 27.925 ;
        RECT 133.930 27.395 134.100 27.565 ;
        RECT 133.930 23.005 134.100 23.175 ;
        RECT 133.930 22.645 134.100 22.815 ;
        RECT 133.930 22.285 134.100 22.455 ;
        RECT 133.930 21.925 134.100 22.095 ;
        RECT 133.930 17.535 134.100 17.705 ;
        RECT 145.380 38.775 145.550 38.945 ;
        RECT 145.380 38.415 145.550 38.585 ;
        RECT 145.380 34.025 145.550 34.195 ;
        RECT 145.380 33.665 145.550 33.835 ;
        RECT 145.380 33.305 145.550 33.475 ;
        RECT 145.380 32.945 145.550 33.115 ;
        RECT 145.380 28.555 145.550 28.725 ;
        RECT 145.380 28.195 145.550 28.365 ;
        RECT 145.380 27.835 145.550 28.005 ;
        RECT 145.380 27.475 145.550 27.645 ;
        RECT 145.380 23.085 145.550 23.255 ;
        RECT 145.380 22.725 145.550 22.895 ;
        RECT 145.380 22.365 145.550 22.535 ;
        RECT 145.380 22.005 145.550 22.175 ;
        RECT 145.380 17.615 145.550 17.785 ;
        RECT 112.770 17.175 112.940 17.345 ;
        RECT 112.770 16.815 112.940 16.985 ;
        RECT 123.350 17.175 123.520 17.345 ;
        RECT 123.350 16.815 123.520 16.985 ;
        RECT 155.960 39.135 156.130 39.305 ;
        RECT 177.930 39.525 178.100 39.695 ;
        RECT 166.540 39.135 166.710 39.305 ;
        RECT 177.930 39.165 178.100 39.335 ;
        RECT 188.510 39.525 188.680 39.695 ;
        RECT 199.090 39.525 199.260 39.695 ;
        RECT 376.370 39.655 376.540 39.825 ;
        RECT 386.950 39.655 387.120 39.825 ;
        RECT 397.530 39.655 397.700 39.825 ;
        RECT 155.960 38.775 156.130 38.945 ;
        RECT 155.960 38.415 156.130 38.585 ;
        RECT 155.960 34.025 156.130 34.195 ;
        RECT 155.960 33.665 156.130 33.835 ;
        RECT 155.960 33.305 156.130 33.475 ;
        RECT 155.960 32.945 156.130 33.115 ;
        RECT 155.960 28.555 156.130 28.725 ;
        RECT 155.960 28.195 156.130 28.365 ;
        RECT 155.960 27.835 156.130 28.005 ;
        RECT 155.960 27.475 156.130 27.645 ;
        RECT 155.960 23.085 156.130 23.255 ;
        RECT 155.960 22.725 156.130 22.895 ;
        RECT 155.960 22.365 156.130 22.535 ;
        RECT 155.960 22.005 156.130 22.175 ;
        RECT 155.960 17.615 156.130 17.785 ;
        RECT 166.540 38.775 166.710 38.945 ;
        RECT 166.540 38.415 166.710 38.585 ;
        RECT 166.540 34.025 166.710 34.195 ;
        RECT 166.540 33.665 166.710 33.835 ;
        RECT 166.540 33.305 166.710 33.475 ;
        RECT 166.540 32.945 166.710 33.115 ;
        RECT 166.540 28.555 166.710 28.725 ;
        RECT 166.540 28.195 166.710 28.365 ;
        RECT 166.540 27.835 166.710 28.005 ;
        RECT 166.540 27.475 166.710 27.645 ;
        RECT 166.540 23.085 166.710 23.255 ;
        RECT 166.540 22.725 166.710 22.895 ;
        RECT 166.540 22.365 166.710 22.535 ;
        RECT 166.540 22.005 166.710 22.175 ;
        RECT 166.540 17.615 166.710 17.785 ;
        RECT 177.930 38.805 178.100 38.975 ;
        RECT 177.930 38.445 178.100 38.615 ;
        RECT 177.930 34.055 178.100 34.225 ;
        RECT 177.930 33.695 178.100 33.865 ;
        RECT 177.930 33.335 178.100 33.505 ;
        RECT 177.930 32.975 178.100 33.145 ;
        RECT 177.930 28.585 178.100 28.755 ;
        RECT 177.930 28.225 178.100 28.395 ;
        RECT 177.930 27.865 178.100 28.035 ;
        RECT 177.930 27.505 178.100 27.675 ;
        RECT 177.930 23.115 178.100 23.285 ;
        RECT 177.930 22.755 178.100 22.925 ;
        RECT 177.930 22.395 178.100 22.565 ;
        RECT 177.930 22.035 178.100 22.205 ;
        RECT 177.930 17.645 178.100 17.815 ;
        RECT 133.930 17.175 134.100 17.345 ;
        RECT 133.930 16.815 134.100 16.985 ;
        RECT 145.380 17.255 145.550 17.425 ;
        RECT 145.380 16.895 145.550 17.065 ;
        RECT 155.960 17.255 156.130 17.425 ;
        RECT 112.770 16.455 112.940 16.625 ;
        RECT 123.350 16.455 123.520 16.625 ;
        RECT 133.930 16.455 134.100 16.625 ;
        RECT 155.960 16.895 156.130 17.065 ;
        RECT 188.510 39.165 188.680 39.335 ;
        RECT 188.510 38.805 188.680 38.975 ;
        RECT 188.510 38.445 188.680 38.615 ;
        RECT 188.510 34.055 188.680 34.225 ;
        RECT 188.510 33.695 188.680 33.865 ;
        RECT 188.510 33.335 188.680 33.505 ;
        RECT 188.510 32.975 188.680 33.145 ;
        RECT 188.510 28.585 188.680 28.755 ;
        RECT 188.510 28.225 188.680 28.395 ;
        RECT 188.510 27.865 188.680 28.035 ;
        RECT 188.510 27.505 188.680 27.675 ;
        RECT 188.510 23.115 188.680 23.285 ;
        RECT 188.510 22.755 188.680 22.925 ;
        RECT 188.510 22.395 188.680 22.565 ;
        RECT 188.510 22.035 188.680 22.205 ;
        RECT 188.510 17.645 188.680 17.815 ;
        RECT 199.090 39.165 199.260 39.335 ;
        RECT 199.090 38.805 199.260 38.975 ;
        RECT 199.090 38.445 199.260 38.615 ;
        RECT 199.090 34.055 199.260 34.225 ;
        RECT 199.090 33.695 199.260 33.865 ;
        RECT 199.090 33.335 199.260 33.505 ;
        RECT 199.090 32.975 199.260 33.145 ;
        RECT 199.090 28.585 199.260 28.755 ;
        RECT 199.090 28.225 199.260 28.395 ;
        RECT 199.090 27.865 199.260 28.035 ;
        RECT 199.090 27.505 199.260 27.675 ;
        RECT 199.090 23.115 199.260 23.285 ;
        RECT 199.090 22.755 199.260 22.925 ;
        RECT 199.090 22.395 199.260 22.565 ;
        RECT 199.090 22.035 199.260 22.205 ;
        RECT 199.090 17.645 199.260 17.815 ;
        RECT 376.370 39.295 376.540 39.465 ;
        RECT 408.730 39.645 408.900 39.815 ;
        RECT 376.370 38.935 376.540 39.105 ;
        RECT 376.370 38.575 376.540 38.745 ;
        RECT 386.950 39.295 387.120 39.465 ;
        RECT 386.950 38.935 387.120 39.105 ;
        RECT 386.950 38.575 387.120 38.745 ;
        RECT 376.370 34.185 376.540 34.355 ;
        RECT 376.370 33.825 376.540 33.995 ;
        RECT 376.370 33.465 376.540 33.635 ;
        RECT 376.370 33.105 376.540 33.275 ;
        RECT 386.950 34.185 387.120 34.355 ;
        RECT 386.950 33.825 387.120 33.995 ;
        RECT 386.950 33.465 387.120 33.635 ;
        RECT 386.950 33.105 387.120 33.275 ;
        RECT 376.370 28.715 376.540 28.885 ;
        RECT 376.370 28.355 376.540 28.525 ;
        RECT 376.370 27.995 376.540 28.165 ;
        RECT 376.370 27.635 376.540 27.805 ;
        RECT 386.950 28.715 387.120 28.885 ;
        RECT 386.950 28.355 387.120 28.525 ;
        RECT 386.950 27.995 387.120 28.165 ;
        RECT 386.950 27.635 387.120 27.805 ;
        RECT 376.370 23.245 376.540 23.415 ;
        RECT 376.370 22.885 376.540 23.055 ;
        RECT 376.370 22.525 376.540 22.695 ;
        RECT 376.370 22.165 376.540 22.335 ;
        RECT 386.950 23.245 387.120 23.415 ;
        RECT 386.950 22.885 387.120 23.055 ;
        RECT 386.950 22.525 387.120 22.695 ;
        RECT 386.950 22.165 387.120 22.335 ;
        RECT 376.370 17.775 376.540 17.945 ;
        RECT 386.950 17.775 387.120 17.945 ;
        RECT 397.530 39.295 397.700 39.465 ;
        RECT 397.530 38.935 397.700 39.105 ;
        RECT 397.530 38.575 397.700 38.745 ;
        RECT 397.530 34.185 397.700 34.355 ;
        RECT 397.530 33.825 397.700 33.995 ;
        RECT 397.530 33.465 397.700 33.635 ;
        RECT 397.530 33.105 397.700 33.275 ;
        RECT 397.530 28.715 397.700 28.885 ;
        RECT 397.530 28.355 397.700 28.525 ;
        RECT 397.530 27.995 397.700 28.165 ;
        RECT 397.530 27.635 397.700 27.805 ;
        RECT 397.530 23.245 397.700 23.415 ;
        RECT 397.530 22.885 397.700 23.055 ;
        RECT 397.530 22.525 397.700 22.695 ;
        RECT 397.530 22.165 397.700 22.335 ;
        RECT 397.530 17.775 397.700 17.945 ;
        RECT 419.310 39.645 419.480 39.815 ;
        RECT 429.890 39.645 430.060 39.815 ;
        RECT 408.730 39.285 408.900 39.455 ;
        RECT 408.730 38.925 408.900 39.095 ;
        RECT 408.730 38.565 408.900 38.735 ;
        RECT 419.310 39.285 419.480 39.455 ;
        RECT 419.310 38.925 419.480 39.095 ;
        RECT 419.310 38.565 419.480 38.735 ;
        RECT 408.730 34.175 408.900 34.345 ;
        RECT 408.730 33.815 408.900 33.985 ;
        RECT 408.730 33.455 408.900 33.625 ;
        RECT 408.730 33.095 408.900 33.265 ;
        RECT 419.310 34.175 419.480 34.345 ;
        RECT 419.310 33.815 419.480 33.985 ;
        RECT 419.310 33.455 419.480 33.625 ;
        RECT 419.310 33.095 419.480 33.265 ;
        RECT 408.730 28.705 408.900 28.875 ;
        RECT 408.730 28.345 408.900 28.515 ;
        RECT 408.730 27.985 408.900 28.155 ;
        RECT 408.730 27.625 408.900 27.795 ;
        RECT 419.310 28.705 419.480 28.875 ;
        RECT 419.310 28.345 419.480 28.515 ;
        RECT 419.310 27.985 419.480 28.155 ;
        RECT 419.310 27.625 419.480 27.795 ;
        RECT 408.730 23.235 408.900 23.405 ;
        RECT 408.730 22.875 408.900 23.045 ;
        RECT 408.730 22.515 408.900 22.685 ;
        RECT 408.730 22.155 408.900 22.325 ;
        RECT 419.310 23.235 419.480 23.405 ;
        RECT 419.310 22.875 419.480 23.045 ;
        RECT 419.310 22.515 419.480 22.685 ;
        RECT 419.310 22.155 419.480 22.325 ;
        RECT 166.540 17.255 166.710 17.425 ;
        RECT 166.540 16.895 166.710 17.065 ;
        RECT 177.930 17.285 178.100 17.455 ;
        RECT 177.930 16.925 178.100 17.095 ;
        RECT 188.510 17.285 188.680 17.455 ;
        RECT 145.380 16.535 145.550 16.705 ;
        RECT 155.960 16.535 156.130 16.705 ;
        RECT 166.540 16.535 166.710 16.705 ;
        RECT 188.510 16.925 188.680 17.095 ;
        RECT 199.090 17.285 199.260 17.455 ;
        RECT 199.090 16.925 199.260 17.095 ;
        RECT 376.370 17.415 376.540 17.585 ;
        RECT 376.370 17.055 376.540 17.225 ;
        RECT 177.930 16.565 178.100 16.735 ;
        RECT 188.510 16.565 188.680 16.735 ;
        RECT 199.090 16.565 199.260 16.735 ;
        RECT 376.370 16.695 376.540 16.865 ;
        RECT 386.950 17.415 387.120 17.585 ;
        RECT 386.950 17.055 387.120 17.225 ;
        RECT 386.950 16.695 387.120 16.865 ;
        RECT 408.730 17.765 408.900 17.935 ;
        RECT 419.310 17.765 419.480 17.935 ;
        RECT 429.890 39.285 430.060 39.455 ;
        RECT 429.890 38.925 430.060 39.095 ;
        RECT 429.890 38.565 430.060 38.735 ;
        RECT 429.890 34.175 430.060 34.345 ;
        RECT 429.890 33.815 430.060 33.985 ;
        RECT 429.890 33.455 430.060 33.625 ;
        RECT 429.890 33.095 430.060 33.265 ;
        RECT 429.890 28.705 430.060 28.875 ;
        RECT 429.890 28.345 430.060 28.515 ;
        RECT 429.890 27.985 430.060 28.155 ;
        RECT 429.890 27.625 430.060 27.795 ;
        RECT 429.890 23.235 430.060 23.405 ;
        RECT 429.890 22.875 430.060 23.045 ;
        RECT 429.890 22.515 430.060 22.685 ;
        RECT 429.890 22.155 430.060 22.325 ;
        RECT 429.890 17.765 430.060 17.935 ;
        RECT 397.530 17.415 397.700 17.585 ;
        RECT 397.530 17.055 397.700 17.225 ;
        RECT 397.530 16.695 397.700 16.865 ;
        RECT 408.730 17.405 408.900 17.575 ;
        RECT 408.730 17.045 408.900 17.215 ;
        RECT 408.730 16.685 408.900 16.855 ;
        RECT 419.310 17.405 419.480 17.575 ;
        RECT 419.310 17.045 419.480 17.215 ;
        RECT 419.310 16.685 419.480 16.855 ;
        RECT 429.890 17.405 430.060 17.575 ;
        RECT 429.890 17.045 430.060 17.215 ;
        RECT 429.890 16.685 430.060 16.855 ;
        RECT -95.840 15.015 -95.670 15.185 ;
        RECT -95.840 14.655 -95.670 14.825 ;
        RECT -95.840 14.295 -95.670 14.465 ;
        RECT -95.840 13.935 -95.670 14.105 ;
        RECT -93.260 15.015 -93.090 15.185 ;
        RECT -93.260 14.655 -93.090 14.825 ;
        RECT -93.260 14.295 -93.090 14.465 ;
        RECT -93.260 13.935 -93.090 14.105 ;
        RECT -90.680 15.015 -90.510 15.185 ;
        RECT -90.680 14.655 -90.510 14.825 ;
        RECT -90.680 14.295 -90.510 14.465 ;
        RECT -90.680 13.935 -90.510 14.105 ;
        RECT -88.100 15.015 -87.930 15.185 ;
        RECT -88.100 14.655 -87.930 14.825 ;
        RECT -88.100 14.295 -87.930 14.465 ;
        RECT -88.100 13.935 -87.930 14.105 ;
        RECT -85.520 15.015 -85.350 15.185 ;
        RECT -85.520 14.655 -85.350 14.825 ;
        RECT -85.520 14.295 -85.350 14.465 ;
        RECT -85.520 13.935 -85.350 14.105 ;
        RECT -82.940 15.015 -82.770 15.185 ;
        RECT -82.940 14.655 -82.770 14.825 ;
        RECT -82.940 14.295 -82.770 14.465 ;
        RECT -82.940 13.935 -82.770 14.105 ;
        RECT -80.360 15.015 -80.190 15.185 ;
        RECT -80.360 14.655 -80.190 14.825 ;
        RECT -80.360 14.295 -80.190 14.465 ;
        RECT -80.360 13.935 -80.190 14.105 ;
        RECT -77.780 15.015 -77.610 15.185 ;
        RECT -77.780 14.655 -77.610 14.825 ;
        RECT -77.780 14.295 -77.610 14.465 ;
        RECT -77.780 13.935 -77.610 14.105 ;
        RECT -75.200 15.015 -75.030 15.185 ;
        RECT -75.200 14.655 -75.030 14.825 ;
        RECT -75.200 14.295 -75.030 14.465 ;
        RECT -75.200 13.935 -75.030 14.105 ;
        RECT -72.620 15.015 -72.450 15.185 ;
        RECT -72.620 14.655 -72.450 14.825 ;
        RECT -72.620 14.295 -72.450 14.465 ;
        RECT -72.620 13.935 -72.450 14.105 ;
        RECT -50.930 14.560 -50.760 14.730 ;
        RECT -50.930 14.200 -50.760 14.370 ;
        RECT -50.930 13.840 -50.760 14.010 ;
        RECT -50.930 13.480 -50.760 13.650 ;
        RECT -48.350 14.560 -48.180 14.730 ;
        RECT -48.350 14.200 -48.180 14.370 ;
        RECT -48.350 13.840 -48.180 14.010 ;
        RECT -48.350 13.480 -48.180 13.650 ;
        RECT -45.770 14.560 -45.600 14.730 ;
        RECT -45.770 14.200 -45.600 14.370 ;
        RECT -45.770 13.840 -45.600 14.010 ;
        RECT -45.770 13.480 -45.600 13.650 ;
        RECT -43.190 14.560 -43.020 14.730 ;
        RECT -43.190 14.200 -43.020 14.370 ;
        RECT -43.190 13.840 -43.020 14.010 ;
        RECT -43.190 13.480 -43.020 13.650 ;
        RECT -40.610 14.560 -40.440 14.730 ;
        RECT -40.610 14.200 -40.440 14.370 ;
        RECT -40.610 13.840 -40.440 14.010 ;
        RECT -40.610 13.480 -40.440 13.650 ;
        RECT -38.030 14.560 -37.860 14.730 ;
        RECT -38.030 14.200 -37.860 14.370 ;
        RECT -38.030 13.840 -37.860 14.010 ;
        RECT -38.030 13.480 -37.860 13.650 ;
        RECT -35.450 14.560 -35.280 14.730 ;
        RECT -35.450 14.200 -35.280 14.370 ;
        RECT -35.450 13.840 -35.280 14.010 ;
        RECT -35.450 13.480 -35.280 13.650 ;
        RECT -32.870 14.560 -32.700 14.730 ;
        RECT -32.870 14.200 -32.700 14.370 ;
        RECT -32.870 13.840 -32.700 14.010 ;
        RECT -32.870 13.480 -32.700 13.650 ;
        RECT -30.290 14.560 -30.120 14.730 ;
        RECT -30.290 14.200 -30.120 14.370 ;
        RECT -30.290 13.840 -30.120 14.010 ;
        RECT -30.290 13.480 -30.120 13.650 ;
        RECT -27.710 14.560 -27.540 14.730 ;
        RECT -27.710 14.200 -27.540 14.370 ;
        RECT -27.710 13.840 -27.540 14.010 ;
        RECT -27.710 13.480 -27.540 13.650 ;
      LAYER met1 ;
        RECT 112.600 213.740 112.830 215.320 ;
        RECT 123.180 213.740 123.410 215.320 ;
        RECT 133.760 213.740 133.990 215.320 ;
        RECT 145.210 213.820 145.440 215.400 ;
        RECT 155.790 213.820 156.020 215.400 ;
        RECT 166.370 213.820 166.600 215.400 ;
        RECT 177.760 213.850 177.990 215.430 ;
        RECT 188.340 213.850 188.570 215.430 ;
        RECT 198.920 213.850 199.150 215.430 ;
        RECT 112.600 208.270 112.830 209.850 ;
        RECT 123.180 208.270 123.410 209.850 ;
        RECT 133.760 208.270 133.990 209.850 ;
        RECT 145.210 208.350 145.440 209.930 ;
        RECT 155.790 208.350 156.020 209.930 ;
        RECT 166.370 208.350 166.600 209.930 ;
        RECT 177.760 208.380 177.990 209.960 ;
        RECT 188.340 208.380 188.570 209.960 ;
        RECT 198.920 208.380 199.150 209.960 ;
        RECT 112.600 202.800 112.830 204.380 ;
        RECT 123.180 202.800 123.410 204.380 ;
        RECT 133.760 202.800 133.990 204.380 ;
        RECT 145.210 202.880 145.440 204.460 ;
        RECT 155.790 202.880 156.020 204.460 ;
        RECT 166.370 202.880 166.600 204.460 ;
        RECT 177.760 202.910 177.990 204.490 ;
        RECT 188.340 202.910 188.570 204.490 ;
        RECT 198.920 202.910 199.150 204.490 ;
        RECT 112.600 197.330 112.830 198.910 ;
        RECT 123.180 197.330 123.410 198.910 ;
        RECT 133.760 197.330 133.990 198.910 ;
        RECT 145.210 197.410 145.440 198.990 ;
        RECT 155.790 197.410 156.020 198.990 ;
        RECT 166.370 197.410 166.600 198.990 ;
        RECT 177.760 197.440 177.990 199.020 ;
        RECT 188.340 197.440 188.570 199.020 ;
        RECT 198.920 197.440 199.150 199.020 ;
        RECT 112.600 191.860 112.830 193.440 ;
        RECT 123.180 191.860 123.410 193.440 ;
        RECT 133.760 191.860 133.990 193.440 ;
        RECT 145.210 191.940 145.440 193.520 ;
        RECT 155.790 191.940 156.020 193.520 ;
        RECT 166.370 191.940 166.600 193.520 ;
        RECT 177.760 191.970 177.990 193.550 ;
        RECT 188.340 191.970 188.570 193.550 ;
        RECT 198.920 191.970 199.150 193.550 ;
        RECT 112.600 184.660 112.830 186.240 ;
        RECT 123.180 184.660 123.410 186.240 ;
        RECT 133.760 184.660 133.990 186.240 ;
        RECT 145.210 184.740 145.440 186.320 ;
        RECT 155.790 184.740 156.020 186.320 ;
        RECT 166.370 184.740 166.600 186.320 ;
        RECT 177.760 184.770 177.990 186.350 ;
        RECT 188.340 184.770 188.570 186.350 ;
        RECT 198.920 184.770 199.150 186.350 ;
        RECT 112.600 179.190 112.830 180.770 ;
        RECT 123.180 179.190 123.410 180.770 ;
        RECT 133.760 179.190 133.990 180.770 ;
        RECT 145.210 179.270 145.440 180.850 ;
        RECT 155.790 179.270 156.020 180.850 ;
        RECT 166.370 179.270 166.600 180.850 ;
        RECT 177.760 179.300 177.990 180.880 ;
        RECT 188.340 179.300 188.570 180.880 ;
        RECT 198.920 179.300 199.150 180.880 ;
        RECT 112.600 173.720 112.830 175.300 ;
        RECT 123.180 173.720 123.410 175.300 ;
        RECT 133.760 173.720 133.990 175.300 ;
        RECT 145.210 173.800 145.440 175.380 ;
        RECT 155.790 173.800 156.020 175.380 ;
        RECT 166.370 173.800 166.600 175.380 ;
        RECT 177.760 173.830 177.990 175.410 ;
        RECT 188.340 173.830 188.570 175.410 ;
        RECT 198.920 173.830 199.150 175.410 ;
        RECT 112.600 168.250 112.830 169.830 ;
        RECT 123.180 168.250 123.410 169.830 ;
        RECT 133.760 168.250 133.990 169.830 ;
        RECT 145.210 168.330 145.440 169.910 ;
        RECT 155.790 168.330 156.020 169.910 ;
        RECT 166.370 168.330 166.600 169.910 ;
        RECT 177.760 168.360 177.990 169.940 ;
        RECT 188.340 168.360 188.570 169.940 ;
        RECT 198.920 168.360 199.150 169.940 ;
        RECT 112.600 162.780 112.830 164.360 ;
        RECT 123.180 162.780 123.410 164.360 ;
        RECT 133.760 162.780 133.990 164.360 ;
        RECT 145.210 162.860 145.440 164.440 ;
        RECT 155.790 162.860 156.020 164.440 ;
        RECT 166.370 162.860 166.600 164.440 ;
        RECT 177.760 162.890 177.990 164.470 ;
        RECT 188.340 162.890 188.570 164.470 ;
        RECT 198.920 162.890 199.150 164.470 ;
        RECT 112.600 155.490 112.830 157.070 ;
        RECT 123.180 155.490 123.410 157.070 ;
        RECT 133.760 155.490 133.990 157.070 ;
        RECT 145.210 155.570 145.440 157.150 ;
        RECT 155.790 155.570 156.020 157.150 ;
        RECT 166.370 155.570 166.600 157.150 ;
        RECT 177.760 155.600 177.990 157.180 ;
        RECT 188.340 155.600 188.570 157.180 ;
        RECT 198.920 155.600 199.150 157.180 ;
        RECT 112.600 150.020 112.830 151.600 ;
        RECT 123.180 150.020 123.410 151.600 ;
        RECT 133.760 150.020 133.990 151.600 ;
        RECT 145.210 150.100 145.440 151.680 ;
        RECT 155.790 150.100 156.020 151.680 ;
        RECT 166.370 150.100 166.600 151.680 ;
        RECT 177.760 150.130 177.990 151.710 ;
        RECT 188.340 150.130 188.570 151.710 ;
        RECT 198.920 150.130 199.150 151.710 ;
        RECT 112.600 144.550 112.830 146.130 ;
        RECT 123.180 144.550 123.410 146.130 ;
        RECT 133.760 144.550 133.990 146.130 ;
        RECT 145.210 144.630 145.440 146.210 ;
        RECT 155.790 144.630 156.020 146.210 ;
        RECT 166.370 144.630 166.600 146.210 ;
        RECT 177.760 144.660 177.990 146.240 ;
        RECT 188.340 144.660 188.570 146.240 ;
        RECT 198.920 144.660 199.150 146.240 ;
        RECT 112.600 139.080 112.830 140.660 ;
        RECT 123.180 139.080 123.410 140.660 ;
        RECT 133.760 139.080 133.990 140.660 ;
        RECT 145.210 139.160 145.440 140.740 ;
        RECT 155.790 139.160 156.020 140.740 ;
        RECT 166.370 139.160 166.600 140.740 ;
        RECT 177.760 139.190 177.990 140.770 ;
        RECT 188.340 139.190 188.570 140.770 ;
        RECT 198.920 139.190 199.150 140.770 ;
        RECT 112.600 133.610 112.830 135.190 ;
        RECT 123.180 133.610 123.410 135.190 ;
        RECT 133.760 133.610 133.990 135.190 ;
        RECT 145.210 133.690 145.440 135.270 ;
        RECT 155.790 133.690 156.020 135.270 ;
        RECT 166.370 133.690 166.600 135.270 ;
        RECT 177.760 133.720 177.990 135.300 ;
        RECT 188.340 133.720 188.570 135.300 ;
        RECT 198.920 133.720 199.150 135.300 ;
        RECT 112.600 126.310 112.830 127.890 ;
        RECT 123.180 126.310 123.410 127.890 ;
        RECT 133.760 126.310 133.990 127.890 ;
        RECT 145.210 126.390 145.440 127.970 ;
        RECT 155.790 126.390 156.020 127.970 ;
        RECT 166.370 126.390 166.600 127.970 ;
        RECT 177.760 126.420 177.990 128.000 ;
        RECT 188.340 126.420 188.570 128.000 ;
        RECT 198.920 126.420 199.150 128.000 ;
        RECT 376.310 126.180 376.540 127.760 ;
        RECT 386.890 126.180 387.120 127.760 ;
        RECT 397.470 126.180 397.700 127.760 ;
        RECT 408.620 126.170 408.850 127.750 ;
        RECT 419.200 126.170 419.430 127.750 ;
        RECT 429.780 126.170 430.010 127.750 ;
        RECT 112.600 120.840 112.830 122.420 ;
        RECT 123.180 120.840 123.410 122.420 ;
        RECT 133.760 120.840 133.990 122.420 ;
        RECT 145.210 120.920 145.440 122.500 ;
        RECT 155.790 120.920 156.020 122.500 ;
        RECT 166.370 120.920 166.600 122.500 ;
        RECT 177.760 120.950 177.990 122.530 ;
        RECT 188.340 120.950 188.570 122.530 ;
        RECT 198.920 120.950 199.150 122.530 ;
        RECT 376.310 120.710 376.540 122.290 ;
        RECT 386.890 120.710 387.120 122.290 ;
        RECT 397.470 120.710 397.700 122.290 ;
        RECT 408.620 120.700 408.850 122.280 ;
        RECT 419.200 120.700 419.430 122.280 ;
        RECT 429.780 120.700 430.010 122.280 ;
        RECT 112.600 115.370 112.830 116.950 ;
        RECT 123.180 115.370 123.410 116.950 ;
        RECT 133.760 115.370 133.990 116.950 ;
        RECT 145.210 115.450 145.440 117.030 ;
        RECT 155.790 115.450 156.020 117.030 ;
        RECT 166.370 115.450 166.600 117.030 ;
        RECT 177.760 115.480 177.990 117.060 ;
        RECT 188.340 115.480 188.570 117.060 ;
        RECT 198.920 115.480 199.150 117.060 ;
        RECT 376.310 115.240 376.540 116.820 ;
        RECT 386.890 115.240 387.120 116.820 ;
        RECT 397.470 115.240 397.700 116.820 ;
        RECT 408.620 115.230 408.850 116.810 ;
        RECT 419.200 115.230 419.430 116.810 ;
        RECT 429.780 115.230 430.010 116.810 ;
        RECT 112.600 109.900 112.830 111.480 ;
        RECT 123.180 109.900 123.410 111.480 ;
        RECT 133.760 109.900 133.990 111.480 ;
        RECT 145.210 109.980 145.440 111.560 ;
        RECT 155.790 109.980 156.020 111.560 ;
        RECT 166.370 109.980 166.600 111.560 ;
        RECT 177.760 110.010 177.990 111.590 ;
        RECT 188.340 110.010 188.570 111.590 ;
        RECT 198.920 110.010 199.150 111.590 ;
        RECT 376.310 109.770 376.540 111.350 ;
        RECT 386.890 109.770 387.120 111.350 ;
        RECT 397.470 109.770 397.700 111.350 ;
        RECT 408.620 109.760 408.850 111.340 ;
        RECT 419.200 109.760 419.430 111.340 ;
        RECT 429.780 109.760 430.010 111.340 ;
        RECT 112.600 104.430 112.830 106.010 ;
        RECT 123.180 104.430 123.410 106.010 ;
        RECT 133.760 104.430 133.990 106.010 ;
        RECT 145.210 104.510 145.440 106.090 ;
        RECT 155.790 104.510 156.020 106.090 ;
        RECT 166.370 104.510 166.600 106.090 ;
        RECT 177.760 104.540 177.990 106.120 ;
        RECT 188.340 104.540 188.570 106.120 ;
        RECT 198.920 104.540 199.150 106.120 ;
        RECT 376.310 104.920 376.540 105.880 ;
        RECT 112.600 96.990 112.830 98.570 ;
        RECT 123.180 96.990 123.410 98.570 ;
        RECT 133.760 96.990 133.990 98.570 ;
        RECT 145.210 97.070 145.440 98.650 ;
        RECT 155.790 97.070 156.020 98.650 ;
        RECT 166.370 97.070 166.600 98.650 ;
        RECT 177.760 97.100 177.990 98.680 ;
        RECT 188.340 97.100 188.570 98.680 ;
        RECT 198.920 97.100 199.150 98.680 ;
        RECT 376.180 97.660 376.680 104.920 ;
        RECT 386.890 104.300 387.120 105.880 ;
        RECT 397.470 104.300 397.700 105.880 ;
        RECT 408.620 105.190 408.850 105.870 ;
        RECT 376.340 96.990 376.570 97.660 ;
        RECT 386.920 96.990 387.150 98.570 ;
        RECT 397.500 96.990 397.730 98.570 ;
        RECT 408.590 97.930 409.090 105.190 ;
        RECT 419.200 104.290 419.430 105.870 ;
        RECT 429.780 104.290 430.010 105.870 ;
        RECT 408.660 97.050 408.890 97.930 ;
        RECT 419.240 97.050 419.470 98.630 ;
        RECT 429.820 97.050 430.050 98.630 ;
        RECT 112.600 91.520 112.830 93.100 ;
        RECT 123.180 91.520 123.410 93.100 ;
        RECT 133.760 91.520 133.990 93.100 ;
        RECT 145.210 91.600 145.440 93.180 ;
        RECT 155.790 91.600 156.020 93.180 ;
        RECT 166.370 91.600 166.600 93.180 ;
        RECT 177.760 91.630 177.990 93.210 ;
        RECT 188.340 91.630 188.570 93.210 ;
        RECT 198.920 91.630 199.150 93.210 ;
        RECT 376.340 91.520 376.570 93.100 ;
        RECT 386.920 91.520 387.150 93.100 ;
        RECT 397.500 91.520 397.730 93.100 ;
        RECT 408.660 91.580 408.890 93.160 ;
        RECT 419.240 91.580 419.470 93.160 ;
        RECT 429.820 91.580 430.050 93.160 ;
        RECT 112.600 86.050 112.830 87.630 ;
        RECT 123.180 86.050 123.410 87.630 ;
        RECT 133.760 86.050 133.990 87.630 ;
        RECT 145.210 86.130 145.440 87.710 ;
        RECT 155.790 86.130 156.020 87.710 ;
        RECT 166.370 86.130 166.600 87.710 ;
        RECT 177.760 86.160 177.990 87.740 ;
        RECT 188.340 86.160 188.570 87.740 ;
        RECT 198.920 86.160 199.150 87.740 ;
        RECT 376.340 86.050 376.570 87.630 ;
        RECT 386.920 86.050 387.150 87.630 ;
        RECT 397.500 86.050 397.730 87.630 ;
        RECT 408.660 86.110 408.890 87.690 ;
        RECT 419.240 86.110 419.470 87.690 ;
        RECT 429.820 86.110 430.050 87.690 ;
        RECT 112.600 80.580 112.830 82.160 ;
        RECT 123.180 80.580 123.410 82.160 ;
        RECT 133.760 80.580 133.990 82.160 ;
        RECT 145.210 80.660 145.440 82.240 ;
        RECT 155.790 80.660 156.020 82.240 ;
        RECT 166.370 80.660 166.600 82.240 ;
        RECT 177.760 80.690 177.990 82.270 ;
        RECT 188.340 80.690 188.570 82.270 ;
        RECT 198.920 80.690 199.150 82.270 ;
        RECT 376.340 80.580 376.570 82.160 ;
        RECT 386.920 80.580 387.150 82.160 ;
        RECT 397.500 80.580 397.730 82.160 ;
        RECT 408.660 80.640 408.890 82.220 ;
        RECT 419.240 80.640 419.470 82.220 ;
        RECT 429.820 80.640 430.050 82.220 ;
        RECT 112.600 75.110 112.830 76.690 ;
        RECT 123.180 75.110 123.410 76.690 ;
        RECT 133.760 75.110 133.990 76.690 ;
        RECT 145.210 75.190 145.440 76.770 ;
        RECT 155.790 75.190 156.020 76.770 ;
        RECT 166.370 75.190 166.600 76.770 ;
        RECT 177.760 75.220 177.990 76.800 ;
        RECT 188.340 75.220 188.570 76.800 ;
        RECT 198.920 75.220 199.150 76.800 ;
        RECT 376.340 75.590 376.570 76.690 ;
        RECT 112.650 67.710 112.880 69.290 ;
        RECT 123.230 67.710 123.460 69.290 ;
        RECT 133.810 67.710 134.040 69.290 ;
        RECT 145.260 67.790 145.490 69.370 ;
        RECT 155.840 67.790 156.070 69.370 ;
        RECT 166.420 67.790 166.650 69.370 ;
        RECT 177.810 67.820 178.040 69.400 ;
        RECT 188.390 67.820 188.620 69.400 ;
        RECT 198.970 67.820 199.200 69.400 ;
        RECT 376.180 68.330 376.680 75.590 ;
        RECT 386.920 75.110 387.150 76.690 ;
        RECT 397.500 75.110 397.730 76.690 ;
        RECT 408.660 75.760 408.890 76.750 ;
        RECT 408.370 75.170 408.890 75.760 ;
        RECT 419.240 75.170 419.470 76.750 ;
        RECT 429.820 75.170 430.050 76.750 ;
        RECT 376.340 67.700 376.570 68.330 ;
        RECT 386.920 67.700 387.150 69.280 ;
        RECT 397.500 67.700 397.730 69.280 ;
        RECT 408.370 69.270 408.870 75.170 ;
        RECT 408.370 68.500 408.910 69.270 ;
        RECT 408.680 67.690 408.910 68.500 ;
        RECT 419.260 67.690 419.490 69.270 ;
        RECT 429.840 67.690 430.070 69.270 ;
        RECT 112.650 62.240 112.880 63.820 ;
        RECT 123.230 62.240 123.460 63.820 ;
        RECT 133.810 62.240 134.040 63.820 ;
        RECT 145.260 62.320 145.490 63.900 ;
        RECT 155.840 62.320 156.070 63.900 ;
        RECT 166.420 62.320 166.650 63.900 ;
        RECT 177.810 62.350 178.040 63.930 ;
        RECT 188.390 62.350 188.620 63.930 ;
        RECT 198.970 62.350 199.200 63.930 ;
        RECT 376.340 62.230 376.570 63.810 ;
        RECT 386.920 62.230 387.150 63.810 ;
        RECT 397.500 62.230 397.730 63.810 ;
        RECT 408.680 62.220 408.910 63.800 ;
        RECT 419.260 62.220 419.490 63.800 ;
        RECT 429.840 62.220 430.070 63.800 ;
        RECT 112.650 56.770 112.880 58.350 ;
        RECT 123.230 56.770 123.460 58.350 ;
        RECT 133.810 56.770 134.040 58.350 ;
        RECT 145.260 56.850 145.490 58.430 ;
        RECT 155.840 56.850 156.070 58.430 ;
        RECT 166.420 56.850 166.650 58.430 ;
        RECT 177.810 56.880 178.040 58.460 ;
        RECT 188.390 56.880 188.620 58.460 ;
        RECT 198.970 56.880 199.200 58.460 ;
        RECT 376.340 56.760 376.570 58.340 ;
        RECT 386.920 56.760 387.150 58.340 ;
        RECT 397.500 56.760 397.730 58.340 ;
        RECT 408.680 56.750 408.910 58.330 ;
        RECT 419.260 56.750 419.490 58.330 ;
        RECT 429.840 56.750 430.070 58.330 ;
        RECT 112.650 51.300 112.880 52.880 ;
        RECT 123.230 51.300 123.460 52.880 ;
        RECT 133.810 51.300 134.040 52.880 ;
        RECT 145.260 51.380 145.490 52.960 ;
        RECT 155.840 51.380 156.070 52.960 ;
        RECT 166.420 51.380 166.650 52.960 ;
        RECT 177.810 51.410 178.040 52.990 ;
        RECT 188.390 51.410 188.620 52.990 ;
        RECT 198.970 51.410 199.200 52.990 ;
        RECT 376.340 51.290 376.570 52.870 ;
        RECT 386.920 51.290 387.150 52.870 ;
        RECT 397.500 51.290 397.730 52.870 ;
        RECT 408.680 51.280 408.910 52.860 ;
        RECT 419.260 51.280 419.490 52.860 ;
        RECT 429.840 51.280 430.070 52.860 ;
        RECT 112.650 45.830 112.880 47.410 ;
        RECT 123.230 45.830 123.460 47.410 ;
        RECT 133.810 45.830 134.040 47.410 ;
        RECT 145.260 45.910 145.490 47.490 ;
        RECT 155.840 45.910 156.070 47.490 ;
        RECT 166.420 45.910 166.650 47.490 ;
        RECT 177.810 45.940 178.040 47.520 ;
        RECT 188.390 45.940 188.620 47.520 ;
        RECT 198.970 45.940 199.200 47.520 ;
        RECT 376.340 46.320 376.570 47.400 ;
        RECT 112.740 38.170 112.970 39.750 ;
        RECT 123.320 38.170 123.550 39.750 ;
        RECT 133.900 38.170 134.130 39.750 ;
        RECT 145.350 38.250 145.580 39.830 ;
        RECT 155.930 38.250 156.160 39.830 ;
        RECT 166.510 38.250 166.740 39.830 ;
        RECT 177.900 38.280 178.130 39.860 ;
        RECT 188.480 38.280 188.710 39.860 ;
        RECT 199.060 38.280 199.290 39.860 ;
        RECT 376.240 39.060 376.740 46.320 ;
        RECT 386.920 45.820 387.150 47.400 ;
        RECT 397.500 45.820 397.730 47.400 ;
        RECT 408.680 46.600 408.910 47.390 ;
        RECT 376.340 38.410 376.570 39.060 ;
        RECT 386.920 38.410 387.150 39.990 ;
        RECT 397.500 38.410 397.730 39.990 ;
        RECT 408.530 39.340 409.030 46.600 ;
        RECT 419.260 45.810 419.490 47.390 ;
        RECT 429.840 45.810 430.070 47.390 ;
        RECT 408.700 38.400 408.930 39.340 ;
        RECT 419.280 38.400 419.510 39.980 ;
        RECT 429.860 38.400 430.090 39.980 ;
        RECT 112.740 32.700 112.970 34.280 ;
        RECT 123.320 32.700 123.550 34.280 ;
        RECT 133.900 32.700 134.130 34.280 ;
        RECT 145.350 32.780 145.580 34.360 ;
        RECT 155.930 32.780 156.160 34.360 ;
        RECT 166.510 32.780 166.740 34.360 ;
        RECT 177.900 32.810 178.130 34.390 ;
        RECT 188.480 32.810 188.710 34.390 ;
        RECT 199.060 32.810 199.290 34.390 ;
        RECT 376.340 32.940 376.570 34.520 ;
        RECT 386.920 32.940 387.150 34.520 ;
        RECT 397.500 32.940 397.730 34.520 ;
        RECT 408.700 32.930 408.930 34.510 ;
        RECT 419.280 32.930 419.510 34.510 ;
        RECT 429.860 32.930 430.090 34.510 ;
        RECT 112.740 27.230 112.970 28.810 ;
        RECT 123.320 27.230 123.550 28.810 ;
        RECT 133.900 27.230 134.130 28.810 ;
        RECT 145.350 27.310 145.580 28.890 ;
        RECT 155.930 27.310 156.160 28.890 ;
        RECT 166.510 27.310 166.740 28.890 ;
        RECT 177.900 27.340 178.130 28.920 ;
        RECT 188.480 27.340 188.710 28.920 ;
        RECT 199.060 27.340 199.290 28.920 ;
        RECT 376.340 27.470 376.570 29.050 ;
        RECT 386.920 27.470 387.150 29.050 ;
        RECT 397.500 27.470 397.730 29.050 ;
        RECT 408.700 27.460 408.930 29.040 ;
        RECT 419.280 27.460 419.510 29.040 ;
        RECT 429.860 27.460 430.090 29.040 ;
        RECT 112.740 21.760 112.970 23.340 ;
        RECT 123.320 21.760 123.550 23.340 ;
        RECT 133.900 21.760 134.130 23.340 ;
        RECT 145.350 21.840 145.580 23.420 ;
        RECT 155.930 21.840 156.160 23.420 ;
        RECT 166.510 21.840 166.740 23.420 ;
        RECT 177.900 21.870 178.130 23.450 ;
        RECT 188.480 21.870 188.710 23.450 ;
        RECT 199.060 21.870 199.290 23.450 ;
        RECT 376.340 22.000 376.570 23.580 ;
        RECT 386.920 22.000 387.150 23.580 ;
        RECT 397.500 22.000 397.730 23.580 ;
        RECT 408.700 21.990 408.930 23.570 ;
        RECT 419.280 21.990 419.510 23.570 ;
        RECT 429.860 21.990 430.090 23.570 ;
        RECT -75.245 16.500 -75.015 18.685 ;
        RECT -96.080 15.920 -72.130 16.500 ;
        RECT 112.740 16.290 112.970 17.870 ;
        RECT 123.320 16.290 123.550 17.870 ;
        RECT 133.900 16.290 134.130 17.870 ;
        RECT 145.350 16.370 145.580 17.950 ;
        RECT 155.930 16.370 156.160 17.950 ;
        RECT 166.510 16.370 166.740 17.950 ;
        RECT 177.900 16.400 178.130 17.980 ;
        RECT 188.480 16.400 188.710 17.980 ;
        RECT 199.060 16.950 199.290 17.980 ;
        RECT 376.340 17.080 376.570 18.110 ;
        RECT -95.875 15.350 -95.665 15.920 ;
        RECT -93.295 15.350 -93.085 15.920 ;
        RECT -90.725 15.350 -90.515 15.920 ;
        RECT -88.165 15.350 -87.955 15.920 ;
        RECT -85.525 15.350 -85.315 15.920 ;
        RECT -95.875 15.015 -95.640 15.350 ;
        RECT -93.295 15.055 -93.060 15.350 ;
        RECT -90.725 15.055 -90.480 15.350 ;
        RECT -95.870 13.770 -95.640 15.015 ;
        RECT -93.290 13.770 -93.060 15.055 ;
        RECT -90.710 13.770 -90.480 15.055 ;
        RECT -88.165 15.035 -87.900 15.350 ;
        RECT -88.130 13.770 -87.900 15.035 ;
        RECT -85.550 15.015 -85.315 15.350 ;
        RECT -82.985 15.350 -82.775 15.920 ;
        RECT -80.345 15.350 -80.135 15.920 ;
        RECT -77.795 15.350 -77.585 15.920 ;
        RECT -75.245 15.905 -75.015 15.920 ;
        RECT -75.235 15.350 -75.025 15.905 ;
        RECT -72.615 15.350 -72.405 15.920 ;
        RECT -85.550 13.770 -85.320 15.015 ;
        RECT -82.985 14.985 -82.740 15.350 ;
        RECT -82.970 13.770 -82.740 14.985 ;
        RECT -80.390 14.885 -80.135 15.350 ;
        RECT -80.390 13.770 -80.160 14.885 ;
        RECT -77.810 13.770 -77.580 15.350 ;
        RECT -75.235 14.925 -75.000 15.350 ;
        RECT -75.230 13.770 -75.000 14.925 ;
        RECT -72.650 15.015 -72.405 15.350 ;
        RECT -72.650 13.770 -72.420 15.015 ;
        RECT -50.960 13.570 -50.730 14.895 ;
        RECT -50.965 12.640 -50.725 13.570 ;
        RECT -48.380 13.490 -48.150 14.895 ;
        RECT -45.800 13.510 -45.570 14.895 ;
        RECT -43.220 13.570 -42.990 14.895 ;
        RECT -48.405 13.315 -48.150 13.490 ;
        RECT -48.405 12.640 -48.165 13.315 ;
        RECT -45.805 12.640 -45.565 13.510 ;
        RECT -43.245 13.315 -42.990 13.570 ;
        RECT -40.640 13.530 -40.410 14.895 ;
        RECT -38.060 13.570 -37.830 14.895 ;
        RECT -40.665 13.315 -40.410 13.530 ;
        RECT -43.245 12.640 -43.005 13.315 ;
        RECT -40.665 12.640 -40.425 13.315 ;
        RECT -38.065 12.640 -37.825 13.570 ;
        RECT -35.480 13.550 -35.250 14.895 ;
        RECT -35.485 12.640 -35.245 13.550 ;
        RECT -32.900 13.490 -32.670 14.895 ;
        RECT -30.320 13.530 -30.090 14.895 ;
        RECT -32.905 12.640 -32.665 13.490 ;
        RECT -30.345 13.315 -30.090 13.530 ;
        RECT -27.740 13.510 -27.510 14.895 ;
        RECT -27.740 13.315 -27.455 13.510 ;
        RECT -30.345 12.640 -30.105 13.315 ;
        RECT -27.695 12.640 -27.455 13.315 ;
        RECT 198.450 12.970 199.910 16.950 ;
        RECT 207.210 12.970 209.990 13.850 ;
        RECT 375.710 12.970 376.900 17.080 ;
        RECT 386.920 16.530 387.150 18.110 ;
        RECT 397.500 16.530 397.730 18.110 ;
        RECT 408.700 16.520 408.930 18.100 ;
        RECT 419.280 16.520 419.510 18.100 ;
        RECT 429.860 16.520 430.090 18.100 ;
        RECT -51.310 11.950 -27.060 12.640 ;
        RECT 198.440 11.960 376.900 12.970 ;
        RECT -27.765 10.030 -27.455 11.950 ;
        RECT 207.210 11.050 209.990 11.960 ;
        RECT 375.710 11.420 376.900 11.960 ;
      LAYER via ;
        RECT -95.915 15.920 -72.295 16.500 ;
        RECT -51.155 12.005 -27.215 12.585 ;
        RECT 207.350 11.200 209.850 13.700 ;
      LAYER met2 ;
        RECT -97.290 16.550 -93.120 16.630 ;
        RECT -76.720 16.550 -59.520 16.590 ;
        RECT -97.290 16.000 -59.520 16.550 ;
        RECT -97.290 15.870 -72.180 16.000 ;
        RECT -97.290 15.640 -93.120 15.870 ;
        RECT -60.370 12.440 -59.570 16.000 ;
        RECT 207.260 13.170 209.940 13.900 ;
        RECT -29.020 12.690 209.940 13.170 ;
        RECT -51.260 12.440 209.940 12.690 ;
        RECT -60.370 12.060 209.940 12.440 ;
        RECT -60.370 12.050 -4.870 12.060 ;
        RECT -60.370 11.900 -27.110 12.050 ;
        RECT -60.370 11.850 -43.170 11.900 ;
        RECT 207.260 11.000 209.940 12.060 ;
      LAYER via2 ;
        RECT -97.145 15.795 -93.265 16.475 ;
      LAYER met3 ;
        RECT -129.710 16.605 -96.060 17.210 ;
        RECT -129.710 15.665 -93.070 16.605 ;
        RECT -129.710 15.080 -96.060 15.665 ;
    END
  END vcap
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -98.220 351.200 -70.530 358.370 ;
        RECT 653.990 351.075 655.320 352.275 ;
        RECT 657.570 351.935 659.795 352.435 ;
        RECT 663.040 351.935 670.640 352.265 ;
        RECT 653.840 350.645 655.540 351.075 ;
        RECT 657.570 351.065 672.890 351.935 ;
        RECT 675.620 351.895 677.845 352.395 ;
        RECT 681.090 351.895 688.690 352.225 ;
        RECT 693.210 351.915 695.435 352.415 ;
        RECT 698.680 351.915 706.280 352.245 ;
        RECT 711.060 351.915 713.285 352.415 ;
        RECT 716.530 351.915 724.130 352.245 ;
        RECT 729.320 351.915 731.545 352.415 ;
        RECT 734.790 351.915 742.390 352.245 ;
        RECT 657.420 350.635 673.040 351.065 ;
        RECT 675.620 351.025 690.940 351.895 ;
        RECT 693.210 351.045 708.530 351.915 ;
        RECT 711.060 351.045 726.380 351.915 ;
        RECT 729.320 351.045 744.640 351.915 ;
        RECT 747.090 351.885 749.315 352.385 ;
        RECT 752.560 351.885 760.160 352.215 ;
        RECT 675.470 350.595 691.090 351.025 ;
        RECT 693.060 350.615 708.680 351.045 ;
        RECT 710.910 350.615 726.530 351.045 ;
        RECT 729.170 350.615 744.790 351.045 ;
        RECT 747.090 351.015 762.410 351.885 ;
        RECT 765.130 351.805 767.355 352.305 ;
        RECT 770.600 351.805 778.200 352.135 ;
        RECT 783.290 351.845 785.515 352.345 ;
        RECT 788.760 351.845 796.360 352.175 ;
        RECT 801.670 351.855 803.895 352.355 ;
        RECT 807.140 351.855 814.740 352.185 ;
        RECT 746.940 350.585 762.560 351.015 ;
        RECT 765.130 350.935 780.450 351.805 ;
        RECT 783.290 350.975 798.610 351.845 ;
        RECT 801.670 350.985 816.990 351.855 ;
        RECT 820.470 351.835 822.695 352.335 ;
        RECT 825.940 351.835 833.540 352.165 ;
        RECT 764.980 350.505 780.600 350.935 ;
        RECT 783.140 350.545 798.760 350.975 ;
        RECT 801.520 350.555 817.140 350.985 ;
        RECT 820.470 350.965 835.790 351.835 ;
        RECT 820.320 350.535 835.940 350.965 ;
        RECT 838.940 350.945 840.270 352.145 ;
        RECT 838.790 350.515 840.490 350.945 ;
        RECT 783.850 343.675 785.160 344.005 ;
        RECT 783.850 342.805 787.170 343.675 ;
        RECT 790.410 342.835 791.740 344.035 ;
        RECT 793.870 343.765 796.095 344.265 ;
        RECT 799.340 343.765 806.940 344.095 ;
        RECT 793.870 342.895 809.190 343.765 ;
        RECT 813.230 343.675 815.455 344.175 ;
        RECT 818.700 343.675 826.300 344.005 ;
        RECT 783.700 342.375 787.320 342.805 ;
        RECT 790.260 342.405 791.960 342.835 ;
        RECT 793.720 342.465 809.340 342.895 ;
        RECT 813.230 342.805 828.550 343.675 ;
        RECT 813.080 342.375 828.700 342.805 ;
        RECT 665.220 329.585 666.530 329.915 ;
        RECT 670.850 329.585 672.160 329.915 ;
        RECT 678.220 329.815 679.260 329.820 ;
        RECT 663.210 328.715 666.530 329.585 ;
        RECT 668.840 328.715 672.160 329.585 ;
        RECT 676.590 329.485 679.260 329.815 ;
        RECT 674.870 328.790 679.260 329.485 ;
        RECT 595.390 326.925 596.720 328.125 ;
        RECT 635.350 327.375 636.680 328.575 ;
        RECT 639.540 327.465 640.870 328.665 ;
        RECT 643.640 328.640 644.970 328.645 ;
        RECT 595.240 326.495 596.940 326.925 ;
        RECT 605.200 323.670 606.350 327.180 ;
        RECT 610.210 325.140 613.920 326.660 ;
        RECT 617.800 325.140 621.510 326.630 ;
        RECT 610.210 323.670 621.510 325.140 ;
        RECT 625.380 323.670 626.560 327.310 ;
        RECT 635.130 326.945 636.830 327.375 ;
        RECT 639.320 327.035 641.020 327.465 ;
        RECT 643.640 327.445 646.720 328.640 ;
        RECT 663.060 328.285 666.680 328.715 ;
        RECT 668.690 328.285 672.310 328.715 ;
        RECT 674.870 328.615 678.070 328.790 ;
        RECT 681.675 328.655 685.430 329.855 ;
        RECT 689.500 329.535 690.810 329.865 ;
        RECT 687.490 328.665 690.810 329.535 ;
        RECT 674.450 328.185 678.070 328.615 ;
        RECT 681.480 328.225 685.580 328.655 ;
        RECT 687.340 328.235 690.960 328.665 ;
        RECT 852.430 327.550 855.560 338.360 ;
        RECT 643.420 327.070 646.720 327.445 ;
        RECT 643.420 327.015 645.120 327.070 ;
        RECT 605.200 322.550 626.560 323.670 ;
        RECT 605.200 322.460 625.260 322.550 ;
        RECT 605.200 322.450 610.170 322.460 ;
        RECT 606.460 322.410 610.170 322.450 ;
        RECT 614.040 322.430 625.260 322.460 ;
        RECT 614.040 322.410 617.750 322.430 ;
        RECT 621.550 322.410 625.260 322.430 ;
        RECT 658.850 322.415 660.180 323.615 ;
        RECT 658.630 321.985 660.330 322.415 ;
        RECT 663.750 322.375 665.080 323.575 ;
        RECT 668.340 322.405 669.670 323.605 ;
        RECT 670.580 322.405 671.420 323.340 ;
        RECT 663.530 321.945 665.230 322.375 ;
        RECT 668.120 322.240 671.420 322.405 ;
        RECT 672.880 322.385 674.210 323.585 ;
        RECT 676.285 322.395 680.040 323.595 ;
        RECT 684.020 323.265 685.330 323.595 ;
        RECT 689.470 323.330 690.780 323.595 ;
        RECT 689.470 323.285 692.270 323.330 ;
        RECT 694.760 323.285 696.090 323.615 ;
        RECT 689.470 323.265 696.090 323.285 ;
        RECT 682.010 322.395 685.330 323.265 ;
        RECT 687.460 322.415 696.090 323.265 ;
        RECT 687.460 322.395 696.240 322.415 ;
        RECT 668.120 321.975 669.820 322.240 ;
        RECT 672.660 321.955 674.360 322.385 ;
        RECT 676.090 321.965 680.190 322.395 ;
        RECT 681.860 321.965 685.480 322.395 ;
        RECT 687.310 322.330 696.240 322.395 ;
        RECT 687.310 321.965 690.930 322.330 ;
        RECT 692.620 321.985 696.240 322.330 ;
        RECT 661.465 316.535 665.220 317.735 ;
        RECT 669.250 317.415 670.560 317.745 ;
        RECT 674.690 317.425 676.000 317.755 ;
        RECT 679.990 317.425 681.320 317.755 ;
        RECT 685.360 317.425 686.670 317.755 ;
        RECT 667.240 317.310 670.560 317.415 ;
        RECT 672.680 317.310 676.000 317.425 ;
        RECT 667.240 316.555 676.000 317.310 ;
        RECT 678.270 317.260 681.320 317.425 ;
        RECT 683.350 317.260 686.670 317.425 ;
        RECT 690.215 317.405 691.525 317.735 ;
        RECT 694.615 317.405 695.925 317.735 ;
        RECT 678.270 316.555 686.670 317.260 ;
        RECT 689.215 317.270 691.525 317.405 ;
        RECT 693.615 317.270 695.925 317.405 ;
        RECT 667.240 316.545 676.150 316.555 ;
        RECT 661.270 316.105 665.370 316.535 ;
        RECT 667.090 316.380 676.150 316.545 ;
        RECT 667.090 316.115 670.710 316.380 ;
        RECT 672.530 316.125 676.150 316.380 ;
        RECT 677.850 316.360 686.820 316.555 ;
        RECT 689.215 316.535 695.925 317.270 ;
        RECT 677.850 316.125 681.470 316.360 ;
        RECT 683.200 316.125 686.820 316.360 ;
        RECT 689.020 316.400 696.080 316.535 ;
        RECT 689.020 316.105 691.680 316.400 ;
        RECT 693.420 316.105 696.080 316.400 ;
        RECT 851.380 315.550 855.560 327.550 ;
        RECT 852.430 313.580 855.560 315.550 ;
        RECT 873.030 320.570 876.160 321.220 ;
        RECT 873.030 314.490 877.570 320.570 ;
        RECT 873.030 314.080 876.160 314.490 ;
        RECT 595.240 308.755 596.570 309.955 ;
        RECT 635.200 309.205 636.530 310.405 ;
        RECT 639.390 309.295 640.720 310.495 ;
        RECT 595.090 308.325 596.790 308.755 ;
        RECT 605.050 305.500 606.200 309.010 ;
        RECT 610.060 306.970 613.770 308.490 ;
        RECT 617.650 306.970 621.360 308.460 ;
        RECT 610.060 305.500 621.360 306.970 ;
        RECT 625.230 305.500 626.410 309.140 ;
        RECT 634.980 308.775 636.680 309.205 ;
        RECT 639.170 308.865 640.870 309.295 ;
        RECT 643.490 309.275 644.820 310.475 ;
        RECT 643.270 308.845 644.970 309.275 ;
        RECT 605.050 304.380 626.410 305.500 ;
        RECT 798.750 305.115 806.350 305.445 ;
        RECT 809.595 305.115 811.820 305.615 ;
        RECT 816.510 305.115 824.110 305.445 ;
        RECT 827.355 305.115 829.580 305.615 ;
        RECT 605.050 304.290 625.110 304.380 ;
        RECT 605.050 304.280 610.020 304.290 ;
        RECT 606.310 304.240 610.020 304.280 ;
        RECT 613.890 304.260 625.110 304.290 ;
        RECT 613.890 304.240 617.600 304.260 ;
        RECT 621.400 304.240 625.110 304.260 ;
        RECT 796.500 304.245 811.820 305.115 ;
        RECT 814.260 304.245 829.580 305.115 ;
        RECT 796.350 303.815 811.970 304.245 ;
        RECT 814.110 303.815 829.730 304.245 ;
        RECT 831.870 304.215 833.200 305.415 ;
        RECT 835.440 304.275 840.410 305.475 ;
        RECT 842.780 304.275 844.110 305.475 ;
        RECT 831.650 303.785 833.350 304.215 ;
        RECT 835.290 303.845 840.830 304.275 ;
        RECT 842.560 303.845 844.260 304.275 ;
        RECT 682.330 296.055 689.930 296.385 ;
        RECT 693.175 296.055 695.400 296.555 ;
        RECT 680.080 295.185 695.400 296.055 ;
        RECT 699.820 296.015 707.420 296.345 ;
        RECT 710.665 296.015 712.890 296.515 ;
        RECT 717.430 296.075 725.030 296.405 ;
        RECT 728.275 296.075 730.500 296.575 ;
        RECT 679.930 294.755 695.550 295.185 ;
        RECT 697.570 295.145 712.890 296.015 ;
        RECT 715.180 295.205 730.500 296.075 ;
        RECT 735.130 296.025 742.730 296.355 ;
        RECT 745.975 296.025 748.200 296.525 ;
        RECT 697.420 294.715 713.040 295.145 ;
        RECT 715.030 294.775 730.650 295.205 ;
        RECT 732.880 295.155 748.200 296.025 ;
        RECT 752.870 296.015 760.470 296.345 ;
        RECT 763.715 296.015 765.940 296.515 ;
        RECT 732.730 294.725 748.350 295.155 ;
        RECT 750.620 295.145 765.940 296.015 ;
        RECT 857.830 295.375 859.140 295.705 ;
        RECT 750.470 294.715 766.090 295.145 ;
        RECT 855.820 294.505 859.140 295.375 ;
        RECT 855.670 294.075 859.290 294.505 ;
        RECT 841.420 293.395 842.730 293.725 ;
        RECT 839.410 292.525 842.730 293.395 ;
        RECT 839.260 292.095 842.880 292.525 ;
        RECT 847.100 291.745 848.430 292.075 ;
        RECT 152.750 290.980 154.770 291.050 ;
        RECT 114.320 288.150 154.770 290.980 ;
        RECT 595.190 289.575 596.520 290.775 ;
        RECT 635.150 290.025 636.480 291.225 ;
        RECT 639.340 290.115 640.670 291.315 ;
        RECT 643.440 291.200 644.770 291.295 ;
        RECT 595.040 289.145 596.740 289.575 ;
        RECT 114.320 280.460 151.460 288.150 ;
        RECT 114.320 278.140 116.340 280.460 ;
        RECT 121.240 278.140 125.940 280.460 ;
        RECT 143.300 279.110 148.010 280.460 ;
        RECT 114.320 271.010 151.490 278.140 ;
        RECT 114.320 268.430 116.340 271.010 ;
        RECT 121.270 268.430 125.970 271.010 ;
        RECT 143.330 269.660 148.040 271.010 ;
        RECT 114.320 261.150 151.570 268.430 ;
        RECT 152.750 261.150 154.770 288.150 ;
        RECT 605.000 286.320 606.150 289.830 ;
        RECT 610.010 287.790 613.720 289.310 ;
        RECT 617.600 287.790 621.310 289.280 ;
        RECT 610.010 286.320 621.310 287.790 ;
        RECT 625.180 286.320 626.360 289.960 ;
        RECT 634.930 289.595 636.630 290.025 ;
        RECT 639.120 289.685 640.820 290.115 ;
        RECT 643.440 290.095 646.510 291.200 ;
        RECT 845.380 290.875 848.430 291.745 ;
        RECT 863.190 291.475 864.520 291.805 ;
        RECT 820.970 290.385 822.280 290.715 ;
        RECT 844.960 290.445 848.580 290.875 ;
        RECT 861.470 290.605 864.520 291.475 ;
        RECT 643.220 289.665 646.510 290.095 ;
        RECT 645.600 289.630 646.510 289.665 ;
        RECT 818.960 289.515 822.280 290.385 ;
        RECT 861.050 290.175 864.670 290.605 ;
        RECT 857.870 289.845 859.180 290.175 ;
        RECT 818.810 289.085 822.430 289.515 ;
        RECT 855.860 288.975 859.180 289.845 ;
        RECT 826.420 288.215 827.730 288.545 ;
        RECT 824.410 287.345 827.730 288.215 ;
        RECT 829.950 287.365 834.920 288.565 ;
        RECT 841.430 288.275 842.740 288.605 ;
        RECT 855.710 288.545 859.330 288.975 ;
        RECT 839.420 287.405 842.740 288.275 ;
        RECT 824.260 286.915 827.880 287.345 ;
        RECT 829.800 286.935 835.340 287.365 ;
        RECT 839.270 286.975 842.890 287.405 ;
        RECT 605.000 285.200 626.360 286.320 ;
        RECT 820.940 285.225 822.250 285.555 ;
        RECT 605.000 285.110 625.060 285.200 ;
        RECT 605.000 285.100 609.970 285.110 ;
        RECT 606.260 285.060 609.970 285.100 ;
        RECT 613.840 285.080 625.060 285.110 ;
        RECT 613.840 285.060 617.550 285.080 ;
        RECT 621.350 285.060 625.060 285.080 ;
        RECT 818.930 284.355 822.250 285.225 ;
        RECT 857.940 284.445 859.250 284.775 ;
        RECT 818.780 283.925 822.400 284.355 ;
        RECT 855.930 283.575 859.250 284.445 ;
        RECT 855.780 283.145 859.400 283.575 ;
        RECT 863.270 282.425 864.600 282.755 ;
        RECT 861.550 281.555 864.600 282.425 ;
        RECT 861.130 281.125 864.750 281.555 ;
        RECT 799.620 279.665 800.950 280.865 ;
        RECT 679.410 278.445 684.380 279.645 ;
        RECT 696.690 278.455 701.660 279.655 ;
        RECT 714.460 278.455 719.430 279.655 ;
        RECT 731.700 278.455 736.670 279.655 ;
        RECT 749.180 278.465 754.150 279.665 ;
        RECT 799.400 279.235 801.100 279.665 ;
        RECT 819.370 279.325 824.340 280.525 ;
        RECT 829.990 280.105 831.300 280.435 ;
        RECT 819.220 278.895 824.760 279.325 ;
        RECT 827.980 279.235 831.300 280.105 ;
        RECT 833.270 279.235 838.240 280.435 ;
        RECT 840.525 279.235 844.280 280.435 ;
        RECT 846.320 279.235 851.290 280.435 ;
        RECT 827.830 278.805 831.450 279.235 ;
        RECT 833.120 278.805 838.660 279.235 ;
        RECT 840.330 278.805 844.430 279.235 ;
        RECT 846.170 278.805 851.710 279.235 ;
        RECT 857.960 278.985 859.270 279.315 ;
        RECT 679.260 278.015 684.800 278.445 ;
        RECT 696.540 278.025 702.080 278.455 ;
        RECT 714.310 278.025 719.850 278.455 ;
        RECT 731.550 278.025 737.090 278.455 ;
        RECT 749.030 278.035 754.570 278.465 ;
        RECT 855.950 278.115 859.270 278.985 ;
        RECT 855.800 277.685 859.420 278.115 ;
        RECT 595.110 271.105 596.440 272.305 ;
        RECT 635.070 271.555 636.400 272.755 ;
        RECT 639.260 271.645 640.590 272.845 ;
        RECT 594.960 270.675 596.660 271.105 ;
        RECT 604.920 267.850 606.070 271.360 ;
        RECT 609.930 269.320 613.640 270.840 ;
        RECT 617.520 269.320 621.230 270.810 ;
        RECT 609.930 267.850 621.230 269.320 ;
        RECT 625.100 267.850 626.280 271.490 ;
        RECT 634.850 271.125 636.550 271.555 ;
        RECT 639.040 271.215 640.740 271.645 ;
        RECT 643.360 271.625 644.690 272.825 ;
        RECT 679.820 272.785 684.790 273.985 ;
        RECT 679.670 272.355 685.210 272.785 ;
        RECT 687.060 272.745 692.030 273.945 ;
        RECT 697.050 272.805 702.020 274.005 ;
        RECT 686.910 272.315 692.450 272.745 ;
        RECT 696.900 272.375 702.440 272.805 ;
        RECT 704.290 272.765 709.260 273.965 ;
        RECT 714.620 272.905 719.590 274.105 ;
        RECT 704.140 272.335 709.680 272.765 ;
        RECT 714.470 272.475 720.010 272.905 ;
        RECT 721.860 272.865 726.830 274.065 ;
        RECT 731.790 272.935 736.760 274.135 ;
        RECT 721.710 272.435 727.250 272.865 ;
        RECT 731.640 272.505 737.180 272.935 ;
        RECT 739.030 272.895 744.000 274.095 ;
        RECT 749.600 272.995 754.570 274.195 ;
        RECT 738.880 272.465 744.420 272.895 ;
        RECT 749.450 272.565 754.990 272.995 ;
        RECT 756.840 272.955 761.810 274.155 ;
        RECT 756.690 272.525 762.230 272.955 ;
        RECT 783.230 272.495 790.830 272.825 ;
        RECT 794.075 272.495 796.300 272.995 ;
        RECT 780.980 271.625 796.300 272.495 ;
        RECT 802.120 272.485 809.720 272.815 ;
        RECT 812.965 272.485 815.190 272.985 ;
        RECT 643.140 271.195 644.840 271.625 ;
        RECT 780.830 271.195 796.450 271.625 ;
        RECT 799.870 271.615 815.190 272.485 ;
        RECT 820.970 272.455 828.570 272.785 ;
        RECT 831.815 272.455 834.040 272.955 ;
        RECT 799.720 271.185 815.340 271.615 ;
        RECT 818.720 271.585 834.040 272.455 ;
        RECT 838.485 271.625 842.240 272.825 ;
        RECT 857.960 272.445 859.270 272.775 ;
        RECT 818.570 271.155 834.190 271.585 ;
        RECT 838.290 271.195 842.390 271.625 ;
        RECT 855.950 271.575 859.270 272.445 ;
        RECT 855.800 271.145 859.420 271.575 ;
        RECT 846.700 270.235 848.010 270.565 ;
        RECT 844.690 269.365 848.010 270.235 ;
        RECT 850.170 269.375 851.500 270.575 ;
        RECT 844.540 268.935 848.160 269.365 ;
        RECT 849.950 268.945 851.650 269.375 ;
        RECT 863.260 269.055 864.590 269.385 ;
        RECT 681.950 267.975 683.260 268.305 ;
        RECT 687.610 267.985 688.920 268.315 ;
        RECT 692.940 268.005 694.270 268.335 ;
        RECT 604.920 266.730 626.280 267.850 ;
        RECT 679.940 267.105 683.260 267.975 ;
        RECT 685.600 267.115 688.920 267.985 ;
        RECT 691.220 267.135 694.270 268.005 ;
        RECT 699.180 267.995 700.490 268.325 ;
        RECT 704.840 268.005 706.150 268.335 ;
        RECT 710.170 268.025 711.500 268.355 ;
        RECT 716.750 268.095 718.060 268.425 ;
        RECT 722.410 268.105 723.720 268.435 ;
        RECT 727.740 268.125 729.070 268.455 ;
        RECT 733.920 268.125 735.230 268.455 ;
        RECT 739.580 268.135 740.890 268.465 ;
        RECT 744.910 268.155 746.240 268.485 ;
        RECT 751.730 268.185 753.040 268.515 ;
        RECT 757.390 268.195 758.700 268.525 ;
        RECT 762.720 268.215 764.050 268.545 ;
        RECT 604.920 266.640 624.980 266.730 ;
        RECT 679.790 266.675 683.410 267.105 ;
        RECT 685.450 266.685 689.070 267.115 ;
        RECT 690.800 266.705 694.420 267.135 ;
        RECT 697.170 267.125 700.490 267.995 ;
        RECT 702.830 267.135 706.150 268.005 ;
        RECT 708.450 267.155 711.500 268.025 ;
        RECT 714.740 267.225 718.060 268.095 ;
        RECT 720.400 267.235 723.720 268.105 ;
        RECT 726.020 267.255 729.070 268.125 ;
        RECT 731.910 267.255 735.230 268.125 ;
        RECT 737.570 267.265 740.890 268.135 ;
        RECT 743.190 267.285 746.240 268.155 ;
        RECT 749.720 267.315 753.040 268.185 ;
        RECT 755.380 267.325 758.700 268.195 ;
        RECT 761.000 267.345 764.050 268.215 ;
        RECT 861.540 268.185 864.590 269.055 ;
        RECT 861.120 267.755 864.740 268.185 ;
        RECT 697.020 266.695 700.640 267.125 ;
        RECT 702.680 266.705 706.300 267.135 ;
        RECT 708.030 266.725 711.650 267.155 ;
        RECT 714.590 266.795 718.210 267.225 ;
        RECT 720.250 266.805 723.870 267.235 ;
        RECT 725.600 266.825 729.220 267.255 ;
        RECT 731.760 266.825 735.380 267.255 ;
        RECT 737.420 266.835 741.040 267.265 ;
        RECT 742.770 266.855 746.390 267.285 ;
        RECT 749.570 266.885 753.190 267.315 ;
        RECT 755.230 266.895 758.850 267.325 ;
        RECT 760.580 266.915 764.200 267.345 ;
        RECT 840.460 266.935 841.770 267.265 ;
        RECT 604.920 266.630 609.890 266.640 ;
        RECT 606.180 266.590 609.890 266.630 ;
        RECT 613.760 266.610 624.980 266.640 ;
        RECT 613.760 266.590 617.470 266.610 ;
        RECT 621.270 266.590 624.980 266.610 ;
        RECT 838.450 266.065 841.770 266.935 ;
        RECT 838.300 265.635 841.920 266.065 ;
        RECT 858.040 265.775 859.350 266.105 ;
        RECT 783.240 264.935 790.840 265.265 ;
        RECT 794.085 264.935 796.310 265.435 ;
        RECT 801.770 264.995 809.370 265.325 ;
        RECT 812.615 264.995 814.840 265.495 ;
        RECT 780.990 264.065 796.310 264.935 ;
        RECT 799.520 264.125 814.840 264.995 ;
        RECT 856.030 264.905 859.350 265.775 ;
        RECT 855.880 264.475 859.500 264.905 ;
        RECT 780.840 263.635 796.460 264.065 ;
        RECT 799.370 263.695 814.990 264.125 ;
        RECT 114.320 258.460 154.770 261.150 ;
        RECT 114.320 258.390 154.630 258.460 ;
        RECT 115.200 258.320 154.630 258.390 ;
        RECT 679.390 256.915 684.360 258.115 ;
        RECT 696.670 256.925 701.640 258.125 ;
        RECT 714.440 256.925 719.410 258.125 ;
        RECT 731.680 256.925 736.650 258.125 ;
        RECT 749.160 256.935 754.130 258.135 ;
        RECT 679.240 256.485 684.780 256.915 ;
        RECT 696.520 256.495 702.060 256.925 ;
        RECT 714.290 256.495 719.830 256.925 ;
        RECT 731.530 256.495 737.070 256.925 ;
        RECT 749.010 256.505 754.550 256.935 ;
        RECT 857.910 256.465 859.220 256.795 ;
        RECT 855.900 255.595 859.220 256.465 ;
        RECT 855.750 255.165 859.370 255.595 ;
        RECT 594.960 253.375 596.290 254.575 ;
        RECT 634.920 253.825 636.250 255.025 ;
        RECT 639.110 253.915 640.440 255.115 ;
        RECT 594.810 252.945 596.510 253.375 ;
        RECT 604.770 250.120 605.920 253.630 ;
        RECT 609.780 251.590 613.490 253.110 ;
        RECT 617.370 251.590 621.080 253.080 ;
        RECT 609.780 250.120 621.080 251.590 ;
        RECT 624.950 250.120 626.130 253.760 ;
        RECT 634.700 253.395 636.400 253.825 ;
        RECT 638.890 253.485 640.590 253.915 ;
        RECT 643.210 253.895 644.540 255.095 ;
        RECT 645.520 253.895 646.430 255.070 ;
        RECT 863.200 253.975 864.530 254.305 ;
        RECT 642.990 253.500 646.430 253.895 ;
        RECT 642.990 253.465 644.690 253.500 ;
        RECT 861.480 253.105 864.530 253.975 ;
        RECT 861.060 252.675 864.680 253.105 ;
        RECT 679.800 251.255 684.770 252.455 ;
        RECT 679.650 250.825 685.190 251.255 ;
        RECT 687.040 251.215 692.010 252.415 ;
        RECT 697.030 251.275 702.000 252.475 ;
        RECT 686.890 250.785 692.430 251.215 ;
        RECT 696.880 250.845 702.420 251.275 ;
        RECT 704.270 251.235 709.240 252.435 ;
        RECT 714.600 251.375 719.570 252.575 ;
        RECT 704.120 250.805 709.660 251.235 ;
        RECT 714.450 250.945 719.990 251.375 ;
        RECT 721.840 251.335 726.810 252.535 ;
        RECT 731.770 251.405 736.740 252.605 ;
        RECT 721.690 250.905 727.230 251.335 ;
        RECT 731.620 250.975 737.160 251.405 ;
        RECT 739.010 251.365 743.980 252.565 ;
        RECT 749.580 251.465 754.550 252.665 ;
        RECT 738.860 250.935 744.400 251.365 ;
        RECT 749.430 251.035 754.970 251.465 ;
        RECT 756.820 251.425 761.790 252.625 ;
        RECT 756.670 250.995 762.210 251.425 ;
        RECT 857.970 250.695 859.280 251.025 ;
        RECT 604.770 249.000 626.130 250.120 ;
        RECT 855.960 249.825 859.280 250.695 ;
        RECT 855.810 249.395 859.430 249.825 ;
        RECT 604.770 248.910 624.830 249.000 ;
        RECT 604.770 248.900 609.740 248.910 ;
        RECT 606.030 248.860 609.740 248.900 ;
        RECT 613.610 248.880 624.830 248.910 ;
        RECT 613.610 248.860 617.320 248.880 ;
        RECT 621.120 248.860 624.830 248.880 ;
        RECT 681.930 246.445 683.240 246.775 ;
        RECT 687.590 246.455 688.900 246.785 ;
        RECT 692.920 246.475 694.250 246.805 ;
        RECT 679.920 245.575 683.240 246.445 ;
        RECT 685.580 245.585 688.900 246.455 ;
        RECT 691.200 245.605 694.250 246.475 ;
        RECT 699.160 246.465 700.470 246.795 ;
        RECT 704.820 246.475 706.130 246.805 ;
        RECT 710.150 246.495 711.480 246.825 ;
        RECT 716.730 246.565 718.040 246.895 ;
        RECT 722.390 246.575 723.700 246.905 ;
        RECT 727.720 246.595 729.050 246.925 ;
        RECT 733.900 246.595 735.210 246.925 ;
        RECT 739.560 246.605 740.870 246.935 ;
        RECT 744.890 246.625 746.220 246.955 ;
        RECT 751.710 246.655 753.020 246.985 ;
        RECT 757.370 246.665 758.680 246.995 ;
        RECT 762.700 246.685 764.030 247.015 ;
        RECT 679.770 245.145 683.390 245.575 ;
        RECT 685.430 245.155 689.050 245.585 ;
        RECT 690.780 245.175 694.400 245.605 ;
        RECT 697.150 245.595 700.470 246.465 ;
        RECT 702.810 245.605 706.130 246.475 ;
        RECT 708.430 245.625 711.480 246.495 ;
        RECT 714.720 245.695 718.040 246.565 ;
        RECT 720.380 245.705 723.700 246.575 ;
        RECT 726.000 245.725 729.050 246.595 ;
        RECT 731.890 245.725 735.210 246.595 ;
        RECT 737.550 245.735 740.870 246.605 ;
        RECT 743.170 245.755 746.220 246.625 ;
        RECT 749.700 245.785 753.020 246.655 ;
        RECT 755.360 245.795 758.680 246.665 ;
        RECT 760.980 245.815 764.030 246.685 ;
        RECT 697.000 245.165 700.620 245.595 ;
        RECT 702.660 245.175 706.280 245.605 ;
        RECT 708.010 245.195 711.630 245.625 ;
        RECT 714.570 245.265 718.190 245.695 ;
        RECT 720.230 245.275 723.850 245.705 ;
        RECT 725.580 245.295 729.200 245.725 ;
        RECT 731.740 245.295 735.360 245.725 ;
        RECT 737.400 245.305 741.020 245.735 ;
        RECT 742.750 245.325 746.370 245.755 ;
        RECT 749.550 245.355 753.170 245.785 ;
        RECT 755.210 245.365 758.830 245.795 ;
        RECT 760.560 245.385 764.180 245.815 ;
        RECT -98.710 230.000 -71.020 237.170 ;
        RECT -0.130 227.160 301.170 227.290 ;
        RECT -98.020 217.900 -70.330 225.070 ;
        RECT -0.130 220.340 301.320 227.160 ;
        RECT -98.420 130.150 -70.730 137.320 ;
        RECT -97.990 10.820 -70.300 17.990 ;
        RECT 0.110 6.550 8.640 220.340 ;
        RECT 297.660 217.450 301.320 220.340 ;
        RECT 309.970 218.590 369.870 220.330 ;
        RECT 42.170 211.080 69.170 217.200 ;
        RECT 172.310 214.240 199.310 217.270 ;
        RECT 37.850 190.060 69.170 211.080 ;
        RECT 71.370 208.580 72.670 208.610 ;
        RECT 37.850 188.120 41.390 190.060 ;
        RECT 37.850 160.980 69.170 188.120 ;
        RECT 37.850 158.950 41.390 160.980 ;
        RECT 37.850 131.810 69.170 158.950 ;
        RECT 37.850 129.770 41.390 131.810 ;
        RECT 37.850 102.630 69.170 129.770 ;
        RECT 37.850 100.450 41.390 102.630 ;
        RECT 37.850 73.310 69.170 100.450 ;
        RECT 37.850 71.170 41.390 73.310 ;
        RECT 37.850 44.030 69.220 71.170 ;
        RECT 37.850 24.730 41.390 44.030 ;
        RECT 70.100 41.630 73.560 208.580 ;
        RECT 102.670 41.670 106.130 209.600 ;
        RECT 38.980 24.130 40.280 24.730 ;
        RECT 42.310 16.760 73.560 41.630 ;
        RECT 74.840 17.780 106.130 41.670 ;
        RECT 42.310 14.490 69.310 16.760 ;
        RECT 74.840 14.530 101.840 17.780 ;
        RECT 135.280 17.520 138.570 213.980 ;
        RECT 167.820 190.130 199.310 214.240 ;
        RECT 167.820 188.190 171.520 190.130 ;
        RECT 167.820 161.050 199.310 188.190 ;
        RECT 167.820 159.020 171.520 161.050 ;
        RECT 167.820 131.880 199.310 159.020 ;
        RECT 167.820 129.840 171.520 131.880 ;
        RECT 167.820 102.700 199.310 129.840 ;
        RECT 167.820 100.520 171.520 102.700 ;
        RECT 167.820 73.380 199.310 100.520 ;
        RECT 167.820 71.240 171.520 73.380 ;
        RECT 167.820 44.100 199.360 71.240 ;
        RECT 167.820 18.810 171.520 44.100 ;
        RECT 200.330 27.810 203.820 212.960 ;
        RECT 201.570 24.200 202.870 27.810 ;
        RECT 232.850 26.900 236.590 212.250 ;
        RECT 265.550 71.350 269.290 212.100 ;
        RECT 270.270 190.310 301.320 217.450 ;
        RECT 310.230 216.740 312.160 218.590 ;
        RECT 367.830 216.820 369.860 218.590 ;
        RECT 310.230 213.640 329.350 216.740 ;
        RECT 331.320 213.710 348.320 216.750 ;
        RECT 350.360 215.140 369.860 216.820 ;
        RECT 350.360 213.710 369.880 215.140 ;
        RECT 331.320 213.640 369.880 213.710 ;
        RECT 310.230 203.900 369.880 213.640 ;
        RECT 310.230 203.830 348.320 203.900 ;
        RECT 310.230 199.600 329.350 203.830 ;
        RECT 331.320 199.610 348.320 203.830 ;
        RECT 350.360 203.210 369.880 203.900 ;
        RECT 350.360 199.680 369.860 203.210 ;
        RECT 310.230 198.450 312.160 199.600 ;
        RECT 367.830 198.450 369.860 199.680 ;
        RECT 310.190 196.930 369.860 198.450 ;
        RECT 382.570 198.400 435.910 200.330 ;
        RECT 382.490 197.850 435.910 198.400 ;
        RECT 310.190 196.580 369.650 196.930 ;
        RECT 382.490 196.670 385.190 197.850 ;
        RECT 297.660 188.370 301.320 190.310 ;
        RECT 270.270 161.230 301.320 188.370 ;
        RECT 382.490 195.510 399.370 196.670 ;
        RECT 432.980 196.640 435.680 197.850 ;
        RECT 402.290 195.510 416.000 196.640 ;
        RECT 418.840 195.510 435.680 196.640 ;
        RECT 382.490 177.490 435.680 195.510 ;
        RECT 382.490 176.060 399.370 177.490 ;
        RECT 382.490 175.010 385.190 176.060 ;
        RECT 402.290 176.030 416.000 177.490 ;
        RECT 418.840 176.030 435.680 177.490 ;
        RECT 432.760 175.120 435.680 176.030 ;
        RECT 432.760 175.010 435.610 175.120 ;
        RECT 382.490 173.270 435.610 175.010 ;
        RECT 382.940 173.190 435.610 173.270 ;
        RECT 432.760 173.050 435.610 173.190 ;
        RECT 297.660 159.200 301.320 161.230 ;
        RECT 270.270 132.060 301.320 159.200 ;
        RECT 304.160 137.810 309.830 137.950 ;
        RECT 304.160 134.480 507.050 137.810 ;
        RECT 304.160 133.870 507.390 134.480 ;
        RECT 304.160 132.070 309.830 133.870 ;
        RECT 297.660 130.020 301.320 132.060 ;
        RECT 270.270 102.880 301.320 130.020 ;
        RECT 297.660 100.700 301.320 102.880 ;
        RECT 270.270 73.560 301.320 100.700 ;
        RECT 297.660 71.420 301.320 73.560 ;
        RECT 237.750 44.210 269.290 71.350 ;
        RECT 270.320 44.280 301.320 71.420 ;
        RECT 265.550 41.810 269.290 44.210 ;
        RECT 297.660 41.880 301.320 44.280 ;
        RECT 234.510 24.310 235.810 26.900 ;
        RECT 237.840 26.750 269.290 41.810 ;
        RECT 237.840 14.670 264.840 26.750 ;
        RECT 267.080 24.380 268.380 26.750 ;
        RECT 270.410 14.740 301.320 41.880 ;
        RECT 297.660 6.550 301.320 14.740 ;
        RECT 304.480 129.740 309.810 132.070 ;
        RECT 304.480 102.600 337.370 129.740 ;
        RECT 304.480 100.550 309.810 102.600 ;
        RECT 304.480 73.410 337.400 100.550 ;
        RECT 304.480 71.260 309.810 73.410 ;
        RECT 304.480 44.120 337.400 71.260 ;
        RECT 304.480 41.970 309.810 44.120 ;
        RECT 304.480 14.830 337.400 41.970 ;
        RECT 338.330 23.830 341.750 126.940 ;
        RECT 376.150 124.880 403.150 129.600 ;
        RECT 408.460 124.880 435.460 129.590 ;
        RECT 502.060 129.550 507.390 133.870 ;
        RECT 437.970 125.650 441.250 125.660 ;
        RECT 376.150 124.540 435.460 124.880 ;
        RECT 371.270 102.460 435.460 124.540 ;
        RECT 371.270 100.410 375.460 102.460 ;
        RECT 403.460 102.450 435.460 102.460 ;
        RECT 403.460 100.410 407.650 102.450 ;
        RECT 371.270 73.270 407.650 100.410 ;
        RECT 371.270 71.120 375.460 73.270 ;
        RECT 403.460 71.120 407.650 73.270 ;
        RECT 371.270 43.980 407.650 71.120 ;
        RECT 371.270 41.830 375.460 43.980 ;
        RECT 403.460 41.830 407.650 43.980 ;
        RECT 371.270 17.270 407.650 41.830 ;
        RECT 436.690 18.060 441.250 125.650 ;
        RECT 470.250 21.080 473.530 125.140 ;
        RECT 474.630 102.410 507.390 129.550 ;
        RECT 502.060 100.430 507.390 102.410 ;
        RECT 474.670 73.290 507.390 100.430 ;
        RECT 502.060 71.070 507.390 73.290 ;
        RECT 474.690 43.930 507.390 71.070 ;
        RECT 502.060 41.780 507.390 43.930 ;
        RECT 436.690 17.710 439.490 18.060 ;
        RECT 371.270 16.930 403.180 17.270 ;
        RECT 304.480 13.030 309.810 14.830 ;
        RECT 376.180 14.690 403.180 16.930 ;
        RECT 474.710 14.640 507.390 41.780 ;
        RECT 502.060 13.030 507.390 14.640 ;
        RECT 304.410 11.920 507.390 13.030 ;
        RECT 304.410 9.090 507.300 11.920 ;
        RECT 0.110 0.020 301.590 6.550 ;
        RECT 297.660 -0.130 301.320 0.020 ;
      LAYER li1 ;
        RECT -91.040 358.010 -77.710 358.180 ;
        RECT -98.030 353.245 -97.860 356.325 ;
        RECT -97.360 354.130 -97.190 355.750 ;
        RECT -94.780 354.130 -94.610 355.750 ;
        RECT -92.200 354.130 -92.030 355.750 ;
        RECT -89.620 354.130 -89.450 355.750 ;
        RECT -87.040 354.130 -86.870 355.750 ;
        RECT -84.460 354.130 -84.290 355.750 ;
        RECT -81.880 354.130 -81.710 355.750 ;
        RECT -79.300 354.130 -79.130 355.750 ;
        RECT -76.720 354.130 -76.550 355.750 ;
        RECT -74.140 354.130 -73.970 355.750 ;
        RECT -71.560 354.130 -71.390 355.750 ;
        RECT -70.890 353.245 -70.720 356.325 ;
        RECT -96.585 352.250 -72.085 352.285 ;
        RECT -96.920 352.080 -71.830 352.250 ;
        RECT -96.585 352.035 -72.085 352.080 ;
        RECT -81.845 351.750 -81.675 352.035 ;
        RECT -90.980 351.560 -77.510 351.750 ;
        RECT -91.040 351.390 -77.510 351.560 ;
        RECT -90.980 349.630 -77.510 351.390 ;
        RECT 654.730 351.225 655.320 352.185 ;
        RECT 658.225 351.215 659.175 352.345 ;
        RECT 660.830 351.215 661.780 351.765 ;
        RECT 664.800 351.215 665.750 351.795 ;
        RECT 670.120 351.215 670.710 352.095 ;
        RECT 671.400 351.215 672.350 351.845 ;
        RECT 676.275 351.175 677.225 352.305 ;
        RECT 678.880 351.175 679.830 351.725 ;
        RECT 682.850 351.175 683.800 351.755 ;
        RECT 688.170 351.175 688.760 352.055 ;
        RECT 689.450 351.175 690.400 351.805 ;
        RECT 693.865 351.195 694.815 352.325 ;
        RECT 696.470 351.195 697.420 351.745 ;
        RECT 700.440 351.195 701.390 351.775 ;
        RECT 705.760 351.195 706.350 352.075 ;
        RECT 707.040 351.195 707.990 351.825 ;
        RECT 711.715 351.195 712.665 352.325 ;
        RECT 714.320 351.195 715.270 351.745 ;
        RECT 718.290 351.195 719.240 351.775 ;
        RECT 723.610 351.195 724.200 352.075 ;
        RECT 724.890 351.195 725.840 351.825 ;
        RECT 729.975 351.195 730.925 352.325 ;
        RECT 732.580 351.195 733.530 351.745 ;
        RECT 736.550 351.195 737.500 351.775 ;
        RECT 741.870 351.195 742.460 352.075 ;
        RECT 743.150 351.195 744.100 351.825 ;
        RECT 747.745 351.165 748.695 352.295 ;
        RECT 750.350 351.165 751.300 351.715 ;
        RECT 754.320 351.165 755.270 351.745 ;
        RECT 759.640 351.165 760.230 352.045 ;
        RECT 760.920 351.165 761.870 351.795 ;
        RECT 765.785 351.085 766.735 352.215 ;
        RECT 768.390 351.085 769.340 351.635 ;
        RECT 772.360 351.085 773.310 351.665 ;
        RECT 777.680 351.085 778.270 351.965 ;
        RECT 778.960 351.085 779.910 351.715 ;
        RECT 783.945 351.125 784.895 352.255 ;
        RECT 786.550 351.125 787.500 351.675 ;
        RECT 790.520 351.125 791.470 351.705 ;
        RECT 795.840 351.125 796.430 352.005 ;
        RECT 797.120 351.125 798.070 351.755 ;
        RECT 802.325 351.135 803.275 352.265 ;
        RECT 804.930 351.135 805.880 351.685 ;
        RECT 808.900 351.135 809.850 351.715 ;
        RECT 814.220 351.135 814.810 352.015 ;
        RECT 815.500 351.135 816.450 351.765 ;
        RECT 821.125 351.115 822.075 352.245 ;
        RECT 823.730 351.115 824.680 351.665 ;
        RECT 827.700 351.115 828.650 351.695 ;
        RECT 833.020 351.115 833.610 351.995 ;
        RECT 834.300 351.115 835.250 351.745 ;
        RECT 839.680 351.095 840.270 352.055 ;
        RECT 653.970 350.775 655.410 350.945 ;
        RECT 657.550 350.765 672.910 350.935 ;
        RECT 675.600 350.725 690.960 350.895 ;
        RECT 693.190 350.745 708.550 350.915 ;
        RECT 711.040 350.745 726.400 350.915 ;
        RECT 729.300 350.745 744.660 350.915 ;
        RECT 747.070 350.715 762.430 350.885 ;
        RECT 765.110 350.635 780.470 350.805 ;
        RECT 783.270 350.675 798.630 350.845 ;
        RECT 801.650 350.685 817.010 350.855 ;
        RECT 820.450 350.665 835.810 350.835 ;
        RECT 838.920 350.645 840.360 350.815 ;
        RECT 784.565 342.955 785.555 343.915 ;
        RECT 791.150 342.985 791.740 343.945 ;
        RECT 794.525 343.045 795.475 344.175 ;
        RECT 797.130 343.045 798.080 343.595 ;
        RECT 801.100 343.045 802.050 343.625 ;
        RECT 806.420 343.045 807.010 343.925 ;
        RECT 807.700 343.045 808.650 343.675 ;
        RECT 813.885 342.955 814.835 344.085 ;
        RECT 816.490 342.955 817.440 343.505 ;
        RECT 820.460 342.955 821.410 343.535 ;
        RECT 825.780 342.955 826.370 343.835 ;
        RECT 827.060 342.955 828.010 343.585 ;
        RECT 783.830 342.505 787.190 342.675 ;
        RECT 790.390 342.535 791.830 342.705 ;
        RECT 793.850 342.595 809.210 342.765 ;
        RECT 813.210 342.505 828.570 342.675 ;
        RECT 853.910 337.520 854.080 337.940 ;
        RECT 853.910 336.050 854.080 336.470 ;
        RECT 853.910 334.580 854.080 335.000 ;
        RECT 853.910 333.110 854.080 333.530 ;
        RECT 853.910 331.640 854.080 332.060 ;
        RECT 853.910 330.170 854.080 330.590 ;
        RECT 664.825 328.865 665.815 329.825 ;
        RECT 670.455 328.865 671.445 329.825 ;
        RECT 674.670 328.765 675.580 329.395 ;
        RECT 676.620 328.765 677.210 329.725 ;
        RECT 678.350 328.920 679.130 329.690 ;
        RECT 684.045 328.805 684.850 329.765 ;
        RECT 689.105 328.815 690.095 329.775 ;
        RECT 853.910 328.700 854.080 329.120 ;
        RECT 596.130 327.075 596.720 328.035 ;
        RECT 635.350 327.525 635.940 328.485 ;
        RECT 639.540 327.615 640.130 328.575 ;
        RECT 643.640 327.595 644.230 328.555 ;
        RECT 595.370 326.625 596.810 326.795 ;
        RECT 596.610 325.840 597.180 326.140 ;
        RECT 605.330 322.580 606.220 327.050 ;
        RECT 615.020 324.300 615.190 324.720 ;
        RECT 616.600 324.300 616.770 324.720 ;
        RECT 615.020 322.830 615.190 323.250 ;
        RECT 616.600 322.830 616.770 323.250 ;
        RECT 625.510 322.680 626.430 327.180 ;
        RECT 635.260 327.075 636.700 327.245 ;
        RECT 639.450 327.165 640.890 327.335 ;
        RECT 643.550 327.145 644.990 327.315 ;
        RECT 645.940 327.200 646.590 328.510 ;
        RECT 663.190 328.415 666.550 328.585 ;
        RECT 668.820 328.415 672.180 328.585 ;
        RECT 674.580 328.315 677.940 328.485 ;
        RECT 681.610 328.355 685.450 328.525 ;
        RECT 687.470 328.365 690.830 328.535 ;
        RECT 640.370 323.410 640.540 323.830 ;
        RECT 644.420 323.460 644.590 323.880 ;
        RECT 658.850 322.565 659.440 323.525 ;
        RECT 663.750 322.525 664.340 323.485 ;
        RECT 668.340 322.555 668.930 323.515 ;
        RECT 670.710 322.370 671.290 323.210 ;
        RECT 672.880 322.535 673.470 323.495 ;
        RECT 678.655 322.545 679.460 323.505 ;
        RECT 683.625 322.545 684.615 323.505 ;
        RECT 689.075 322.545 690.065 323.505 ;
        RECT 691.410 322.460 692.140 323.200 ;
        RECT 692.840 322.565 693.750 323.195 ;
        RECT 694.790 322.565 695.380 323.525 ;
        RECT 658.760 322.115 660.200 322.285 ;
        RECT 663.660 322.075 665.100 322.245 ;
        RECT 668.250 322.105 669.690 322.275 ;
        RECT 672.790 322.085 674.230 322.255 ;
        RECT 676.220 322.095 680.060 322.265 ;
        RECT 681.990 322.095 685.350 322.265 ;
        RECT 687.440 322.095 690.800 322.265 ;
        RECT 692.750 322.115 696.110 322.285 ;
        RECT 663.835 316.685 664.640 317.645 ;
        RECT 668.855 316.695 669.845 317.655 ;
        RECT 671.050 316.510 671.780 317.180 ;
        RECT 674.295 316.705 675.285 317.665 ;
        RECT 678.070 316.705 678.980 317.335 ;
        RECT 680.020 316.705 680.610 317.665 ;
        RECT 681.900 316.490 682.670 317.130 ;
        RECT 684.965 316.705 685.955 317.665 ;
        RECT 689.755 316.685 691.005 317.255 ;
        RECT 692.160 316.530 693.000 317.140 ;
        RECT 694.155 316.685 695.405 317.255 ;
        RECT 661.400 316.235 665.240 316.405 ;
        RECT 667.220 316.245 670.580 316.415 ;
        RECT 672.660 316.255 676.020 316.425 ;
        RECT 677.980 316.255 681.340 316.425 ;
        RECT 683.330 316.255 686.690 316.425 ;
        RECT 689.150 316.235 691.550 316.405 ;
        RECT 693.550 316.235 695.950 316.405 ;
        RECT 851.510 315.680 852.180 327.420 ;
        RECT 853.910 327.230 854.080 327.650 ;
        RECT 853.910 325.760 854.080 326.180 ;
        RECT 853.910 324.290 854.080 324.710 ;
        RECT 853.910 322.820 854.080 323.240 ;
        RECT 853.910 321.350 854.080 321.770 ;
        RECT 874.510 320.380 874.680 320.800 ;
        RECT 853.910 319.880 854.080 320.300 ;
        RECT 874.510 318.910 874.680 319.330 ;
        RECT 853.910 318.410 854.080 318.830 ;
        RECT 874.510 317.440 874.680 317.860 ;
        RECT 853.910 316.940 854.080 317.360 ;
        RECT 874.510 315.970 874.680 316.390 ;
        RECT 853.910 315.470 854.080 315.890 ;
        RECT 874.510 314.500 874.680 314.920 ;
        RECT 876.590 314.620 877.440 320.440 ;
        RECT 853.910 314.000 854.080 314.420 ;
        RECT 595.980 308.905 596.570 309.865 ;
        RECT 635.200 309.355 635.790 310.315 ;
        RECT 639.390 309.445 639.980 310.405 ;
        RECT 643.490 309.425 644.080 310.385 ;
        RECT 595.220 308.455 596.660 308.625 ;
        RECT 596.460 307.670 597.030 307.970 ;
        RECT 605.180 304.410 606.070 308.880 ;
        RECT 614.870 306.130 615.040 306.550 ;
        RECT 616.450 306.130 616.620 306.550 ;
        RECT 614.870 304.660 615.040 305.080 ;
        RECT 616.450 304.660 616.620 305.080 ;
        RECT 625.360 304.510 626.280 309.010 ;
        RECT 635.110 308.905 636.550 309.075 ;
        RECT 639.300 308.995 640.740 309.165 ;
        RECT 643.400 308.975 644.840 309.145 ;
        RECT 640.220 305.240 640.390 305.660 ;
        RECT 644.270 305.290 644.440 305.710 ;
        RECT 797.040 304.395 797.990 305.025 ;
        RECT 798.680 304.395 799.270 305.275 ;
        RECT 803.640 304.395 804.590 304.975 ;
        RECT 807.610 304.395 808.560 304.945 ;
        RECT 810.215 304.395 811.165 305.525 ;
        RECT 814.800 304.395 815.750 305.025 ;
        RECT 816.440 304.395 817.030 305.275 ;
        RECT 821.400 304.395 822.350 304.975 ;
        RECT 825.370 304.395 826.320 304.945 ;
        RECT 827.975 304.395 828.925 305.525 ;
        RECT 831.870 304.365 832.460 305.325 ;
        RECT 835.510 304.425 836.100 305.305 ;
        RECT 836.760 304.425 839.090 305.305 ;
        RECT 839.970 304.425 840.560 305.385 ;
        RECT 842.780 304.425 843.370 305.385 ;
        RECT 796.480 303.945 811.840 304.115 ;
        RECT 814.240 303.945 829.600 304.115 ;
        RECT 831.780 303.915 833.220 304.085 ;
        RECT 835.420 303.975 840.700 304.145 ;
        RECT 842.690 303.975 844.130 304.145 ;
        RECT 680.620 295.335 681.570 295.965 ;
        RECT 682.260 295.335 682.850 296.215 ;
        RECT 687.220 295.335 688.170 295.915 ;
        RECT 691.190 295.335 692.140 295.885 ;
        RECT 693.795 295.335 694.745 296.465 ;
        RECT 698.110 295.295 699.060 295.925 ;
        RECT 699.750 295.295 700.340 296.175 ;
        RECT 704.710 295.295 705.660 295.875 ;
        RECT 708.680 295.295 709.630 295.845 ;
        RECT 711.285 295.295 712.235 296.425 ;
        RECT 715.720 295.355 716.670 295.985 ;
        RECT 717.360 295.355 717.950 296.235 ;
        RECT 722.320 295.355 723.270 295.935 ;
        RECT 726.290 295.355 727.240 295.905 ;
        RECT 728.895 295.355 729.845 296.485 ;
        RECT 733.420 295.305 734.370 295.935 ;
        RECT 735.060 295.305 735.650 296.185 ;
        RECT 740.020 295.305 740.970 295.885 ;
        RECT 743.990 295.305 744.940 295.855 ;
        RECT 746.595 295.305 747.545 296.435 ;
        RECT 751.160 295.295 752.110 295.925 ;
        RECT 752.800 295.295 753.390 296.175 ;
        RECT 757.760 295.295 758.710 295.875 ;
        RECT 761.730 295.295 762.680 295.845 ;
        RECT 764.335 295.295 765.285 296.425 ;
        RECT 680.060 294.885 695.420 295.055 ;
        RECT 697.550 294.845 712.910 295.015 ;
        RECT 715.160 294.905 730.520 295.075 ;
        RECT 732.860 294.855 748.220 295.025 ;
        RECT 750.600 294.845 765.960 295.015 ;
        RECT 857.435 294.655 858.425 295.615 ;
        RECT 855.800 294.205 859.160 294.375 ;
        RECT 841.025 292.675 842.015 293.635 ;
        RECT 839.390 292.225 842.750 292.395 ;
        RECT 595.930 289.725 596.520 290.685 ;
        RECT 635.150 290.175 635.740 291.135 ;
        RECT 639.340 290.265 639.930 291.225 ;
        RECT 643.440 290.245 644.030 291.205 ;
        RECT 595.170 289.275 596.610 289.445 ;
        RECT 596.410 288.490 596.980 288.790 ;
        RECT 150.750 287.440 151.030 287.460 ;
        RECT 150.110 287.430 151.040 287.440 ;
        RECT 118.630 287.400 151.040 287.430 ;
        RECT 118.090 287.230 151.040 287.400 ;
        RECT 118.630 287.160 151.040 287.230 ;
        RECT 118.630 287.120 150.200 287.160 ;
        RECT 150.750 284.160 151.030 287.160 ;
        RECT 605.130 285.230 606.020 289.700 ;
        RECT 614.820 286.950 614.990 287.370 ;
        RECT 616.400 286.950 616.570 287.370 ;
        RECT 614.820 285.480 614.990 285.900 ;
        RECT 616.400 285.480 616.570 285.900 ;
        RECT 625.310 285.330 626.230 289.830 ;
        RECT 635.060 289.725 636.500 289.895 ;
        RECT 639.250 289.815 640.690 289.985 ;
        RECT 643.350 289.795 644.790 289.965 ;
        RECT 645.730 289.760 646.380 291.070 ;
        RECT 845.180 291.025 846.090 291.655 ;
        RECT 847.130 291.025 847.720 291.985 ;
        RECT 861.270 290.755 862.180 291.385 ;
        RECT 863.220 290.755 863.810 291.715 ;
        RECT 820.575 289.665 821.565 290.625 ;
        RECT 845.090 290.575 848.450 290.745 ;
        RECT 861.180 290.305 864.540 290.475 ;
        RECT 818.940 289.215 822.300 289.385 ;
        RECT 857.475 289.125 858.465 290.085 ;
        RECT 855.840 288.675 859.200 288.845 ;
        RECT 826.025 287.495 827.015 288.455 ;
        RECT 830.020 287.515 830.610 288.395 ;
        RECT 831.270 287.515 833.600 288.395 ;
        RECT 834.480 287.515 835.070 288.475 ;
        RECT 841.035 287.555 842.025 288.515 ;
        RECT 824.390 287.045 827.750 287.215 ;
        RECT 829.930 287.065 835.210 287.235 ;
        RECT 839.400 287.105 842.760 287.275 ;
        RECT 640.170 286.060 640.340 286.480 ;
        RECT 644.220 286.110 644.390 286.530 ;
        RECT 820.545 284.505 821.535 285.465 ;
        RECT 151.610 284.160 152.080 284.350 ;
        RECT 117.410 284.150 118.800 284.160 ;
        RECT 150.750 284.150 152.080 284.160 ;
        RECT 117.410 283.950 152.080 284.150 ;
        RECT 818.910 284.055 822.270 284.225 ;
        RECT 117.410 283.940 151.150 283.950 ;
        RECT 117.410 283.840 150.210 283.940 ;
        RECT 117.410 283.820 118.800 283.840 ;
        RECT 150.750 280.900 151.030 283.940 ;
        RECT 151.610 283.750 152.080 283.950 ;
        RECT 857.545 283.725 858.535 284.685 ;
        RECT 855.910 283.275 859.270 283.445 ;
        RECT 861.350 281.705 862.260 282.335 ;
        RECT 863.300 281.705 863.890 282.665 ;
        RECT 861.260 281.255 864.620 281.425 ;
        RECT 149.970 280.880 151.030 280.900 ;
        RECT 118.530 280.820 151.030 280.880 ;
        RECT 118.090 280.650 151.030 280.820 ;
        RECT 118.530 280.600 151.030 280.650 ;
        RECT 118.530 280.590 151.010 280.600 ;
        RECT 118.530 280.570 150.100 280.590 ;
        RECT 147.030 279.950 147.670 280.570 ;
        RECT 121.370 278.660 125.810 279.540 ;
        RECT 143.430 279.240 147.880 279.950 ;
        RECT 799.620 279.815 800.210 280.775 ;
        RECT 679.480 278.595 680.070 279.475 ;
        RECT 680.730 278.595 683.060 279.475 ;
        RECT 683.940 278.595 684.530 279.555 ;
        RECT 696.760 278.605 697.350 279.485 ;
        RECT 698.010 278.605 700.340 279.485 ;
        RECT 701.220 278.605 701.810 279.565 ;
        RECT 714.530 278.605 715.120 279.485 ;
        RECT 715.780 278.605 718.110 279.485 ;
        RECT 718.990 278.605 719.580 279.565 ;
        RECT 731.770 278.605 732.360 279.485 ;
        RECT 733.020 278.605 735.350 279.485 ;
        RECT 736.230 278.605 736.820 279.565 ;
        RECT 749.250 278.615 749.840 279.495 ;
        RECT 750.500 278.615 752.830 279.495 ;
        RECT 753.710 278.615 754.300 279.575 ;
        RECT 799.530 279.365 800.970 279.535 ;
        RECT 819.440 279.475 820.030 280.355 ;
        RECT 820.690 279.475 823.020 280.355 ;
        RECT 823.900 279.475 824.490 280.435 ;
        RECT 829.595 279.385 830.585 280.345 ;
        RECT 833.340 279.385 833.930 280.265 ;
        RECT 834.590 279.385 836.920 280.265 ;
        RECT 837.800 279.385 838.390 280.345 ;
        RECT 842.895 279.385 843.700 280.345 ;
        RECT 846.390 279.385 846.980 280.265 ;
        RECT 847.640 279.385 849.970 280.265 ;
        RECT 850.850 279.385 851.440 280.345 ;
        RECT 819.350 279.025 824.630 279.195 ;
        RECT 827.960 278.935 831.320 279.105 ;
        RECT 833.250 278.935 838.530 279.105 ;
        RECT 840.460 278.935 844.300 279.105 ;
        RECT 846.300 278.935 851.580 279.105 ;
        RECT 679.390 278.145 684.670 278.315 ;
        RECT 696.670 278.155 701.950 278.325 ;
        RECT 714.440 278.155 719.720 278.325 ;
        RECT 731.680 278.155 736.960 278.325 ;
        RECT 749.160 278.165 754.440 278.335 ;
        RECT 857.565 278.265 858.555 279.225 ;
        RECT 855.930 277.815 859.290 277.985 ;
        RECT 114.580 275.350 116.010 276.880 ;
        RECT 114.580 274.870 117.420 275.350 ;
        RECT 114.580 274.710 117.690 274.870 ;
        RECT 114.580 274.700 118.830 274.710 ;
        RECT 114.580 274.660 150.240 274.700 ;
        RECT 114.580 274.490 150.370 274.660 ;
        RECT 751.625 274.555 752.815 274.930 ;
        RECT 114.580 274.460 150.240 274.490 ;
        RECT 114.580 274.300 116.010 274.460 ;
        RECT 116.580 274.390 150.240 274.460 ;
        RECT 116.580 274.370 118.830 274.390 ;
        RECT 116.580 274.220 117.690 274.370 ;
        RECT 679.890 272.935 680.480 273.815 ;
        RECT 681.140 272.935 683.470 273.815 ;
        RECT 684.350 272.935 684.940 273.895 ;
        RECT 687.130 272.895 687.720 273.775 ;
        RECT 688.380 272.895 690.710 273.775 ;
        RECT 691.590 272.895 692.180 273.855 ;
        RECT 697.120 272.955 697.710 273.835 ;
        RECT 698.370 272.955 700.700 273.835 ;
        RECT 701.580 272.955 702.170 273.915 ;
        RECT 704.360 272.915 704.950 273.795 ;
        RECT 705.610 272.915 707.940 273.795 ;
        RECT 708.820 272.915 709.410 273.875 ;
        RECT 714.690 273.055 715.280 273.935 ;
        RECT 715.940 273.055 718.270 273.935 ;
        RECT 719.150 273.055 719.740 274.015 ;
        RECT 721.930 273.015 722.520 273.895 ;
        RECT 723.180 273.015 725.510 273.895 ;
        RECT 726.390 273.015 726.980 273.975 ;
        RECT 731.860 273.085 732.450 273.965 ;
        RECT 733.110 273.085 735.440 273.965 ;
        RECT 736.320 273.085 736.910 274.045 ;
        RECT 739.100 273.045 739.690 273.925 ;
        RECT 740.350 273.045 742.680 273.925 ;
        RECT 743.560 273.045 744.150 274.005 ;
        RECT 749.670 273.145 750.260 274.025 ;
        RECT 750.920 273.145 753.250 274.025 ;
        RECT 754.130 273.145 754.720 274.105 ;
        RECT 756.910 273.105 757.500 273.985 ;
        RECT 758.160 273.105 760.490 273.985 ;
        RECT 761.370 273.105 761.960 274.065 ;
        RECT 595.850 271.255 596.440 272.215 ;
        RECT 635.070 271.705 635.660 272.665 ;
        RECT 639.260 271.795 639.850 272.755 ;
        RECT 643.360 271.775 643.950 272.735 ;
        RECT 679.800 272.485 685.080 272.655 ;
        RECT 687.040 272.445 692.320 272.615 ;
        RECT 697.030 272.505 702.310 272.675 ;
        RECT 704.270 272.465 709.550 272.635 ;
        RECT 714.600 272.605 719.880 272.775 ;
        RECT 721.840 272.565 727.120 272.735 ;
        RECT 731.770 272.635 737.050 272.805 ;
        RECT 739.010 272.595 744.290 272.765 ;
        RECT 749.580 272.695 754.860 272.865 ;
        RECT 756.820 272.655 762.100 272.825 ;
        RECT 781.520 271.775 782.470 272.405 ;
        RECT 783.160 271.775 783.750 272.655 ;
        RECT 788.120 271.775 789.070 272.355 ;
        RECT 792.090 271.775 793.040 272.325 ;
        RECT 794.695 271.775 795.645 272.905 ;
        RECT 800.410 271.765 801.360 272.395 ;
        RECT 802.050 271.765 802.640 272.645 ;
        RECT 807.010 271.765 807.960 272.345 ;
        RECT 810.980 271.765 811.930 272.315 ;
        RECT 813.585 271.765 814.535 272.895 ;
        RECT 819.260 271.735 820.210 272.365 ;
        RECT 820.900 271.735 821.490 272.615 ;
        RECT 825.860 271.735 826.810 272.315 ;
        RECT 829.830 271.735 830.780 272.285 ;
        RECT 832.435 271.735 833.385 272.865 ;
        RECT 840.855 271.775 841.660 272.735 ;
        RECT 857.565 271.725 858.555 272.685 ;
        RECT 595.090 270.805 596.530 270.975 ;
        RECT 143.460 270.470 147.910 270.500 ;
        RECT 121.400 269.210 125.840 270.090 ;
        RECT 143.460 269.890 149.260 270.470 ;
        RECT 596.330 270.020 596.900 270.320 ;
        RECT 143.460 269.790 147.910 269.890 ;
        RECT 150.860 268.280 151.140 268.300 ;
        RECT 150.220 268.270 151.150 268.280 ;
        RECT 118.740 268.240 151.150 268.270 ;
        RECT 118.200 268.070 151.150 268.240 ;
        RECT 118.740 268.000 151.150 268.070 ;
        RECT 118.740 267.960 150.310 268.000 ;
        RECT 150.860 265.010 151.140 268.000 ;
        RECT 605.050 266.760 605.940 271.230 ;
        RECT 614.740 268.480 614.910 268.900 ;
        RECT 616.320 268.480 616.490 268.900 ;
        RECT 614.740 267.010 614.910 267.430 ;
        RECT 616.320 267.010 616.490 267.430 ;
        RECT 625.230 266.860 626.150 271.360 ;
        RECT 634.980 271.255 636.420 271.425 ;
        RECT 639.170 271.345 640.610 271.515 ;
        RECT 643.270 271.325 644.710 271.495 ;
        RECT 780.960 271.325 796.320 271.495 ;
        RECT 799.850 271.315 815.210 271.485 ;
        RECT 818.700 271.285 834.060 271.455 ;
        RECT 838.420 271.325 842.260 271.495 ;
        RECT 855.930 271.275 859.290 271.445 ;
        RECT 846.305 269.515 847.295 270.475 ;
        RECT 850.170 269.525 850.760 270.485 ;
        RECT 844.670 269.065 848.030 269.235 ;
        RECT 850.080 269.075 851.520 269.245 ;
        RECT 640.090 267.590 640.260 268.010 ;
        RECT 644.140 267.640 644.310 268.060 ;
        RECT 681.555 267.255 682.545 268.215 ;
        RECT 687.215 267.265 688.205 268.225 ;
        RECT 691.020 267.285 691.930 267.915 ;
        RECT 692.970 267.285 693.560 268.245 ;
        RECT 698.785 267.275 699.775 268.235 ;
        RECT 704.445 267.285 705.435 268.245 ;
        RECT 708.250 267.305 709.160 267.935 ;
        RECT 710.200 267.305 710.790 268.265 ;
        RECT 716.355 267.375 717.345 268.335 ;
        RECT 722.015 267.385 723.005 268.345 ;
        RECT 725.820 267.405 726.730 268.035 ;
        RECT 727.770 267.405 728.360 268.365 ;
        RECT 733.525 267.405 734.515 268.365 ;
        RECT 739.185 267.415 740.175 268.375 ;
        RECT 742.990 267.435 743.900 268.065 ;
        RECT 744.940 267.435 745.530 268.395 ;
        RECT 749.825 268.275 750.235 268.945 ;
        RECT 751.335 267.465 752.325 268.425 ;
        RECT 756.995 267.475 757.985 268.435 ;
        RECT 760.800 267.495 761.710 268.125 ;
        RECT 762.750 267.495 763.340 268.455 ;
        RECT 861.340 268.335 862.250 268.965 ;
        RECT 863.290 268.335 863.880 269.295 ;
        RECT 861.250 267.885 864.610 268.055 ;
        RECT 679.920 266.805 683.280 266.975 ;
        RECT 685.580 266.815 688.940 266.985 ;
        RECT 690.930 266.835 694.290 267.005 ;
        RECT 697.150 266.825 700.510 266.995 ;
        RECT 702.810 266.835 706.170 267.005 ;
        RECT 708.160 266.855 711.520 267.025 ;
        RECT 714.720 266.925 718.080 267.095 ;
        RECT 720.380 266.935 723.740 267.105 ;
        RECT 725.730 266.955 729.090 267.125 ;
        RECT 731.890 266.955 735.250 267.125 ;
        RECT 737.550 266.965 740.910 267.135 ;
        RECT 742.900 266.985 746.260 267.155 ;
        RECT 749.700 267.015 753.060 267.185 ;
        RECT 755.360 267.025 758.720 267.195 ;
        RECT 760.710 267.045 764.070 267.215 ;
        RECT 840.065 266.215 841.055 267.175 ;
        RECT 838.430 265.765 841.790 265.935 ;
        RECT 151.800 265.010 152.550 265.530 ;
        RECT 117.520 264.990 118.910 265.000 ;
        RECT 150.170 264.990 152.550 265.010 ;
        RECT 117.520 264.700 152.550 264.990 ;
        RECT 117.520 264.680 150.320 264.700 ;
        RECT 117.520 264.660 118.910 264.680 ;
        RECT 150.860 261.740 151.140 264.700 ;
        RECT 151.800 264.460 152.550 264.700 ;
        RECT 781.530 264.215 782.480 264.845 ;
        RECT 783.170 264.215 783.760 265.095 ;
        RECT 788.130 264.215 789.080 264.795 ;
        RECT 792.100 264.215 793.050 264.765 ;
        RECT 794.705 264.215 795.655 265.345 ;
        RECT 800.060 264.275 801.010 264.905 ;
        RECT 801.700 264.275 802.290 265.155 ;
        RECT 806.660 264.275 807.610 264.855 ;
        RECT 810.630 264.275 811.580 264.825 ;
        RECT 813.235 264.275 814.185 265.405 ;
        RECT 857.645 265.055 858.635 266.015 ;
        RECT 856.010 264.605 859.370 264.775 ;
        RECT 780.970 263.765 796.330 263.935 ;
        RECT 799.500 263.825 814.860 263.995 ;
        RECT 147.420 261.720 147.790 261.730 ;
        RECT 150.080 261.720 151.140 261.740 ;
        RECT 118.640 261.660 151.140 261.720 ;
        RECT 118.200 261.490 151.140 261.660 ;
        RECT 118.640 261.440 151.140 261.490 ;
        RECT 118.640 261.430 151.120 261.440 ;
        RECT 118.640 261.410 150.210 261.430 ;
        RECT 147.420 260.790 147.790 261.410 ;
        RECT 121.480 259.500 125.920 260.380 ;
        RECT 143.540 260.080 147.990 260.790 ;
        RECT -91.530 236.810 -78.200 236.980 ;
        RECT -98.520 232.045 -98.350 235.125 ;
        RECT -97.850 232.930 -97.680 234.550 ;
        RECT -95.270 232.930 -95.100 234.550 ;
        RECT -92.690 232.930 -92.520 234.550 ;
        RECT -90.110 232.930 -89.940 234.550 ;
        RECT -87.530 232.930 -87.360 234.550 ;
        RECT -84.950 232.930 -84.780 234.550 ;
        RECT -82.370 232.930 -82.200 234.550 ;
        RECT -79.790 232.930 -79.620 234.550 ;
        RECT -77.210 232.930 -77.040 234.550 ;
        RECT -74.630 232.930 -74.460 234.550 ;
        RECT -72.050 232.930 -71.880 234.550 ;
        RECT -71.380 232.045 -71.210 235.125 ;
        RECT -97.075 231.050 -72.575 231.085 ;
        RECT -97.410 230.880 -72.320 231.050 ;
        RECT -97.075 230.835 -72.575 230.880 ;
        RECT -82.335 230.470 -82.165 230.835 ;
        RECT -91.610 227.850 -78.120 230.470 ;
        RECT 122.490 225.350 124.280 259.500 ;
        RECT 699.530 258.860 699.860 258.870 ;
        RECT 717.320 258.860 717.650 258.910 ;
        RECT 734.580 258.860 734.910 258.940 ;
        RECT 752.050 258.870 752.380 258.930 ;
        RECT 681.415 258.475 682.605 258.850 ;
        RECT 698.695 258.485 699.885 258.860 ;
        RECT 716.465 258.485 717.655 258.860 ;
        RECT 733.705 258.660 734.910 258.860 ;
        RECT 733.705 258.485 734.895 258.660 ;
        RECT 751.185 258.650 752.380 258.870 ;
        RECT 751.185 258.495 752.375 258.650 ;
        RECT 679.460 257.065 680.050 257.945 ;
        RECT 680.710 257.065 683.040 257.945 ;
        RECT 683.920 257.065 684.510 258.025 ;
        RECT 696.740 257.075 697.330 257.955 ;
        RECT 697.990 257.075 700.320 257.955 ;
        RECT 701.200 257.075 701.790 258.035 ;
        RECT 714.510 257.075 715.100 257.955 ;
        RECT 715.760 257.075 718.090 257.955 ;
        RECT 718.970 257.075 719.560 258.035 ;
        RECT 731.750 257.075 732.340 257.955 ;
        RECT 733.000 257.075 735.330 257.955 ;
        RECT 736.210 257.075 736.800 258.035 ;
        RECT 749.230 257.085 749.820 257.965 ;
        RECT 750.480 257.085 752.810 257.965 ;
        RECT 753.690 257.085 754.280 258.045 ;
        RECT 679.370 256.615 684.650 256.785 ;
        RECT 696.650 256.625 701.930 256.795 ;
        RECT 714.420 256.625 719.700 256.795 ;
        RECT 731.660 256.625 736.940 256.795 ;
        RECT 749.140 256.635 754.420 256.805 ;
        RECT 857.515 255.745 858.505 256.705 ;
        RECT 855.880 255.295 859.240 255.465 ;
        RECT 595.700 253.525 596.290 254.485 ;
        RECT 634.920 253.975 635.510 254.935 ;
        RECT 639.110 254.065 639.700 255.025 ;
        RECT 643.210 254.045 643.800 255.005 ;
        RECT 594.940 253.075 596.380 253.245 ;
        RECT 596.180 252.290 596.750 252.590 ;
        RECT 604.900 249.030 605.790 253.500 ;
        RECT 614.590 250.750 614.760 251.170 ;
        RECT 616.170 250.750 616.340 251.170 ;
        RECT 614.590 249.280 614.760 249.700 ;
        RECT 616.170 249.280 616.340 249.700 ;
        RECT 625.080 249.130 626.000 253.630 ;
        RECT 634.830 253.525 636.270 253.695 ;
        RECT 639.020 253.615 640.460 253.785 ;
        RECT 643.120 253.595 644.560 253.765 ;
        RECT 645.650 253.630 646.300 254.940 ;
        RECT 681.825 252.815 683.015 253.190 ;
        RECT 751.605 253.025 752.795 253.400 ;
        RECT 757.360 252.985 758.310 253.265 ;
        RECT 861.280 253.255 862.190 253.885 ;
        RECT 863.230 253.255 863.820 254.215 ;
        RECT 758.140 252.805 758.310 252.985 ;
        RECT 760.215 252.805 760.515 253.045 ;
        RECT 861.190 252.805 864.550 252.975 ;
        RECT 758.140 252.715 760.515 252.805 ;
        RECT 758.140 252.635 760.385 252.715 ;
        RECT 679.870 251.405 680.460 252.285 ;
        RECT 681.120 251.405 683.450 252.285 ;
        RECT 684.330 251.405 684.920 252.365 ;
        RECT 687.110 251.365 687.700 252.245 ;
        RECT 688.360 251.365 690.690 252.245 ;
        RECT 691.570 251.365 692.160 252.325 ;
        RECT 697.100 251.425 697.690 252.305 ;
        RECT 698.350 251.425 700.680 252.305 ;
        RECT 701.560 251.425 702.150 252.385 ;
        RECT 704.340 251.385 704.930 252.265 ;
        RECT 705.590 251.385 707.920 252.265 ;
        RECT 708.800 251.385 709.390 252.345 ;
        RECT 714.670 251.525 715.260 252.405 ;
        RECT 715.920 251.525 718.250 252.405 ;
        RECT 719.130 251.525 719.720 252.485 ;
        RECT 721.910 251.485 722.500 252.365 ;
        RECT 723.160 251.485 725.490 252.365 ;
        RECT 726.370 251.485 726.960 252.445 ;
        RECT 731.840 251.555 732.430 252.435 ;
        RECT 733.090 251.555 735.420 252.435 ;
        RECT 736.300 251.555 736.890 252.515 ;
        RECT 739.080 251.515 739.670 252.395 ;
        RECT 740.330 251.515 742.660 252.395 ;
        RECT 743.540 251.515 744.130 252.475 ;
        RECT 749.650 251.615 750.240 252.495 ;
        RECT 750.900 251.615 753.230 252.495 ;
        RECT 754.110 251.615 754.700 252.575 ;
        RECT 756.890 251.575 757.480 252.455 ;
        RECT 758.140 251.575 760.470 252.455 ;
        RECT 761.350 251.575 761.940 252.535 ;
        RECT 679.780 250.955 685.060 251.125 ;
        RECT 687.020 250.915 692.300 251.085 ;
        RECT 697.010 250.975 702.290 251.145 ;
        RECT 704.250 250.935 709.530 251.105 ;
        RECT 714.580 251.075 719.860 251.245 ;
        RECT 721.820 251.035 727.100 251.205 ;
        RECT 731.750 251.105 737.030 251.275 ;
        RECT 738.990 251.065 744.270 251.235 ;
        RECT 749.560 251.165 754.840 251.335 ;
        RECT 756.800 251.125 762.080 251.295 ;
        RECT 639.940 249.860 640.110 250.280 ;
        RECT 643.990 249.910 644.160 250.330 ;
        RECT 857.575 249.975 858.565 250.935 ;
        RECT 855.940 249.525 859.300 249.695 ;
        RECT 601.550 248.380 602.610 248.820 ;
        RECT 591.430 245.220 591.780 247.380 ;
        RECT 680.025 246.535 680.435 247.205 ;
        RECT 681.535 245.725 682.525 246.685 ;
        RECT 687.195 245.735 688.185 246.695 ;
        RECT 691.000 245.755 691.910 246.385 ;
        RECT 692.950 245.755 693.540 246.715 ;
        RECT 698.765 245.745 699.755 246.705 ;
        RECT 704.425 245.755 705.415 246.715 ;
        RECT 708.230 245.775 709.140 246.405 ;
        RECT 710.180 245.775 710.770 246.735 ;
        RECT 716.335 245.845 717.325 246.805 ;
        RECT 721.995 245.855 722.985 246.815 ;
        RECT 725.800 245.875 726.710 246.505 ;
        RECT 727.750 245.875 728.340 246.835 ;
        RECT 733.505 245.875 734.495 246.835 ;
        RECT 739.165 245.885 740.155 246.845 ;
        RECT 742.970 245.905 743.880 246.535 ;
        RECT 744.920 245.905 745.510 246.865 ;
        RECT 749.805 246.745 750.215 247.415 ;
        RECT 756.405 247.110 756.795 247.305 ;
        RECT 751.315 245.935 752.305 246.895 ;
        RECT 756.405 246.530 756.800 247.110 ;
        RECT 756.405 246.390 756.795 246.530 ;
        RECT 756.975 245.945 757.965 246.905 ;
        RECT 760.780 245.965 761.690 246.595 ;
        RECT 762.730 245.965 763.320 246.925 ;
        RECT 679.900 245.275 683.260 245.445 ;
        RECT 685.560 245.285 688.920 245.455 ;
        RECT 690.910 245.305 694.270 245.475 ;
        RECT 697.130 245.295 700.490 245.465 ;
        RECT 702.790 245.305 706.150 245.475 ;
        RECT 708.140 245.325 711.500 245.495 ;
        RECT 714.700 245.395 718.060 245.565 ;
        RECT 720.360 245.405 723.720 245.575 ;
        RECT 725.710 245.425 729.070 245.595 ;
        RECT 731.870 245.425 735.230 245.595 ;
        RECT 737.530 245.435 740.890 245.605 ;
        RECT 742.880 245.455 746.240 245.625 ;
        RECT 749.680 245.485 753.040 245.655 ;
        RECT 755.340 245.495 758.700 245.665 ;
        RECT 760.690 245.515 764.050 245.685 ;
        RECT -90.840 224.710 -77.510 224.880 ;
        RECT -97.830 219.945 -97.660 223.025 ;
        RECT -97.160 220.830 -96.990 222.450 ;
        RECT -94.580 220.830 -94.410 222.450 ;
        RECT -92.000 220.830 -91.830 222.450 ;
        RECT -89.420 220.830 -89.250 222.450 ;
        RECT -86.840 220.830 -86.670 222.450 ;
        RECT -84.260 220.830 -84.090 222.450 ;
        RECT -81.680 220.830 -81.510 222.450 ;
        RECT -79.100 220.830 -78.930 222.450 ;
        RECT -76.520 220.830 -76.350 222.450 ;
        RECT -73.940 220.830 -73.770 222.450 ;
        RECT -71.360 220.830 -71.190 222.450 ;
        RECT -70.690 219.945 -70.520 223.025 ;
        RECT 120.120 222.910 127.210 225.350 ;
        RECT 193.570 221.540 213.970 225.890 ;
        RECT -96.385 218.950 -71.885 218.985 ;
        RECT -96.720 218.780 -71.630 218.950 ;
        RECT -96.385 218.735 -71.885 218.780 ;
        RECT -81.645 218.350 -81.475 218.735 ;
        RECT -90.980 215.730 -77.490 218.350 ;
        RECT 9.550 216.650 10.230 218.130 ;
        RECT 55.080 217.830 56.450 218.870 ;
        RECT 247.270 218.070 250.350 220.020 ;
        RECT 341.380 218.910 345.300 219.920 ;
        RECT 36.200 216.810 36.880 216.950 ;
        RECT 20.240 216.650 20.580 216.730 ;
        RECT 30.860 216.690 43.240 216.810 ;
        RECT 52.810 216.690 53.150 216.770 ;
        RECT 55.390 216.690 55.960 217.830 ;
        RECT 63.430 216.760 63.770 216.850 ;
        RECT 74.820 216.760 75.160 216.780 ;
        RECT 63.120 216.730 77.130 216.760 ;
        RECT 85.340 216.730 85.680 216.810 ;
        RECT 95.960 216.730 96.300 216.890 ;
        RECT 204.880 216.760 205.220 216.810 ;
        RECT 215.400 216.760 215.740 216.840 ;
        RECT 226.020 216.760 226.360 216.920 ;
        RECT 237.820 216.870 238.160 216.920 ;
        RECT 248.210 216.870 249.190 218.070 ;
        RECT 258.960 216.870 259.300 217.030 ;
        RECT 270.390 216.940 270.730 216.990 ;
        RECT 280.910 216.940 281.250 217.020 ;
        RECT 291.530 216.940 291.870 217.100 ;
        RECT 270.390 216.900 291.870 216.940 ;
        RECT 296.740 216.900 297.230 217.280 ;
        RECT 318.960 217.220 321.190 218.260 ;
        RECT 270.390 216.890 297.230 216.900 ;
        RECT 237.820 216.820 259.300 216.870 ;
        RECT 63.120 216.700 96.300 216.730 ;
        RECT 101.270 216.700 101.690 216.750 ;
        RECT 204.880 216.720 226.360 216.760 ;
        RECT 204.340 216.710 226.360 216.720 ;
        RECT 63.120 216.690 101.690 216.700 ;
        RECT 30.860 216.650 101.690 216.690 ;
        RECT 9.550 216.600 101.690 216.650 ;
        RECT 9.030 216.280 101.690 216.600 ;
        RECT 9.030 216.230 95.580 216.280 ;
        RECT 9.030 216.200 77.130 216.230 ;
        RECT 9.030 216.150 30.480 216.200 ;
        RECT 30.820 216.190 77.130 216.200 ;
        RECT 6.520 199.990 7.270 208.220 ;
        RECT 9.550 187.570 10.230 216.150 ;
        RECT 15.080 214.790 15.250 215.340 ;
        RECT 20.240 215.080 20.580 216.150 ;
        RECT 30.820 215.580 43.240 216.190 ;
        RECT 20.240 214.820 20.610 215.080 ;
        RECT 25.660 214.820 25.830 215.340 ;
        RECT 15.060 192.980 15.290 214.790 ;
        RECT 20.320 193.090 20.550 214.820 ;
        RECT 15.080 192.420 15.250 192.980 ;
        RECT 14.980 191.370 15.390 192.420 ;
        RECT 20.370 191.840 20.540 193.090 ;
        RECT 25.660 193.010 25.890 214.820 ;
        RECT 30.820 214.800 31.240 215.580 ;
        RECT 30.920 193.230 31.150 214.800 ;
        RECT 25.660 192.280 25.830 193.010 ;
        RECT 25.610 191.370 26.020 192.280 ;
        RECT 30.950 191.840 31.120 193.230 ;
        RECT 36.200 192.390 36.880 215.580 ;
        RECT 36.120 191.370 36.880 192.390 ;
        RECT 14.980 190.920 37.230 191.370 ;
        RECT 15.040 190.890 37.230 190.920 ;
        RECT 25.610 190.780 26.020 190.890 ;
        RECT 20.240 187.570 20.580 187.650 ;
        RECT 30.860 187.570 31.200 187.730 ;
        RECT 9.550 187.520 31.200 187.570 ;
        RECT 9.030 187.300 31.200 187.520 ;
        RECT 9.030 187.120 31.240 187.300 ;
        RECT 9.030 187.070 30.480 187.120 ;
        RECT 6.520 170.910 7.270 179.140 ;
        RECT 9.550 158.400 10.230 187.070 ;
        RECT 15.080 185.710 15.250 186.260 ;
        RECT 20.240 186.000 20.580 187.070 ;
        RECT 20.240 185.740 20.610 186.000 ;
        RECT 25.660 185.740 25.830 186.260 ;
        RECT 15.060 163.900 15.290 185.710 ;
        RECT 20.320 164.010 20.550 185.740 ;
        RECT 15.080 163.340 15.250 163.900 ;
        RECT 14.980 162.290 15.390 163.340 ;
        RECT 20.370 162.760 20.540 164.010 ;
        RECT 25.660 163.930 25.890 185.740 ;
        RECT 30.820 185.720 31.240 187.120 ;
        RECT 30.920 164.150 31.150 185.720 ;
        RECT 25.660 163.200 25.830 163.930 ;
        RECT 25.610 162.290 26.020 163.200 ;
        RECT 30.950 162.760 31.120 164.150 ;
        RECT 36.200 163.310 36.880 190.890 ;
        RECT 36.120 162.290 36.880 163.310 ;
        RECT 14.980 161.840 37.230 162.290 ;
        RECT 15.040 161.810 37.230 161.840 ;
        RECT 25.610 161.700 26.020 161.810 ;
        RECT 20.240 158.400 20.580 158.480 ;
        RECT 30.860 158.400 31.200 158.560 ;
        RECT 9.550 158.350 31.200 158.400 ;
        RECT 9.030 158.130 31.200 158.350 ;
        RECT 9.030 157.950 31.240 158.130 ;
        RECT 9.030 157.900 30.480 157.950 ;
        RECT 6.520 141.740 7.270 149.970 ;
        RECT -91.240 136.960 -77.910 137.130 ;
        RECT -98.230 132.195 -98.060 135.275 ;
        RECT -97.560 133.080 -97.390 134.700 ;
        RECT -94.980 133.080 -94.810 134.700 ;
        RECT -92.400 133.080 -92.230 134.700 ;
        RECT -89.820 133.080 -89.650 134.700 ;
        RECT -87.240 133.080 -87.070 134.700 ;
        RECT -84.660 133.080 -84.490 134.700 ;
        RECT -82.080 133.080 -81.910 134.700 ;
        RECT -79.500 133.080 -79.330 134.700 ;
        RECT -76.920 133.080 -76.750 134.700 ;
        RECT -74.340 133.080 -74.170 134.700 ;
        RECT -71.760 133.080 -71.590 134.700 ;
        RECT -71.090 132.195 -70.920 135.275 ;
        RECT -96.785 131.200 -72.285 131.235 ;
        RECT -97.120 131.030 -72.030 131.200 ;
        RECT -96.785 130.985 -72.285 131.030 ;
        RECT -82.045 130.510 -81.875 130.985 ;
        RECT -91.440 130.340 -77.910 130.510 ;
        RECT -91.440 127.890 -77.950 130.340 ;
        RECT 9.550 129.220 10.230 157.900 ;
        RECT 15.080 156.540 15.250 157.090 ;
        RECT 20.240 156.830 20.580 157.900 ;
        RECT 20.240 156.570 20.610 156.830 ;
        RECT 25.660 156.570 25.830 157.090 ;
        RECT 15.060 134.730 15.290 156.540 ;
        RECT 20.320 134.840 20.550 156.570 ;
        RECT 15.080 134.170 15.250 134.730 ;
        RECT 14.980 133.120 15.390 134.170 ;
        RECT 20.370 133.590 20.540 134.840 ;
        RECT 25.660 134.760 25.890 156.570 ;
        RECT 30.820 156.550 31.240 157.950 ;
        RECT 30.920 134.980 31.150 156.550 ;
        RECT 25.660 134.030 25.830 134.760 ;
        RECT 25.610 133.120 26.020 134.030 ;
        RECT 30.950 133.590 31.120 134.980 ;
        RECT 36.200 134.140 36.880 161.810 ;
        RECT 36.120 133.120 36.880 134.140 ;
        RECT 14.980 132.670 37.230 133.120 ;
        RECT 15.040 132.640 37.230 132.670 ;
        RECT 25.610 132.530 26.020 132.640 ;
        RECT 20.240 129.220 20.580 129.300 ;
        RECT 30.860 129.220 31.200 129.380 ;
        RECT 9.550 129.170 31.200 129.220 ;
        RECT 9.030 128.950 31.200 129.170 ;
        RECT 9.030 128.770 31.240 128.950 ;
        RECT 9.030 128.720 30.480 128.770 ;
        RECT 6.520 112.560 7.270 120.790 ;
        RECT 9.550 99.900 10.230 128.720 ;
        RECT 15.080 127.360 15.250 127.910 ;
        RECT 20.240 127.650 20.580 128.720 ;
        RECT 20.240 127.390 20.610 127.650 ;
        RECT 25.660 127.390 25.830 127.910 ;
        RECT 15.060 105.550 15.290 127.360 ;
        RECT 20.320 105.660 20.550 127.390 ;
        RECT 15.080 104.990 15.250 105.550 ;
        RECT 14.980 103.940 15.390 104.990 ;
        RECT 20.370 104.410 20.540 105.660 ;
        RECT 25.660 105.580 25.890 127.390 ;
        RECT 30.820 127.370 31.240 128.770 ;
        RECT 30.920 105.800 31.150 127.370 ;
        RECT 25.660 104.850 25.830 105.580 ;
        RECT 25.610 103.940 26.020 104.850 ;
        RECT 30.950 104.410 31.120 105.800 ;
        RECT 36.200 104.960 36.880 132.640 ;
        RECT 36.120 103.940 36.880 104.960 ;
        RECT 14.980 103.490 37.230 103.940 ;
        RECT 15.040 103.460 37.230 103.490 ;
        RECT 25.610 103.350 26.020 103.460 ;
        RECT 20.240 99.900 20.580 99.980 ;
        RECT 30.860 99.900 31.200 100.060 ;
        RECT 9.550 99.850 31.200 99.900 ;
        RECT 9.030 99.630 31.200 99.850 ;
        RECT 9.030 99.450 31.240 99.630 ;
        RECT 9.030 99.400 30.480 99.450 ;
        RECT 6.520 83.240 7.270 91.470 ;
        RECT 9.550 70.620 10.230 99.400 ;
        RECT 15.080 98.040 15.250 98.590 ;
        RECT 20.240 98.330 20.580 99.400 ;
        RECT 20.240 98.070 20.610 98.330 ;
        RECT 25.660 98.070 25.830 98.590 ;
        RECT 15.060 76.230 15.290 98.040 ;
        RECT 20.320 76.340 20.550 98.070 ;
        RECT 15.080 75.670 15.250 76.230 ;
        RECT 14.980 74.620 15.390 75.670 ;
        RECT 20.370 75.090 20.540 76.340 ;
        RECT 25.660 76.260 25.890 98.070 ;
        RECT 30.820 98.050 31.240 99.450 ;
        RECT 30.920 76.480 31.150 98.050 ;
        RECT 25.660 75.530 25.830 76.260 ;
        RECT 25.610 74.620 26.020 75.530 ;
        RECT 30.950 75.090 31.120 76.480 ;
        RECT 36.200 75.640 36.880 103.460 ;
        RECT 36.120 74.620 36.880 75.640 ;
        RECT 14.980 74.170 37.230 74.620 ;
        RECT 15.040 74.140 37.230 74.170 ;
        RECT 25.610 74.030 26.020 74.140 ;
        RECT 20.290 70.620 20.630 70.700 ;
        RECT 30.910 70.620 31.250 70.780 ;
        RECT 9.550 70.570 31.250 70.620 ;
        RECT 9.080 70.350 31.250 70.570 ;
        RECT 9.080 70.170 31.290 70.350 ;
        RECT 9.080 70.120 30.530 70.170 ;
        RECT 6.570 53.960 7.320 62.190 ;
        RECT 9.550 41.080 10.230 70.120 ;
        RECT 15.130 68.760 15.300 69.310 ;
        RECT 20.290 69.050 20.630 70.120 ;
        RECT 20.290 68.790 20.660 69.050 ;
        RECT 25.710 68.790 25.880 69.310 ;
        RECT 15.110 46.950 15.340 68.760 ;
        RECT 20.370 47.060 20.600 68.790 ;
        RECT 15.130 46.390 15.300 46.950 ;
        RECT 15.030 45.340 15.440 46.390 ;
        RECT 20.420 45.810 20.590 47.060 ;
        RECT 25.710 46.980 25.940 68.790 ;
        RECT 30.870 68.770 31.290 70.170 ;
        RECT 30.970 47.200 31.200 68.770 ;
        RECT 25.710 46.250 25.880 46.980 ;
        RECT 25.660 45.340 26.070 46.250 ;
        RECT 31.000 45.810 31.170 47.200 ;
        RECT 36.200 46.360 36.880 74.140 ;
        RECT 36.170 45.340 36.880 46.360 ;
        RECT 15.030 44.890 37.280 45.340 ;
        RECT 15.090 44.860 37.280 44.890 ;
        RECT 25.660 44.750 26.070 44.860 ;
        RECT 20.380 41.080 20.720 41.160 ;
        RECT 31.000 41.080 31.340 41.240 ;
        RECT 9.550 41.030 31.340 41.080 ;
        RECT 9.170 40.810 31.340 41.030 ;
        RECT 9.170 40.630 31.380 40.810 ;
        RECT 9.170 40.580 30.620 40.630 ;
        RECT 9.550 40.040 10.230 40.580 ;
        RECT 9.860 39.180 10.200 40.040 ;
        RECT 15.220 39.220 15.390 39.770 ;
        RECT 20.380 39.510 20.720 40.580 ;
        RECT 20.380 39.250 20.750 39.510 ;
        RECT 25.800 39.250 25.970 39.770 ;
        RECT 9.860 38.150 10.100 39.180 ;
        RECT 9.860 34.300 10.090 38.150 ;
        RECT 9.860 32.680 10.100 34.300 ;
        RECT 6.660 24.420 7.410 32.650 ;
        RECT 9.860 28.830 10.090 32.680 ;
        RECT 9.860 27.210 10.100 28.830 ;
        RECT 9.860 23.360 10.090 27.210 ;
        RECT 9.860 21.740 10.100 23.360 ;
        RECT 9.860 17.890 10.090 21.740 ;
        RECT -90.810 17.630 -77.480 17.800 ;
        RECT 9.860 17.520 10.100 17.890 ;
        RECT 9.930 16.270 10.100 17.520 ;
        RECT 15.200 17.410 15.430 39.220 ;
        RECT 20.460 17.520 20.690 39.250 ;
        RECT 15.220 16.850 15.390 17.410 ;
        RECT -97.800 12.865 -97.630 15.945 ;
        RECT -97.130 13.750 -96.960 15.370 ;
        RECT -94.550 13.750 -94.380 15.370 ;
        RECT -91.970 13.750 -91.800 15.370 ;
        RECT -89.390 13.750 -89.220 15.370 ;
        RECT -86.810 13.750 -86.640 15.370 ;
        RECT -84.230 13.750 -84.060 15.370 ;
        RECT -81.650 13.750 -81.480 15.370 ;
        RECT -79.070 13.750 -78.900 15.370 ;
        RECT -76.490 13.750 -76.320 15.370 ;
        RECT -73.910 13.750 -73.740 15.370 ;
        RECT -71.330 13.750 -71.160 15.370 ;
        RECT -70.660 12.865 -70.490 15.945 ;
        RECT 15.120 15.800 15.530 16.850 ;
        RECT 20.510 16.270 20.680 17.520 ;
        RECT 25.800 17.440 26.030 39.250 ;
        RECT 30.960 39.230 31.380 40.630 ;
        RECT 31.060 17.660 31.290 39.230 ;
        RECT 36.200 38.860 36.880 44.860 ;
        RECT 25.800 16.710 25.970 17.440 ;
        RECT 25.750 15.800 26.160 16.710 ;
        RECT 31.090 16.270 31.260 17.660 ;
        RECT 36.340 17.520 36.570 38.860 ;
        RECT 37.980 24.860 41.260 210.950 ;
        RECT 42.180 187.610 42.860 215.580 ;
        RECT 47.650 214.830 47.820 215.380 ;
        RECT 52.810 215.120 53.150 216.190 ;
        RECT 62.890 216.120 77.130 216.190 ;
        RECT 52.810 214.860 53.180 215.120 ;
        RECT 58.230 214.860 58.400 215.380 ;
        RECT 47.630 193.020 47.860 214.830 ;
        RECT 52.890 193.130 53.120 214.860 ;
        RECT 47.650 192.460 47.820 193.020 ;
        RECT 47.550 191.410 47.960 192.460 ;
        RECT 52.940 191.880 53.110 193.130 ;
        RECT 58.230 193.050 58.460 214.860 ;
        RECT 63.390 214.840 63.810 216.120 ;
        RECT 68.730 215.110 69.440 216.120 ;
        RECT 68.710 215.030 69.440 215.110 ;
        RECT 68.710 214.860 69.370 215.030 ;
        RECT 63.490 193.270 63.720 214.840 ;
        RECT 58.230 192.320 58.400 193.050 ;
        RECT 58.180 191.410 58.590 192.320 ;
        RECT 63.520 191.880 63.690 193.270 ;
        RECT 68.770 193.130 69.370 214.860 ;
        RECT 74.700 214.830 75.160 216.120 ;
        RECT 80.180 214.870 80.350 215.420 ;
        RECT 85.340 215.160 85.680 216.230 ;
        RECT 95.910 216.030 101.690 216.280 ;
        RECT 204.190 216.690 226.360 216.710 ;
        RECT 237.130 216.800 259.300 216.820 ;
        RECT 269.700 216.800 297.230 216.890 ;
        RECT 237.130 216.690 297.230 216.800 ;
        RECT 204.190 216.490 297.230 216.690 ;
        RECT 204.190 216.440 291.150 216.490 ;
        RECT 204.190 216.420 272.480 216.440 ;
        RECT 204.190 216.370 258.580 216.420 ;
        RECT 204.190 216.310 239.500 216.370 ;
        RECT 204.190 216.260 225.640 216.310 ;
        RECT 85.340 214.900 85.710 215.160 ;
        RECT 90.760 214.900 90.930 215.420 ;
        RECT 68.810 192.430 69.370 193.130 ;
        RECT 68.690 191.410 69.370 192.430 ;
        RECT 47.550 190.960 69.800 191.410 ;
        RECT 47.610 190.930 69.800 190.960 ;
        RECT 58.180 190.820 58.590 190.930 ;
        RECT 52.810 187.610 53.150 187.690 ;
        RECT 63.430 187.610 63.770 187.770 ;
        RECT 42.180 187.560 63.770 187.610 ;
        RECT 41.600 187.340 63.770 187.560 ;
        RECT 41.600 187.160 63.810 187.340 ;
        RECT 41.600 187.110 63.050 187.160 ;
        RECT 42.180 158.440 42.860 187.110 ;
        RECT 47.650 185.750 47.820 186.300 ;
        RECT 52.810 186.040 53.150 187.110 ;
        RECT 52.810 185.780 53.180 186.040 ;
        RECT 58.230 185.780 58.400 186.300 ;
        RECT 47.630 163.940 47.860 185.750 ;
        RECT 52.890 164.050 53.120 185.780 ;
        RECT 47.650 163.380 47.820 163.940 ;
        RECT 47.550 162.330 47.960 163.380 ;
        RECT 52.940 162.800 53.110 164.050 ;
        RECT 58.230 163.970 58.460 185.780 ;
        RECT 63.390 185.760 63.810 187.160 ;
        RECT 68.840 186.300 69.370 190.930 ;
        RECT 68.810 185.860 69.370 186.300 ;
        RECT 63.490 164.190 63.720 185.760 ;
        RECT 58.230 163.240 58.400 163.970 ;
        RECT 58.180 162.330 58.590 163.240 ;
        RECT 63.520 162.800 63.690 164.190 ;
        RECT 68.770 164.050 69.370 185.860 ;
        RECT 68.810 163.350 69.370 164.050 ;
        RECT 68.690 162.330 69.370 163.350 ;
        RECT 47.550 161.880 69.800 162.330 ;
        RECT 47.610 161.850 69.800 161.880 ;
        RECT 58.180 161.740 58.590 161.850 ;
        RECT 52.810 158.440 53.150 158.520 ;
        RECT 63.430 158.440 63.770 158.600 ;
        RECT 42.180 158.390 63.770 158.440 ;
        RECT 41.600 158.170 63.770 158.390 ;
        RECT 41.600 157.990 63.810 158.170 ;
        RECT 41.600 157.940 63.050 157.990 ;
        RECT 42.180 129.260 42.860 157.940 ;
        RECT 47.650 156.580 47.820 157.130 ;
        RECT 52.810 156.870 53.150 157.940 ;
        RECT 52.810 156.610 53.180 156.870 ;
        RECT 58.230 156.610 58.400 157.130 ;
        RECT 47.630 134.770 47.860 156.580 ;
        RECT 52.890 134.880 53.120 156.610 ;
        RECT 47.650 134.210 47.820 134.770 ;
        RECT 47.550 133.160 47.960 134.210 ;
        RECT 52.940 133.630 53.110 134.880 ;
        RECT 58.230 134.800 58.460 156.610 ;
        RECT 63.390 156.590 63.810 157.990 ;
        RECT 68.840 157.130 69.370 161.850 ;
        RECT 68.810 156.690 69.370 157.130 ;
        RECT 63.490 135.020 63.720 156.590 ;
        RECT 58.230 134.070 58.400 134.800 ;
        RECT 58.180 133.160 58.590 134.070 ;
        RECT 63.520 133.630 63.690 135.020 ;
        RECT 68.770 134.880 69.370 156.690 ;
        RECT 68.810 134.180 69.370 134.880 ;
        RECT 68.690 133.160 69.370 134.180 ;
        RECT 47.550 132.710 69.800 133.160 ;
        RECT 47.610 132.680 69.800 132.710 ;
        RECT 58.180 132.570 58.590 132.680 ;
        RECT 52.810 129.260 53.150 129.340 ;
        RECT 63.430 129.260 63.770 129.420 ;
        RECT 42.180 129.210 63.770 129.260 ;
        RECT 41.600 128.990 63.770 129.210 ;
        RECT 41.600 128.810 63.810 128.990 ;
        RECT 41.600 128.760 63.050 128.810 ;
        RECT 42.180 99.940 42.860 128.760 ;
        RECT 47.650 127.400 47.820 127.950 ;
        RECT 52.810 127.690 53.150 128.760 ;
        RECT 52.810 127.430 53.180 127.690 ;
        RECT 58.230 127.430 58.400 127.950 ;
        RECT 47.630 105.590 47.860 127.400 ;
        RECT 52.890 105.700 53.120 127.430 ;
        RECT 47.650 105.030 47.820 105.590 ;
        RECT 47.550 103.980 47.960 105.030 ;
        RECT 52.940 104.450 53.110 105.700 ;
        RECT 58.230 105.620 58.460 127.430 ;
        RECT 63.390 127.410 63.810 128.810 ;
        RECT 68.840 127.950 69.370 132.680 ;
        RECT 68.810 127.510 69.370 127.950 ;
        RECT 63.490 105.840 63.720 127.410 ;
        RECT 58.230 104.890 58.400 105.620 ;
        RECT 58.180 103.980 58.590 104.890 ;
        RECT 63.520 104.450 63.690 105.840 ;
        RECT 68.770 105.700 69.370 127.510 ;
        RECT 68.810 105.000 69.370 105.700 ;
        RECT 68.690 103.980 69.370 105.000 ;
        RECT 47.550 103.530 69.800 103.980 ;
        RECT 47.610 103.500 69.800 103.530 ;
        RECT 58.180 103.390 58.590 103.500 ;
        RECT 52.810 99.940 53.150 100.020 ;
        RECT 63.430 99.940 63.770 100.100 ;
        RECT 42.180 99.890 63.770 99.940 ;
        RECT 41.600 99.670 63.770 99.890 ;
        RECT 41.600 99.490 63.810 99.670 ;
        RECT 41.600 99.440 63.050 99.490 ;
        RECT 42.180 70.660 42.860 99.440 ;
        RECT 47.650 98.080 47.820 98.630 ;
        RECT 52.810 98.370 53.150 99.440 ;
        RECT 52.810 98.110 53.180 98.370 ;
        RECT 58.230 98.110 58.400 98.630 ;
        RECT 47.630 76.270 47.860 98.080 ;
        RECT 52.890 76.380 53.120 98.110 ;
        RECT 47.650 75.710 47.820 76.270 ;
        RECT 47.550 74.660 47.960 75.710 ;
        RECT 52.940 75.130 53.110 76.380 ;
        RECT 58.230 76.300 58.460 98.110 ;
        RECT 63.390 98.090 63.810 99.490 ;
        RECT 68.840 98.630 69.370 103.500 ;
        RECT 68.810 98.190 69.370 98.630 ;
        RECT 63.490 76.520 63.720 98.090 ;
        RECT 58.230 75.570 58.400 76.300 ;
        RECT 58.180 74.660 58.590 75.570 ;
        RECT 63.520 75.130 63.690 76.520 ;
        RECT 68.770 76.380 69.370 98.190 ;
        RECT 68.810 75.680 69.370 76.380 ;
        RECT 68.690 74.660 69.370 75.680 ;
        RECT 47.550 74.210 69.800 74.660 ;
        RECT 47.610 74.180 69.800 74.210 ;
        RECT 58.180 74.070 58.590 74.180 ;
        RECT 52.860 70.660 53.200 70.740 ;
        RECT 63.480 70.660 63.820 70.820 ;
        RECT 42.180 70.610 63.820 70.660 ;
        RECT 41.650 70.390 63.820 70.610 ;
        RECT 41.650 70.210 63.860 70.390 ;
        RECT 41.650 70.160 63.100 70.210 ;
        RECT 42.180 41.120 42.860 70.160 ;
        RECT 47.700 68.800 47.870 69.350 ;
        RECT 52.860 69.090 53.200 70.160 ;
        RECT 52.860 68.830 53.230 69.090 ;
        RECT 58.280 68.830 58.450 69.350 ;
        RECT 47.680 46.990 47.910 68.800 ;
        RECT 52.940 47.100 53.170 68.830 ;
        RECT 47.700 46.430 47.870 46.990 ;
        RECT 47.600 45.380 48.010 46.430 ;
        RECT 52.990 45.850 53.160 47.100 ;
        RECT 58.280 47.020 58.510 68.830 ;
        RECT 63.440 68.810 63.860 70.210 ;
        RECT 68.840 68.910 69.370 74.180 ;
        RECT 63.540 47.240 63.770 68.810 ;
        RECT 58.280 46.290 58.450 47.020 ;
        RECT 58.230 45.380 58.640 46.290 ;
        RECT 63.570 45.850 63.740 47.240 ;
        RECT 68.820 47.100 69.370 68.910 ;
        RECT 68.840 46.400 69.370 47.100 ;
        RECT 68.740 45.380 69.370 46.400 ;
        RECT 47.600 44.930 69.850 45.380 ;
        RECT 47.660 44.900 69.850 44.930 ;
        RECT 58.230 44.790 58.640 44.900 ;
        RECT 52.950 41.120 53.290 41.200 ;
        RECT 63.570 41.120 63.910 41.280 ;
        RECT 42.180 41.070 63.910 41.120 ;
        RECT 41.740 40.850 63.910 41.070 ;
        RECT 41.740 40.670 63.950 40.850 ;
        RECT 41.740 40.620 63.190 40.670 ;
        RECT 42.180 38.440 42.860 40.620 ;
        RECT 47.790 39.260 47.960 39.810 ;
        RECT 52.950 39.550 53.290 40.620 ;
        RECT 52.950 39.290 53.320 39.550 ;
        RECT 58.370 39.290 58.540 39.810 ;
        RECT 42.430 38.190 42.670 38.440 ;
        RECT 42.430 34.340 42.660 38.190 ;
        RECT 42.430 32.720 42.670 34.340 ;
        RECT 42.430 28.870 42.660 32.720 ;
        RECT 42.430 27.250 42.670 28.870 ;
        RECT 39.230 24.460 39.980 24.860 ;
        RECT 42.430 23.400 42.660 27.250 ;
        RECT 42.430 21.780 42.670 23.400 ;
        RECT 42.430 17.930 42.660 21.780 ;
        RECT 42.430 17.560 42.670 17.930 ;
        RECT 36.380 16.820 36.550 17.520 ;
        RECT 36.260 15.800 36.670 16.820 ;
        RECT 42.500 16.310 42.670 17.560 ;
        RECT 47.770 17.450 48.000 39.260 ;
        RECT 53.030 17.560 53.260 39.290 ;
        RECT 47.790 16.890 47.960 17.450 ;
        RECT 47.690 15.840 48.100 16.890 ;
        RECT 53.080 16.310 53.250 17.560 ;
        RECT 58.370 17.480 58.600 39.290 ;
        RECT 63.530 39.270 63.950 40.670 ;
        RECT 63.630 17.700 63.860 39.270 ;
        RECT 68.840 39.200 69.370 44.900 ;
        RECT 58.370 16.750 58.540 17.480 ;
        RECT 58.320 15.840 58.730 16.750 ;
        RECT 63.660 16.310 63.830 17.700 ;
        RECT 68.910 17.560 69.140 39.200 ;
        RECT 68.950 16.860 69.120 17.560 ;
        RECT 70.230 16.890 73.430 208.450 ;
        RECT 74.700 187.700 75.140 214.830 ;
        RECT 80.160 193.060 80.390 214.870 ;
        RECT 85.420 193.170 85.650 214.900 ;
        RECT 80.180 192.500 80.350 193.060 ;
        RECT 80.080 191.450 80.490 192.500 ;
        RECT 85.470 191.920 85.640 193.170 ;
        RECT 90.760 193.090 90.990 214.900 ;
        RECT 95.920 214.880 96.340 216.030 ;
        RECT 101.210 214.930 101.690 216.030 ;
        RECT 204.340 215.810 205.650 216.260 ;
        RECT 96.020 193.310 96.250 214.880 ;
        RECT 90.760 192.360 90.930 193.090 ;
        RECT 90.710 191.450 91.120 192.360 ;
        RECT 96.050 191.920 96.220 193.310 ;
        RECT 101.210 191.450 101.680 214.930 ;
        RECT 204.880 214.860 205.220 215.810 ;
        RECT 210.240 214.900 210.410 215.450 ;
        RECT 215.400 215.190 215.740 216.260 ;
        RECT 225.910 216.200 239.500 216.310 ;
        RECT 215.400 214.930 215.770 215.190 ;
        RECT 220.820 214.930 220.990 215.450 ;
        RECT 80.080 191.000 102.330 191.450 ;
        RECT 80.140 190.970 102.330 191.000 ;
        RECT 90.710 190.860 91.120 190.970 ;
        RECT 74.700 187.650 75.160 187.700 ;
        RECT 85.340 187.650 85.680 187.730 ;
        RECT 95.960 187.650 96.300 187.810 ;
        RECT 74.700 187.600 96.300 187.650 ;
        RECT 74.130 187.380 96.300 187.600 ;
        RECT 74.130 187.200 96.340 187.380 ;
        RECT 74.130 187.150 95.580 187.200 ;
        RECT 74.700 185.750 75.160 187.150 ;
        RECT 80.180 185.790 80.350 186.340 ;
        RECT 85.340 186.080 85.680 187.150 ;
        RECT 85.340 185.820 85.710 186.080 ;
        RECT 90.760 185.820 90.930 186.340 ;
        RECT 74.700 158.530 75.140 185.750 ;
        RECT 80.160 163.980 80.390 185.790 ;
        RECT 85.420 164.090 85.650 185.820 ;
        RECT 80.180 163.420 80.350 163.980 ;
        RECT 80.080 162.370 80.490 163.420 ;
        RECT 85.470 162.840 85.640 164.090 ;
        RECT 90.760 164.010 90.990 185.820 ;
        RECT 95.920 185.800 96.340 187.200 ;
        RECT 96.020 164.230 96.250 185.800 ;
        RECT 90.760 163.280 90.930 164.010 ;
        RECT 90.710 162.370 91.120 163.280 ;
        RECT 96.050 162.840 96.220 164.230 ;
        RECT 101.210 163.650 101.680 190.970 ;
        RECT 101.210 162.370 101.900 163.650 ;
        RECT 80.080 161.920 102.330 162.370 ;
        RECT 80.140 161.890 102.330 161.920 ;
        RECT 90.710 161.780 91.120 161.890 ;
        RECT 74.700 158.480 75.160 158.530 ;
        RECT 85.340 158.480 85.680 158.560 ;
        RECT 95.960 158.480 96.300 158.640 ;
        RECT 74.700 158.430 96.300 158.480 ;
        RECT 74.130 158.210 96.300 158.430 ;
        RECT 74.130 158.030 96.340 158.210 ;
        RECT 74.130 157.980 95.580 158.030 ;
        RECT 74.700 156.580 75.160 157.980 ;
        RECT 80.180 156.620 80.350 157.170 ;
        RECT 85.340 156.910 85.680 157.980 ;
        RECT 85.340 156.650 85.710 156.910 ;
        RECT 90.760 156.650 90.930 157.170 ;
        RECT 74.700 129.350 75.140 156.580 ;
        RECT 80.160 134.810 80.390 156.620 ;
        RECT 85.420 134.920 85.650 156.650 ;
        RECT 80.180 134.250 80.350 134.810 ;
        RECT 80.080 133.200 80.490 134.250 ;
        RECT 85.470 133.670 85.640 134.920 ;
        RECT 90.760 134.840 90.990 156.650 ;
        RECT 95.920 156.630 96.340 158.030 ;
        RECT 96.020 135.060 96.250 156.630 ;
        RECT 101.210 156.610 101.900 161.890 ;
        RECT 90.760 134.110 90.930 134.840 ;
        RECT 90.710 133.200 91.120 134.110 ;
        RECT 96.050 133.670 96.220 135.060 ;
        RECT 101.210 134.320 101.680 156.610 ;
        RECT 101.200 133.200 101.860 134.320 ;
        RECT 80.080 132.750 102.330 133.200 ;
        RECT 80.140 132.720 102.330 132.750 ;
        RECT 90.710 132.610 91.120 132.720 ;
        RECT 74.700 129.300 75.160 129.350 ;
        RECT 85.340 129.300 85.680 129.380 ;
        RECT 95.960 129.300 96.300 129.460 ;
        RECT 74.700 129.250 96.300 129.300 ;
        RECT 74.130 129.030 96.300 129.250 ;
        RECT 74.130 128.850 96.340 129.030 ;
        RECT 74.130 128.800 95.580 128.850 ;
        RECT 74.700 127.400 75.160 128.800 ;
        RECT 80.180 127.440 80.350 127.990 ;
        RECT 85.340 127.730 85.680 128.800 ;
        RECT 85.340 127.470 85.710 127.730 ;
        RECT 90.760 127.470 90.930 127.990 ;
        RECT 74.700 100.030 75.140 127.400 ;
        RECT 80.160 105.630 80.390 127.440 ;
        RECT 85.420 105.740 85.650 127.470 ;
        RECT 80.180 105.070 80.350 105.630 ;
        RECT 80.080 104.020 80.490 105.070 ;
        RECT 85.470 104.490 85.640 105.740 ;
        RECT 90.760 105.660 90.990 127.470 ;
        RECT 95.920 127.450 96.340 128.850 ;
        RECT 96.020 105.880 96.250 127.450 ;
        RECT 101.200 127.280 101.860 132.720 ;
        RECT 90.760 104.930 90.930 105.660 ;
        RECT 90.710 104.020 91.120 104.930 ;
        RECT 96.050 104.490 96.220 105.880 ;
        RECT 101.210 104.020 101.680 127.280 ;
        RECT 80.080 103.570 102.330 104.020 ;
        RECT 80.140 103.540 102.330 103.570 ;
        RECT 90.710 103.430 91.120 103.540 ;
        RECT 74.700 99.980 75.160 100.030 ;
        RECT 85.340 99.980 85.680 100.060 ;
        RECT 95.960 99.980 96.300 100.140 ;
        RECT 74.700 99.930 96.300 99.980 ;
        RECT 74.130 99.710 96.300 99.930 ;
        RECT 74.130 99.530 96.340 99.710 ;
        RECT 74.130 99.480 95.580 99.530 ;
        RECT 74.700 98.080 75.160 99.480 ;
        RECT 80.180 98.120 80.350 98.670 ;
        RECT 85.340 98.410 85.680 99.480 ;
        RECT 85.340 98.150 85.710 98.410 ;
        RECT 90.760 98.150 90.930 98.670 ;
        RECT 74.700 70.750 75.140 98.080 ;
        RECT 80.160 76.310 80.390 98.120 ;
        RECT 85.420 76.420 85.650 98.150 ;
        RECT 80.180 75.750 80.350 76.310 ;
        RECT 80.080 74.700 80.490 75.750 ;
        RECT 85.470 75.170 85.640 76.420 ;
        RECT 90.760 76.340 90.990 98.150 ;
        RECT 95.920 98.130 96.340 99.530 ;
        RECT 96.020 76.560 96.250 98.130 ;
        RECT 90.760 75.610 90.930 76.340 ;
        RECT 90.710 74.700 91.120 75.610 ;
        RECT 96.050 75.170 96.220 76.560 ;
        RECT 101.210 74.700 101.680 103.540 ;
        RECT 80.080 74.250 102.330 74.700 ;
        RECT 80.140 74.220 102.330 74.250 ;
        RECT 90.710 74.110 91.120 74.220 ;
        RECT 74.700 70.700 75.210 70.750 ;
        RECT 85.390 70.700 85.730 70.780 ;
        RECT 96.010 70.700 96.350 70.860 ;
        RECT 74.700 70.650 96.350 70.700 ;
        RECT 74.180 70.430 96.350 70.650 ;
        RECT 74.180 70.250 96.390 70.430 ;
        RECT 74.180 70.200 95.630 70.250 ;
        RECT 74.700 68.800 75.210 70.200 ;
        RECT 80.230 68.840 80.400 69.390 ;
        RECT 85.390 69.130 85.730 70.200 ;
        RECT 85.390 68.870 85.760 69.130 ;
        RECT 90.810 68.870 90.980 69.390 ;
        RECT 74.700 46.200 75.140 68.800 ;
        RECT 80.210 47.030 80.440 68.840 ;
        RECT 85.470 47.140 85.700 68.870 ;
        RECT 80.230 46.470 80.400 47.030 ;
        RECT 74.700 41.160 75.360 46.200 ;
        RECT 80.130 45.420 80.540 46.470 ;
        RECT 85.520 45.890 85.690 47.140 ;
        RECT 90.810 47.060 91.040 68.870 ;
        RECT 95.970 68.850 96.390 70.250 ;
        RECT 96.070 47.280 96.300 68.850 ;
        RECT 90.810 46.330 90.980 47.060 ;
        RECT 90.760 45.420 91.170 46.330 ;
        RECT 96.100 45.890 96.270 47.280 ;
        RECT 101.210 46.130 101.680 74.220 ;
        RECT 101.210 45.420 101.900 46.130 ;
        RECT 80.130 44.970 102.380 45.420 ;
        RECT 80.190 44.940 102.380 44.970 ;
        RECT 90.760 44.830 91.170 44.940 ;
        RECT 85.480 41.160 85.820 41.240 ;
        RECT 96.100 41.160 96.440 41.320 ;
        RECT 74.700 41.110 96.440 41.160 ;
        RECT 74.270 40.890 96.440 41.110 ;
        RECT 74.270 40.710 96.480 40.890 ;
        RECT 74.270 40.660 95.720 40.710 ;
        RECT 74.700 39.160 75.360 40.660 ;
        RECT 80.320 39.300 80.490 39.850 ;
        RECT 85.480 39.590 85.820 40.660 ;
        RECT 85.480 39.330 85.850 39.590 ;
        RECT 90.900 39.330 91.070 39.850 ;
        RECT 74.960 38.230 75.200 39.160 ;
        RECT 74.960 34.380 75.190 38.230 ;
        RECT 74.960 32.760 75.200 34.380 ;
        RECT 74.960 28.910 75.190 32.760 ;
        RECT 74.960 27.290 75.200 28.910 ;
        RECT 74.960 23.440 75.190 27.290 ;
        RECT 74.960 21.820 75.200 23.440 ;
        RECT 74.960 17.970 75.190 21.820 ;
        RECT 74.960 17.600 75.200 17.970 ;
        RECT 68.830 15.840 69.240 16.860 ;
        RECT 75.030 16.350 75.200 17.600 ;
        RECT 80.300 17.490 80.530 39.300 ;
        RECT 85.560 17.600 85.790 39.330 ;
        RECT 80.320 16.930 80.490 17.490 ;
        RECT 80.220 15.880 80.630 16.930 ;
        RECT 85.610 16.350 85.780 17.600 ;
        RECT 90.900 17.520 91.130 39.330 ;
        RECT 96.060 39.310 96.480 40.710 ;
        RECT 96.160 17.740 96.390 39.310 ;
        RECT 101.210 39.170 101.900 44.940 ;
        RECT 101.240 39.090 101.900 39.170 ;
        RECT 90.900 16.790 91.070 17.520 ;
        RECT 90.850 15.880 91.260 16.790 ;
        RECT 96.190 16.350 96.360 17.740 ;
        RECT 101.440 17.600 101.670 39.090 ;
        RECT 102.800 17.910 106.000 209.470 ;
        RECT 135.410 17.650 138.440 213.850 ;
        RECT 167.950 18.940 171.390 214.110 ;
        RECT 204.880 213.830 205.120 214.860 ;
        RECT 200.460 27.940 203.690 212.830 ;
        RECT 204.880 209.980 205.110 213.830 ;
        RECT 204.880 208.360 205.120 209.980 ;
        RECT 204.880 204.510 205.110 208.360 ;
        RECT 204.880 202.890 205.120 204.510 ;
        RECT 204.880 199.040 205.110 202.890 ;
        RECT 204.880 197.420 205.120 199.040 ;
        RECT 204.880 193.570 205.110 197.420 ;
        RECT 204.880 193.200 205.120 193.570 ;
        RECT 204.950 192.980 205.120 193.200 ;
        RECT 210.220 193.090 210.450 214.900 ;
        RECT 215.480 193.200 215.710 214.930 ;
        RECT 204.810 187.680 205.440 192.980 ;
        RECT 210.240 192.530 210.410 193.090 ;
        RECT 210.140 191.480 210.550 192.530 ;
        RECT 215.530 191.950 215.700 193.200 ;
        RECT 220.820 193.120 221.050 214.930 ;
        RECT 225.980 214.910 226.400 216.200 ;
        RECT 226.080 193.340 226.310 214.910 ;
        RECT 231.280 212.770 231.930 216.200 ;
        RECT 237.820 214.970 238.160 216.200 ;
        RECT 243.180 215.010 243.350 215.560 ;
        RECT 248.340 215.300 248.680 216.370 ;
        RECT 258.890 216.310 272.480 216.420 ;
        RECT 248.340 215.040 248.710 215.300 ;
        RECT 253.760 215.040 253.930 215.560 ;
        RECT 237.820 213.940 238.060 214.970 ;
        RECT 220.820 192.390 220.990 193.120 ;
        RECT 220.770 191.480 221.180 192.390 ;
        RECT 226.110 191.950 226.280 193.340 ;
        RECT 231.360 193.200 231.590 212.770 ;
        RECT 231.400 192.560 231.570 193.200 ;
        RECT 231.210 191.480 231.840 192.560 ;
        RECT 210.140 191.030 232.390 191.480 ;
        RECT 210.200 191.000 232.390 191.030 ;
        RECT 220.770 190.890 221.180 191.000 ;
        RECT 215.400 187.680 215.740 187.760 ;
        RECT 226.020 187.680 226.360 187.840 ;
        RECT 204.810 187.630 226.360 187.680 ;
        RECT 204.190 187.410 226.360 187.630 ;
        RECT 204.190 187.230 226.400 187.410 ;
        RECT 204.190 187.180 225.640 187.230 ;
        RECT 204.810 186.060 205.440 187.180 ;
        RECT 204.880 185.780 205.220 186.060 ;
        RECT 210.240 185.820 210.410 186.370 ;
        RECT 215.400 186.110 215.740 187.180 ;
        RECT 215.400 185.850 215.770 186.110 ;
        RECT 220.820 185.850 220.990 186.370 ;
        RECT 204.880 184.750 205.120 185.780 ;
        RECT 204.880 180.900 205.110 184.750 ;
        RECT 204.880 179.280 205.120 180.900 ;
        RECT 204.880 175.430 205.110 179.280 ;
        RECT 204.880 173.810 205.120 175.430 ;
        RECT 204.880 169.960 205.110 173.810 ;
        RECT 204.880 168.340 205.120 169.960 ;
        RECT 204.880 164.490 205.110 168.340 ;
        RECT 204.880 164.120 205.120 164.490 ;
        RECT 204.950 163.510 205.120 164.120 ;
        RECT 210.220 164.010 210.450 185.820 ;
        RECT 215.480 164.120 215.710 185.850 ;
        RECT 204.810 158.510 205.440 163.510 ;
        RECT 210.240 163.450 210.410 164.010 ;
        RECT 210.140 162.400 210.550 163.450 ;
        RECT 215.530 162.870 215.700 164.120 ;
        RECT 220.820 164.040 221.050 185.850 ;
        RECT 225.980 185.830 226.400 187.230 ;
        RECT 226.080 164.260 226.310 185.830 ;
        RECT 231.210 185.640 231.840 191.000 ;
        RECT 220.820 163.310 220.990 164.040 ;
        RECT 220.770 162.400 221.180 163.310 ;
        RECT 226.110 162.870 226.280 164.260 ;
        RECT 231.360 164.120 231.590 185.640 ;
        RECT 231.400 163.420 231.570 164.120 ;
        RECT 231.280 163.160 231.690 163.420 ;
        RECT 231.210 162.400 231.840 163.160 ;
        RECT 210.140 161.950 232.390 162.400 ;
        RECT 210.200 161.920 232.390 161.950 ;
        RECT 220.770 161.810 221.180 161.920 ;
        RECT 215.400 158.510 215.740 158.590 ;
        RECT 226.020 158.510 226.360 158.670 ;
        RECT 204.810 158.460 226.360 158.510 ;
        RECT 204.190 158.240 226.360 158.460 ;
        RECT 204.190 158.060 226.400 158.240 ;
        RECT 204.190 158.010 225.640 158.060 ;
        RECT 204.810 156.590 205.440 158.010 ;
        RECT 210.240 156.650 210.410 157.200 ;
        RECT 215.400 156.940 215.740 158.010 ;
        RECT 215.400 156.680 215.770 156.940 ;
        RECT 220.820 156.680 220.990 157.200 ;
        RECT 204.880 155.580 205.120 156.590 ;
        RECT 204.880 151.730 205.110 155.580 ;
        RECT 204.880 150.110 205.120 151.730 ;
        RECT 204.880 146.260 205.110 150.110 ;
        RECT 204.880 144.640 205.120 146.260 ;
        RECT 204.880 140.790 205.110 144.640 ;
        RECT 204.880 139.170 205.120 140.790 ;
        RECT 204.880 135.320 205.110 139.170 ;
        RECT 204.880 134.950 205.120 135.320 ;
        RECT 204.950 134.180 205.120 134.950 ;
        RECT 210.220 134.840 210.450 156.650 ;
        RECT 215.480 134.950 215.710 156.680 ;
        RECT 210.240 134.280 210.410 134.840 ;
        RECT 204.810 129.330 205.440 134.180 ;
        RECT 210.140 133.230 210.550 134.280 ;
        RECT 215.530 133.700 215.700 134.950 ;
        RECT 220.820 134.870 221.050 156.680 ;
        RECT 225.980 156.660 226.400 158.060 ;
        RECT 226.080 135.090 226.310 156.660 ;
        RECT 231.210 156.240 231.840 161.920 ;
        RECT 220.820 134.140 220.990 134.870 ;
        RECT 220.770 133.230 221.180 134.140 ;
        RECT 226.110 133.700 226.280 135.090 ;
        RECT 231.360 134.950 231.590 156.240 ;
        RECT 231.400 134.320 231.570 134.950 ;
        RECT 231.210 133.230 231.840 134.320 ;
        RECT 210.140 132.780 232.390 133.230 ;
        RECT 210.200 132.750 232.390 132.780 ;
        RECT 220.770 132.640 221.180 132.750 ;
        RECT 215.400 129.330 215.740 129.410 ;
        RECT 226.020 129.330 226.360 129.490 ;
        RECT 204.810 129.280 226.360 129.330 ;
        RECT 204.190 129.060 226.360 129.280 ;
        RECT 204.190 128.880 226.400 129.060 ;
        RECT 204.190 128.830 225.640 128.880 ;
        RECT 204.810 127.260 205.440 128.830 ;
        RECT 210.240 127.470 210.410 128.020 ;
        RECT 215.400 127.760 215.740 128.830 ;
        RECT 215.400 127.500 215.770 127.760 ;
        RECT 220.820 127.500 220.990 128.020 ;
        RECT 204.880 126.400 205.120 127.260 ;
        RECT 204.880 122.550 205.110 126.400 ;
        RECT 204.880 120.930 205.120 122.550 ;
        RECT 204.880 117.080 205.110 120.930 ;
        RECT 204.880 115.460 205.120 117.080 ;
        RECT 204.880 111.610 205.110 115.460 ;
        RECT 204.880 109.990 205.120 111.610 ;
        RECT 204.880 106.140 205.110 109.990 ;
        RECT 204.880 105.770 205.120 106.140 ;
        RECT 204.950 105.540 205.120 105.770 ;
        RECT 210.220 105.660 210.450 127.470 ;
        RECT 215.480 105.770 215.710 127.500 ;
        RECT 204.740 100.010 205.370 105.540 ;
        RECT 210.240 105.100 210.410 105.660 ;
        RECT 210.140 104.050 210.550 105.100 ;
        RECT 215.530 104.520 215.700 105.770 ;
        RECT 220.820 105.690 221.050 127.500 ;
        RECT 225.980 127.480 226.400 128.880 ;
        RECT 226.080 105.910 226.310 127.480 ;
        RECT 231.210 127.400 231.840 132.750 ;
        RECT 220.820 104.960 220.990 105.690 ;
        RECT 220.770 104.050 221.180 104.960 ;
        RECT 226.110 104.520 226.280 105.910 ;
        RECT 231.360 105.770 231.590 127.400 ;
        RECT 231.400 105.070 231.570 105.770 ;
        RECT 231.280 104.990 231.690 105.070 ;
        RECT 231.210 104.050 231.840 104.990 ;
        RECT 210.140 103.600 232.390 104.050 ;
        RECT 210.200 103.570 232.390 103.600 ;
        RECT 220.770 103.460 221.180 103.570 ;
        RECT 215.400 100.010 215.740 100.090 ;
        RECT 226.020 100.010 226.360 100.170 ;
        RECT 204.740 99.960 226.360 100.010 ;
        RECT 204.190 99.740 226.360 99.960 ;
        RECT 204.190 99.560 226.400 99.740 ;
        RECT 204.190 99.510 225.640 99.560 ;
        RECT 204.740 98.620 205.370 99.510 ;
        RECT 204.880 98.110 205.220 98.620 ;
        RECT 210.240 98.150 210.410 98.700 ;
        RECT 215.400 98.440 215.740 99.510 ;
        RECT 215.400 98.180 215.770 98.440 ;
        RECT 220.820 98.180 220.990 98.700 ;
        RECT 204.880 97.080 205.120 98.110 ;
        RECT 204.880 93.230 205.110 97.080 ;
        RECT 204.880 91.610 205.120 93.230 ;
        RECT 204.880 87.760 205.110 91.610 ;
        RECT 204.880 86.140 205.120 87.760 ;
        RECT 204.880 82.290 205.110 86.140 ;
        RECT 204.880 80.670 205.120 82.290 ;
        RECT 204.880 76.820 205.110 80.670 ;
        RECT 204.880 76.450 205.120 76.820 ;
        RECT 204.950 76.280 205.120 76.450 ;
        RECT 210.220 76.340 210.450 98.150 ;
        RECT 215.480 76.450 215.710 98.180 ;
        RECT 204.880 70.730 205.510 76.280 ;
        RECT 210.240 75.780 210.410 76.340 ;
        RECT 210.140 74.730 210.550 75.780 ;
        RECT 215.530 75.200 215.700 76.450 ;
        RECT 220.820 76.370 221.050 98.180 ;
        RECT 225.980 98.160 226.400 99.560 ;
        RECT 226.080 76.590 226.310 98.160 ;
        RECT 231.210 98.070 231.840 103.570 ;
        RECT 220.820 75.640 220.990 76.370 ;
        RECT 220.770 74.730 221.180 75.640 ;
        RECT 226.110 75.200 226.280 76.590 ;
        RECT 231.360 76.450 231.590 98.070 ;
        RECT 231.400 75.750 231.570 76.450 ;
        RECT 231.280 75.160 231.690 75.750 ;
        RECT 231.280 74.730 231.910 75.160 ;
        RECT 210.140 74.280 232.390 74.730 ;
        RECT 210.200 74.250 232.390 74.280 ;
        RECT 220.770 74.140 221.180 74.250 ;
        RECT 215.450 70.730 215.790 70.810 ;
        RECT 226.070 70.730 226.410 70.890 ;
        RECT 204.880 70.680 226.410 70.730 ;
        RECT 204.240 70.460 226.410 70.680 ;
        RECT 204.240 70.280 226.450 70.460 ;
        RECT 204.240 70.230 225.690 70.280 ;
        RECT 204.880 69.360 205.510 70.230 ;
        RECT 204.930 68.830 205.270 69.360 ;
        RECT 210.290 68.870 210.460 69.420 ;
        RECT 215.450 69.160 215.790 70.230 ;
        RECT 215.450 68.900 215.820 69.160 ;
        RECT 220.870 68.900 221.040 69.420 ;
        RECT 204.930 67.800 205.170 68.830 ;
        RECT 204.930 63.950 205.160 67.800 ;
        RECT 204.930 62.330 205.170 63.950 ;
        RECT 204.930 58.480 205.160 62.330 ;
        RECT 204.930 56.860 205.170 58.480 ;
        RECT 204.930 53.010 205.160 56.860 ;
        RECT 204.930 51.390 205.170 53.010 ;
        RECT 204.930 47.540 205.160 51.390 ;
        RECT 204.930 47.170 205.170 47.540 ;
        RECT 205.000 46.950 205.170 47.170 ;
        RECT 210.270 47.060 210.500 68.870 ;
        RECT 215.530 47.170 215.760 68.900 ;
        RECT 204.740 41.190 205.370 46.950 ;
        RECT 210.290 46.500 210.460 47.060 ;
        RECT 210.190 45.450 210.600 46.500 ;
        RECT 215.580 45.920 215.750 47.170 ;
        RECT 220.870 47.090 221.100 68.900 ;
        RECT 226.030 68.880 226.450 70.280 ;
        RECT 226.130 47.310 226.360 68.880 ;
        RECT 231.280 68.240 231.910 74.250 ;
        RECT 220.870 46.360 221.040 47.090 ;
        RECT 220.820 45.450 221.230 46.360 ;
        RECT 226.160 45.920 226.330 47.310 ;
        RECT 231.410 47.170 231.640 68.240 ;
        RECT 231.450 46.470 231.620 47.170 ;
        RECT 231.330 45.550 231.740 46.470 ;
        RECT 231.280 45.450 231.910 45.550 ;
        RECT 210.190 45.000 232.440 45.450 ;
        RECT 210.250 44.970 232.440 45.000 ;
        RECT 220.820 44.860 221.230 44.970 ;
        RECT 215.540 41.190 215.880 41.270 ;
        RECT 226.160 41.190 226.500 41.350 ;
        RECT 204.740 41.140 226.500 41.190 ;
        RECT 204.330 40.920 226.500 41.140 ;
        RECT 204.330 40.740 226.540 40.920 ;
        RECT 204.330 40.690 225.780 40.740 ;
        RECT 204.740 40.030 205.370 40.690 ;
        RECT 205.020 39.290 205.360 40.030 ;
        RECT 210.380 39.330 210.550 39.880 ;
        RECT 215.540 39.620 215.880 40.690 ;
        RECT 215.540 39.360 215.910 39.620 ;
        RECT 220.960 39.360 221.130 39.880 ;
        RECT 205.020 38.260 205.260 39.290 ;
        RECT 205.020 34.410 205.250 38.260 ;
        RECT 205.020 32.790 205.260 34.410 ;
        RECT 205.020 28.940 205.250 32.790 ;
        RECT 101.480 16.900 101.650 17.600 ;
        RECT 101.360 15.880 101.770 16.900 ;
        RECT 15.120 15.350 37.370 15.800 ;
        RECT 47.690 15.390 69.940 15.840 ;
        RECT 80.220 15.430 102.470 15.880 ;
        RECT 80.280 15.400 102.470 15.430 ;
        RECT 47.750 15.360 69.940 15.390 ;
        RECT 15.180 15.320 37.370 15.350 ;
        RECT 25.750 15.210 26.160 15.320 ;
        RECT 58.320 15.250 58.730 15.360 ;
        RECT 90.850 15.290 91.260 15.400 ;
        RECT -96.355 11.870 -71.855 11.905 ;
        RECT -96.690 11.700 -71.600 11.870 ;
        RECT -96.355 11.655 -71.855 11.700 ;
        RECT -81.615 11.300 -81.445 11.655 ;
        RECT -90.700 11.180 -77.210 11.300 ;
        RECT -90.810 11.010 -77.210 11.180 ;
        RECT -90.700 8.680 -77.210 11.010 ;
        RECT 201.610 -2.480 202.830 27.940 ;
        RECT 205.020 27.320 205.260 28.940 ;
        RECT 205.020 23.470 205.250 27.320 ;
        RECT 205.020 21.850 205.260 23.470 ;
        RECT 205.020 18.000 205.250 21.850 ;
        RECT 205.020 17.630 205.260 18.000 ;
        RECT 205.090 16.380 205.260 17.630 ;
        RECT 210.360 17.520 210.590 39.330 ;
        RECT 215.620 17.630 215.850 39.360 ;
        RECT 210.380 16.960 210.550 17.520 ;
        RECT 210.280 15.910 210.690 16.960 ;
        RECT 215.670 16.380 215.840 17.630 ;
        RECT 220.960 17.550 221.190 39.360 ;
        RECT 226.120 39.340 226.540 40.740 ;
        RECT 226.220 17.770 226.450 39.340 ;
        RECT 231.280 38.630 231.910 44.970 ;
        RECT 220.960 16.820 221.130 17.550 ;
        RECT 220.910 15.910 221.320 16.820 ;
        RECT 226.250 16.380 226.420 17.770 ;
        RECT 231.500 17.630 231.730 38.630 ;
        RECT 232.980 27.030 236.460 212.120 ;
        RECT 237.820 210.090 238.050 213.940 ;
        RECT 237.820 208.470 238.060 210.090 ;
        RECT 237.820 204.620 238.050 208.470 ;
        RECT 237.820 203.000 238.060 204.620 ;
        RECT 237.820 199.150 238.050 203.000 ;
        RECT 237.820 197.530 238.060 199.150 ;
        RECT 237.820 193.680 238.050 197.530 ;
        RECT 237.820 193.310 238.060 193.680 ;
        RECT 237.890 193.020 238.060 193.310 ;
        RECT 243.160 193.200 243.390 215.010 ;
        RECT 248.420 193.310 248.650 215.040 ;
        RECT 237.740 187.790 238.400 193.020 ;
        RECT 243.180 192.640 243.350 193.200 ;
        RECT 243.080 191.590 243.490 192.640 ;
        RECT 248.470 192.060 248.640 193.310 ;
        RECT 253.760 193.230 253.990 215.040 ;
        RECT 258.920 215.020 259.340 216.310 ;
        RECT 259.020 193.450 259.250 215.020 ;
        RECT 264.150 212.870 264.800 216.310 ;
        RECT 270.390 215.040 270.730 216.310 ;
        RECT 275.750 215.080 275.920 215.630 ;
        RECT 280.910 215.370 281.250 216.440 ;
        RECT 291.480 215.990 297.230 216.490 ;
        RECT 312.490 216.420 312.800 216.470 ;
        RECT 280.910 215.110 281.280 215.370 ;
        RECT 286.330 215.110 286.500 215.630 ;
        RECT 270.390 214.010 270.630 215.040 ;
        RECT 253.760 192.500 253.930 193.230 ;
        RECT 253.710 191.590 254.120 192.500 ;
        RECT 259.050 192.060 259.220 193.450 ;
        RECT 264.300 193.310 264.530 212.870 ;
        RECT 264.340 192.680 264.510 193.310 ;
        RECT 264.250 192.610 264.730 192.680 ;
        RECT 264.220 191.590 264.730 192.610 ;
        RECT 243.080 191.140 265.330 191.590 ;
        RECT 243.140 191.110 265.330 191.140 ;
        RECT 253.710 191.000 254.120 191.110 ;
        RECT 248.340 187.790 248.680 187.870 ;
        RECT 258.960 187.790 259.300 187.950 ;
        RECT 237.740 187.740 259.300 187.790 ;
        RECT 237.130 187.520 259.300 187.740 ;
        RECT 237.130 187.340 259.340 187.520 ;
        RECT 237.130 187.290 258.580 187.340 ;
        RECT 237.740 185.980 238.400 187.290 ;
        RECT 237.820 185.890 238.160 185.980 ;
        RECT 243.180 185.930 243.350 186.480 ;
        RECT 248.340 186.220 248.680 187.290 ;
        RECT 248.340 185.960 248.710 186.220 ;
        RECT 253.760 185.960 253.930 186.480 ;
        RECT 237.820 184.860 238.060 185.890 ;
        RECT 237.820 181.010 238.050 184.860 ;
        RECT 237.820 179.390 238.060 181.010 ;
        RECT 237.820 175.540 238.050 179.390 ;
        RECT 237.820 173.920 238.060 175.540 ;
        RECT 237.820 170.070 238.050 173.920 ;
        RECT 237.820 168.450 238.060 170.070 ;
        RECT 237.820 164.600 238.050 168.450 ;
        RECT 237.820 164.230 238.060 164.600 ;
        RECT 237.890 163.950 238.060 164.230 ;
        RECT 243.160 164.120 243.390 185.930 ;
        RECT 248.420 164.230 248.650 185.960 ;
        RECT 237.620 158.620 238.280 163.950 ;
        RECT 243.180 163.560 243.350 164.120 ;
        RECT 243.080 162.510 243.490 163.560 ;
        RECT 248.470 162.980 248.640 164.230 ;
        RECT 253.760 164.150 253.990 185.960 ;
        RECT 258.920 185.940 259.340 187.340 ;
        RECT 264.250 185.990 264.730 191.110 ;
        RECT 259.020 164.370 259.250 185.940 ;
        RECT 253.760 163.420 253.930 164.150 ;
        RECT 253.710 162.510 254.120 163.420 ;
        RECT 259.050 162.980 259.220 164.370 ;
        RECT 264.300 164.230 264.530 185.990 ;
        RECT 264.340 163.530 264.510 164.230 ;
        RECT 264.220 163.510 264.630 163.530 ;
        RECT 264.210 162.510 264.690 163.510 ;
        RECT 243.080 162.060 265.330 162.510 ;
        RECT 243.140 162.030 265.330 162.060 ;
        RECT 253.710 161.920 254.120 162.030 ;
        RECT 248.340 158.620 248.680 158.700 ;
        RECT 258.960 158.620 259.300 158.780 ;
        RECT 237.620 158.570 259.300 158.620 ;
        RECT 237.130 158.350 259.300 158.570 ;
        RECT 237.130 158.170 259.340 158.350 ;
        RECT 237.130 158.120 258.580 158.170 ;
        RECT 237.620 156.910 238.280 158.120 ;
        RECT 237.820 156.720 238.160 156.910 ;
        RECT 243.180 156.760 243.350 157.310 ;
        RECT 248.340 157.050 248.680 158.120 ;
        RECT 248.340 156.790 248.710 157.050 ;
        RECT 253.760 156.790 253.930 157.310 ;
        RECT 237.820 155.690 238.060 156.720 ;
        RECT 237.820 151.840 238.050 155.690 ;
        RECT 237.820 150.220 238.060 151.840 ;
        RECT 237.820 146.370 238.050 150.220 ;
        RECT 237.820 144.750 238.060 146.370 ;
        RECT 237.820 140.900 238.050 144.750 ;
        RECT 237.820 139.280 238.060 140.900 ;
        RECT 237.820 135.470 238.050 139.280 ;
        RECT 237.700 129.440 238.360 135.470 ;
        RECT 243.160 134.950 243.390 156.760 ;
        RECT 248.420 135.060 248.650 156.790 ;
        RECT 243.180 134.390 243.350 134.950 ;
        RECT 243.080 133.340 243.490 134.390 ;
        RECT 248.470 133.810 248.640 135.060 ;
        RECT 253.760 134.980 253.990 156.790 ;
        RECT 258.920 156.770 259.340 158.170 ;
        RECT 264.210 156.820 264.690 162.030 ;
        RECT 259.020 135.200 259.250 156.770 ;
        RECT 253.760 134.250 253.930 134.980 ;
        RECT 253.710 133.340 254.120 134.250 ;
        RECT 259.050 133.810 259.220 135.200 ;
        RECT 264.300 135.060 264.530 156.820 ;
        RECT 264.340 134.360 264.510 135.060 ;
        RECT 264.220 134.200 264.630 134.360 ;
        RECT 264.180 133.340 264.660 134.200 ;
        RECT 243.080 132.890 265.330 133.340 ;
        RECT 243.140 132.860 265.330 132.890 ;
        RECT 253.710 132.750 254.120 132.860 ;
        RECT 248.340 129.440 248.680 129.520 ;
        RECT 258.960 129.440 259.300 129.600 ;
        RECT 237.700 129.390 259.300 129.440 ;
        RECT 237.130 129.170 259.300 129.390 ;
        RECT 237.130 128.990 259.340 129.170 ;
        RECT 237.130 128.940 258.580 128.990 ;
        RECT 237.700 128.430 238.360 128.940 ;
        RECT 237.820 127.540 238.160 128.430 ;
        RECT 243.180 127.580 243.350 128.130 ;
        RECT 248.340 127.870 248.680 128.940 ;
        RECT 248.340 127.610 248.710 127.870 ;
        RECT 253.760 127.610 253.930 128.130 ;
        RECT 237.820 126.510 238.060 127.540 ;
        RECT 237.820 122.660 238.050 126.510 ;
        RECT 237.820 121.040 238.060 122.660 ;
        RECT 237.820 117.190 238.050 121.040 ;
        RECT 237.820 115.570 238.060 117.190 ;
        RECT 237.820 111.720 238.050 115.570 ;
        RECT 237.820 110.100 238.060 111.720 ;
        RECT 237.820 106.250 238.050 110.100 ;
        RECT 237.820 105.880 238.060 106.250 ;
        RECT 237.890 105.470 238.060 105.880 ;
        RECT 243.160 105.770 243.390 127.580 ;
        RECT 248.420 105.880 248.650 127.610 ;
        RECT 237.740 100.120 238.400 105.470 ;
        RECT 243.180 105.210 243.350 105.770 ;
        RECT 243.080 104.160 243.490 105.210 ;
        RECT 248.470 104.630 248.640 105.880 ;
        RECT 253.760 105.800 253.990 127.610 ;
        RECT 258.920 127.590 259.340 128.990 ;
        RECT 259.020 106.020 259.250 127.590 ;
        RECT 264.180 127.510 264.660 132.860 ;
        RECT 253.760 105.070 253.930 105.800 ;
        RECT 253.710 104.160 254.120 105.070 ;
        RECT 259.050 104.630 259.220 106.020 ;
        RECT 264.300 105.880 264.530 127.510 ;
        RECT 264.340 105.180 264.510 105.880 ;
        RECT 264.220 104.850 264.630 105.180 ;
        RECT 264.220 104.160 264.770 104.850 ;
        RECT 243.080 103.710 265.330 104.160 ;
        RECT 243.140 103.680 265.330 103.710 ;
        RECT 253.710 103.570 254.120 103.680 ;
        RECT 248.340 100.120 248.680 100.200 ;
        RECT 258.960 100.120 259.300 100.280 ;
        RECT 237.740 100.070 259.300 100.120 ;
        RECT 237.130 99.850 259.300 100.070 ;
        RECT 237.130 99.670 259.340 99.850 ;
        RECT 237.130 99.620 258.580 99.670 ;
        RECT 237.740 98.430 238.400 99.620 ;
        RECT 237.820 98.220 238.160 98.430 ;
        RECT 243.180 98.260 243.350 98.810 ;
        RECT 248.340 98.550 248.680 99.620 ;
        RECT 248.340 98.290 248.710 98.550 ;
        RECT 253.760 98.290 253.930 98.810 ;
        RECT 237.820 97.190 238.060 98.220 ;
        RECT 237.820 93.340 238.050 97.190 ;
        RECT 237.820 91.720 238.060 93.340 ;
        RECT 237.820 87.870 238.050 91.720 ;
        RECT 237.820 86.250 238.060 87.870 ;
        RECT 237.820 82.400 238.050 86.250 ;
        RECT 237.820 80.780 238.060 82.400 ;
        RECT 237.820 76.930 238.050 80.780 ;
        RECT 237.820 76.560 238.060 76.930 ;
        RECT 237.890 76.380 238.060 76.560 ;
        RECT 243.160 76.450 243.390 98.260 ;
        RECT 248.420 76.560 248.650 98.290 ;
        RECT 237.640 70.840 238.270 76.380 ;
        RECT 243.180 75.890 243.350 76.450 ;
        RECT 243.080 74.840 243.490 75.890 ;
        RECT 248.470 75.310 248.640 76.560 ;
        RECT 253.760 76.480 253.990 98.290 ;
        RECT 258.920 98.270 259.340 99.670 ;
        RECT 259.020 76.700 259.250 98.270 ;
        RECT 264.290 98.160 264.770 103.680 ;
        RECT 253.760 75.750 253.930 76.480 ;
        RECT 253.710 74.840 254.120 75.750 ;
        RECT 259.050 75.310 259.220 76.700 ;
        RECT 264.300 76.660 264.530 98.160 ;
        RECT 264.150 74.840 264.780 76.660 ;
        RECT 243.080 74.390 265.330 74.840 ;
        RECT 243.140 74.360 265.330 74.390 ;
        RECT 253.710 74.250 254.120 74.360 ;
        RECT 248.390 70.840 248.730 70.920 ;
        RECT 259.010 70.840 259.350 71.000 ;
        RECT 237.640 70.790 259.350 70.840 ;
        RECT 237.180 70.570 259.350 70.790 ;
        RECT 237.180 70.390 259.390 70.570 ;
        RECT 237.180 70.340 258.630 70.390 ;
        RECT 237.640 69.460 238.270 70.340 ;
        RECT 237.870 68.940 238.210 69.460 ;
        RECT 243.230 68.980 243.400 69.530 ;
        RECT 248.390 69.270 248.730 70.340 ;
        RECT 248.390 69.010 248.760 69.270 ;
        RECT 253.810 69.010 253.980 69.530 ;
        RECT 237.870 67.910 238.110 68.940 ;
        RECT 237.870 64.060 238.100 67.910 ;
        RECT 237.870 62.440 238.110 64.060 ;
        RECT 237.870 58.590 238.100 62.440 ;
        RECT 237.870 56.970 238.110 58.590 ;
        RECT 237.870 53.120 238.100 56.970 ;
        RECT 237.870 51.500 238.110 53.120 ;
        RECT 237.870 47.650 238.100 51.500 ;
        RECT 237.870 47.280 238.110 47.650 ;
        RECT 237.940 46.990 238.110 47.280 ;
        RECT 243.210 47.170 243.440 68.980 ;
        RECT 248.470 47.280 248.700 69.010 ;
        RECT 237.710 41.300 238.340 46.990 ;
        RECT 243.230 46.610 243.400 47.170 ;
        RECT 243.130 45.560 243.540 46.610 ;
        RECT 248.520 46.030 248.690 47.280 ;
        RECT 253.810 47.200 254.040 69.010 ;
        RECT 258.970 68.990 259.390 70.390 ;
        RECT 264.150 69.740 264.780 74.360 ;
        RECT 264.390 69.090 264.560 69.530 ;
        RECT 259.070 47.420 259.300 68.990 ;
        RECT 253.810 46.470 253.980 47.200 ;
        RECT 253.760 45.560 254.170 46.470 ;
        RECT 259.100 46.030 259.270 47.420 ;
        RECT 264.350 47.280 264.580 69.090 ;
        RECT 264.390 46.580 264.560 47.280 ;
        RECT 264.270 45.870 264.680 46.580 ;
        RECT 264.270 45.560 264.990 45.870 ;
        RECT 243.130 45.110 265.380 45.560 ;
        RECT 243.190 45.080 265.380 45.110 ;
        RECT 253.760 44.970 254.170 45.080 ;
        RECT 248.480 41.300 248.820 41.380 ;
        RECT 259.100 41.300 259.440 41.460 ;
        RECT 237.710 41.250 259.440 41.300 ;
        RECT 237.270 41.030 259.440 41.250 ;
        RECT 237.270 40.850 259.480 41.030 ;
        RECT 237.270 40.800 258.720 40.850 ;
        RECT 237.710 40.070 238.340 40.800 ;
        RECT 237.960 39.400 238.300 40.070 ;
        RECT 243.320 39.440 243.490 39.990 ;
        RECT 248.480 39.730 248.820 40.800 ;
        RECT 248.480 39.470 248.850 39.730 ;
        RECT 253.900 39.470 254.070 39.990 ;
        RECT 237.960 38.370 238.200 39.400 ;
        RECT 237.960 34.520 238.190 38.370 ;
        RECT 237.960 32.900 238.200 34.520 ;
        RECT 237.960 29.050 238.190 32.900 ;
        RECT 237.960 27.430 238.200 29.050 ;
        RECT 234.760 24.640 235.510 27.030 ;
        RECT 237.960 23.580 238.190 27.430 ;
        RECT 237.960 21.960 238.200 23.580 ;
        RECT 237.960 18.110 238.190 21.960 ;
        RECT 237.960 17.740 238.200 18.110 ;
        RECT 231.540 16.930 231.710 17.630 ;
        RECT 231.420 16.240 231.830 16.930 ;
        RECT 238.030 16.490 238.200 17.740 ;
        RECT 243.300 17.630 243.530 39.440 ;
        RECT 248.560 17.740 248.790 39.470 ;
        RECT 243.320 17.070 243.490 17.630 ;
        RECT 243.220 16.240 243.630 17.070 ;
        RECT 248.610 16.490 248.780 17.740 ;
        RECT 253.900 17.660 254.130 39.470 ;
        RECT 259.060 39.450 259.480 40.850 ;
        RECT 259.160 17.880 259.390 39.450 ;
        RECT 264.360 38.950 264.990 45.080 ;
        RECT 253.900 16.930 254.070 17.660 ;
        RECT 253.850 16.240 254.260 16.930 ;
        RECT 259.190 16.490 259.360 17.880 ;
        RECT 264.440 17.740 264.670 38.950 ;
        RECT 265.680 26.880 269.160 211.970 ;
        RECT 270.390 210.160 270.620 214.010 ;
        RECT 270.390 208.540 270.630 210.160 ;
        RECT 270.390 204.690 270.620 208.540 ;
        RECT 270.390 203.070 270.630 204.690 ;
        RECT 270.390 199.220 270.620 203.070 ;
        RECT 270.390 197.600 270.630 199.220 ;
        RECT 270.390 193.750 270.620 197.600 ;
        RECT 270.390 193.380 270.630 193.750 ;
        RECT 270.460 193.010 270.630 193.380 ;
        RECT 275.730 193.270 275.960 215.080 ;
        RECT 280.990 193.380 281.220 215.110 ;
        RECT 270.310 187.860 270.790 193.010 ;
        RECT 275.750 192.710 275.920 193.270 ;
        RECT 275.650 191.660 276.060 192.710 ;
        RECT 281.040 192.130 281.210 193.380 ;
        RECT 286.330 193.300 286.560 215.110 ;
        RECT 291.490 215.090 291.910 215.990 ;
        RECT 291.590 193.520 291.820 215.090 ;
        RECT 296.740 214.320 297.230 215.990 ;
        RECT 312.390 216.340 312.800 216.420 ;
        RECT 319.210 216.380 319.960 217.220 ;
        RECT 328.880 216.410 329.250 216.430 ;
        RECT 319.080 216.360 319.960 216.380 ;
        RECT 319.040 216.340 319.960 216.360 ;
        RECT 325.330 216.340 329.300 216.410 ;
        RECT 312.390 215.960 329.300 216.340 ;
        RECT 312.390 214.820 312.800 215.960 ;
        RECT 315.830 215.180 316.000 215.620 ;
        RECT 286.330 192.570 286.500 193.300 ;
        RECT 286.280 191.660 286.690 192.570 ;
        RECT 291.620 192.130 291.790 193.520 ;
        RECT 296.870 193.380 297.100 214.320 ;
        RECT 297.650 200.330 299.670 209.760 ;
        RECT 310.740 203.950 311.800 213.500 ;
        RECT 312.490 201.330 312.780 214.820 ;
        RECT 315.780 201.350 316.070 215.180 ;
        RECT 319.040 214.760 319.390 215.960 ;
        RECT 325.330 215.820 329.300 215.960 ;
        RECT 322.410 215.360 322.580 215.620 ;
        RECT 319.040 201.350 319.330 214.760 ;
        RECT 322.350 201.530 322.640 215.360 ;
        RECT 325.550 214.450 326.020 215.820 ;
        RECT 328.880 215.270 329.250 215.820 ;
        RECT 328.870 215.040 329.270 215.270 ;
        RECT 334.800 215.190 334.970 215.630 ;
        RECT 341.380 215.370 341.550 215.630 ;
        RECT 312.540 200.720 312.710 201.330 ;
        RECT 315.790 200.360 316.060 201.350 ;
        RECT 319.120 200.720 319.290 201.350 ;
        RECT 322.410 201.340 322.580 201.530 ;
        RECT 325.620 201.370 325.910 214.450 ;
        RECT 328.940 213.320 329.230 215.040 ;
        RECT 329.430 213.320 331.010 214.590 ;
        RECT 328.940 212.720 331.010 213.320 ;
        RECT 322.380 200.360 322.650 201.340 ;
        RECT 325.700 200.720 325.870 201.370 ;
        RECT 328.940 201.360 329.230 212.720 ;
        RECT 329.430 212.240 331.010 212.720 ;
        RECT 329.710 203.960 330.770 212.240 ;
        RECT 334.750 201.360 335.040 215.190 ;
        RECT 341.320 201.540 341.610 215.370 ;
        RECT 347.890 214.580 348.740 217.740 ;
        RECT 357.850 217.130 359.390 218.190 ;
        RECT 350.500 216.500 350.810 216.550 ;
        RECT 350.400 216.420 350.810 216.500 ;
        RECT 357.090 216.440 357.400 216.460 ;
        RECT 357.050 216.420 357.400 216.440 ;
        RECT 358.280 216.420 358.940 217.130 ;
        RECT 363.560 216.430 364.030 216.440 ;
        RECT 366.820 216.430 367.280 216.440 ;
        RECT 363.560 216.420 367.300 216.430 ;
        RECT 350.400 216.040 367.300 216.420 ;
        RECT 350.400 214.900 350.810 216.040 ;
        RECT 353.840 215.260 354.010 215.700 ;
        RECT 347.910 209.480 348.200 214.580 ;
        RECT 348.750 209.480 349.810 213.580 ;
        RECT 347.840 208.950 349.810 209.480 ;
        RECT 328.920 201.240 329.230 201.360 ;
        RECT 328.920 200.360 329.190 201.240 ;
        RECT 334.760 200.370 335.030 201.360 ;
        RECT 341.380 201.350 341.550 201.540 ;
        RECT 347.910 201.370 348.200 208.950 ;
        RECT 348.750 204.030 349.810 208.950 ;
        RECT 350.500 201.410 350.790 214.900 ;
        RECT 353.790 201.430 354.080 215.260 ;
        RECT 357.050 214.840 357.400 216.040 ;
        RECT 358.280 216.010 358.940 216.040 ;
        RECT 363.560 215.960 367.300 216.040 ;
        RECT 360.420 215.440 360.590 215.700 ;
        RECT 357.050 201.430 357.340 214.840 ;
        RECT 360.360 201.610 360.650 215.440 ;
        RECT 363.560 214.530 364.030 215.960 ;
        RECT 366.820 215.400 367.280 215.960 ;
        RECT 366.820 215.170 367.300 215.400 ;
        RECT 366.870 214.710 367.300 215.170 ;
        RECT 341.350 200.370 341.620 201.350 ;
        RECT 347.890 201.250 348.200 201.370 ;
        RECT 347.890 200.370 348.160 201.250 ;
        RECT 350.550 200.800 350.720 201.410 ;
        RECT 353.800 200.440 354.070 201.430 ;
        RECT 357.130 200.800 357.300 201.430 ;
        RECT 360.420 201.420 360.590 201.610 ;
        RECT 363.630 201.450 363.920 214.530 ;
        RECT 366.950 214.480 367.240 214.710 ;
        RECT 368.050 214.480 369.750 215.010 ;
        RECT 366.950 213.930 369.750 214.480 ;
        RECT 360.390 200.440 360.660 201.420 ;
        RECT 363.710 200.800 363.880 201.450 ;
        RECT 366.950 201.440 367.240 213.930 ;
        RECT 368.050 203.340 369.750 213.930 ;
        RECT 366.930 201.320 367.240 201.440 ;
        RECT 366.930 200.440 367.200 201.320 ;
        RECT 315.710 199.870 329.230 200.360 ;
        RECT 334.680 199.880 348.200 200.370 ;
        RECT 353.720 199.950 367.240 200.440 ;
        RECT 360.390 199.930 360.660 199.950 ;
        RECT 322.380 199.850 322.650 199.870 ;
        RECT 341.350 199.860 341.620 199.880 ;
        RECT 385.440 196.270 386.210 196.990 ;
        RECT 392.480 196.930 394.170 197.640 ;
        RECT 425.140 197.010 426.860 197.710 ;
        RECT 392.380 196.270 392.690 196.320 ;
        RECT 392.870 196.270 393.530 196.930 ;
        RECT 395.500 196.270 396.160 196.470 ;
        RECT 398.880 196.270 399.190 196.420 ;
        RECT 385.440 196.000 399.300 196.270 ;
        RECT 418.620 196.240 419.390 196.960 ;
        RECT 425.470 196.240 426.270 197.010 ;
        RECT 428.740 196.240 429.350 196.300 ;
        RECT 432.060 196.240 432.370 196.390 ;
        RECT 385.440 195.800 386.210 196.000 ;
        RECT 296.910 192.680 297.080 193.380 ;
        RECT 296.790 192.350 297.200 192.680 ;
        RECT 296.710 191.660 297.200 192.350 ;
        RECT 275.650 191.210 297.900 191.660 ;
        RECT 275.710 191.180 297.900 191.210 ;
        RECT 286.280 191.070 286.690 191.180 ;
        RECT 280.910 187.860 281.250 187.940 ;
        RECT 291.530 187.860 291.870 188.020 ;
        RECT 270.310 187.810 291.870 187.860 ;
        RECT 269.700 187.590 291.870 187.810 ;
        RECT 269.700 187.410 291.910 187.590 ;
        RECT 269.700 187.360 291.150 187.410 ;
        RECT 270.310 186.320 270.790 187.360 ;
        RECT 270.390 185.960 270.730 186.320 ;
        RECT 275.750 186.000 275.920 186.550 ;
        RECT 280.910 186.290 281.250 187.360 ;
        RECT 280.910 186.030 281.280 186.290 ;
        RECT 286.330 186.030 286.500 186.550 ;
        RECT 270.390 184.930 270.630 185.960 ;
        RECT 270.390 181.080 270.620 184.930 ;
        RECT 270.390 179.460 270.630 181.080 ;
        RECT 270.390 175.610 270.620 179.460 ;
        RECT 270.390 173.990 270.630 175.610 ;
        RECT 270.390 170.140 270.620 173.990 ;
        RECT 270.390 168.520 270.630 170.140 ;
        RECT 270.390 164.670 270.620 168.520 ;
        RECT 270.390 164.300 270.630 164.670 ;
        RECT 270.460 164.030 270.630 164.300 ;
        RECT 275.730 164.190 275.960 186.000 ;
        RECT 280.990 164.300 281.220 186.030 ;
        RECT 270.060 163.290 270.720 164.030 ;
        RECT 275.750 163.630 275.920 164.190 ;
        RECT 270.060 158.690 270.870 163.290 ;
        RECT 275.650 162.580 276.060 163.630 ;
        RECT 281.040 163.050 281.210 164.300 ;
        RECT 286.330 164.220 286.560 186.030 ;
        RECT 291.490 186.010 291.910 187.410 ;
        RECT 291.590 164.440 291.820 186.010 ;
        RECT 296.710 185.660 297.190 191.180 ;
        RECT 286.330 163.490 286.500 164.220 ;
        RECT 286.280 162.580 286.690 163.490 ;
        RECT 291.620 163.050 291.790 164.440 ;
        RECT 296.870 164.300 297.100 185.660 ;
        RECT 298.000 170.780 300.010 180.420 ;
        RECT 383.170 177.650 384.890 195.410 ;
        RECT 385.720 195.260 386.030 195.800 ;
        RECT 385.720 195.030 386.050 195.260 ;
        RECT 389.140 195.160 389.310 195.550 ;
        RECT 385.800 177.620 386.030 195.030 ;
        RECT 389.100 177.700 389.330 195.160 ;
        RECT 392.380 195.150 392.690 196.000 ;
        RECT 392.870 195.970 393.530 196.000 ;
        RECT 392.390 177.700 392.620 195.150 ;
        RECT 395.500 194.990 396.160 196.000 ;
        RECT 398.880 195.430 399.190 196.000 ;
        RECT 418.620 195.970 432.480 196.240 ;
        RECT 418.620 195.770 419.390 195.970 ;
        RECT 425.470 195.930 426.270 195.970 ;
        RECT 398.880 195.070 399.220 195.430 ;
        RECT 395.690 177.760 395.920 194.990 ;
        RECT 398.990 193.830 399.220 195.070 ;
        RECT 399.800 193.830 401.520 195.380 ;
        RECT 405.770 195.130 405.940 195.520 ;
        RECT 412.350 195.190 412.520 195.520 ;
        RECT 398.970 193.350 401.520 193.830 ;
        RECT 398.990 177.780 399.220 193.350 ;
        RECT 385.850 177.180 386.020 177.620 ;
        RECT 389.140 177.520 389.310 177.700 ;
        RECT 389.040 176.660 389.350 177.520 ;
        RECT 392.430 177.180 392.600 177.700 ;
        RECT 395.720 177.480 395.890 177.760 ;
        RECT 395.600 176.660 395.910 177.480 ;
        RECT 399.010 177.180 399.180 177.780 ;
        RECT 399.800 177.620 401.520 193.350 ;
        RECT 405.730 177.670 405.960 195.130 ;
        RECT 412.320 177.730 412.550 195.190 ;
        RECT 405.770 177.490 405.940 177.670 ;
        RECT 389.040 176.350 395.960 176.660 ;
        RECT 389.100 176.330 395.960 176.350 ;
        RECT 405.670 176.630 405.980 177.490 ;
        RECT 412.350 177.450 412.520 177.730 ;
        RECT 416.350 177.620 418.070 195.380 ;
        RECT 418.900 195.230 419.210 195.770 ;
        RECT 418.900 195.000 419.230 195.230 ;
        RECT 422.320 195.130 422.490 195.520 ;
        RECT 418.980 177.590 419.210 195.000 ;
        RECT 422.280 177.670 422.510 195.130 ;
        RECT 425.560 195.120 425.870 195.930 ;
        RECT 425.570 177.670 425.800 195.120 ;
        RECT 428.740 195.080 429.350 195.970 ;
        RECT 432.060 195.400 432.370 195.970 ;
        RECT 428.870 177.730 429.100 195.080 ;
        RECT 432.060 195.040 432.400 195.400 ;
        RECT 432.170 194.580 432.400 195.040 ;
        RECT 433.480 194.580 435.040 196.940 ;
        RECT 432.150 194.220 435.040 194.580 ;
        RECT 432.170 177.750 432.400 194.220 ;
        RECT 412.230 176.630 412.540 177.450 ;
        RECT 419.030 177.150 419.200 177.590 ;
        RECT 422.320 177.490 422.490 177.670 ;
        RECT 422.220 176.630 422.530 177.490 ;
        RECT 425.610 177.150 425.780 177.670 ;
        RECT 428.900 177.450 429.070 177.730 ;
        RECT 428.780 176.630 429.090 177.450 ;
        RECT 432.190 177.150 432.360 177.750 ;
        RECT 390.980 175.500 391.350 176.330 ;
        RECT 395.600 176.310 395.910 176.330 ;
        RECT 405.670 176.320 412.590 176.630 ;
        RECT 422.220 176.320 429.140 176.630 ;
        RECT 405.730 176.300 412.590 176.320 ;
        RECT 422.280 176.300 429.140 176.320 ;
        RECT 407.610 175.470 407.980 176.300 ;
        RECT 412.230 176.280 412.540 176.300 ;
        RECT 424.160 175.470 424.530 176.300 ;
        RECT 428.780 176.280 429.090 176.300 ;
        RECT 433.480 176.210 435.040 194.220 ;
        RECT 296.910 163.600 297.080 164.300 ;
        RECT 296.790 163.510 297.200 163.600 ;
        RECT 296.750 162.580 297.230 163.510 ;
        RECT 275.650 162.130 297.900 162.580 ;
        RECT 275.710 162.100 297.900 162.130 ;
        RECT 286.280 161.990 286.690 162.100 ;
        RECT 280.910 158.690 281.250 158.770 ;
        RECT 291.530 158.690 291.870 158.850 ;
        RECT 270.060 158.640 291.870 158.690 ;
        RECT 269.700 158.420 291.870 158.640 ;
        RECT 269.700 158.240 291.910 158.420 ;
        RECT 269.700 158.190 291.150 158.240 ;
        RECT 270.060 156.990 270.870 158.190 ;
        RECT 270.390 156.790 270.730 156.990 ;
        RECT 275.750 156.830 275.920 157.380 ;
        RECT 280.910 157.120 281.250 158.190 ;
        RECT 280.910 156.860 281.280 157.120 ;
        RECT 286.330 156.860 286.500 157.380 ;
        RECT 270.390 155.760 270.630 156.790 ;
        RECT 270.390 151.910 270.620 155.760 ;
        RECT 270.390 150.290 270.630 151.910 ;
        RECT 270.390 146.440 270.620 150.290 ;
        RECT 270.390 144.820 270.630 146.440 ;
        RECT 270.390 140.970 270.620 144.820 ;
        RECT 270.390 139.350 270.630 140.970 ;
        RECT 270.390 135.530 270.620 139.350 ;
        RECT 270.390 129.510 270.870 135.530 ;
        RECT 275.730 135.020 275.960 156.830 ;
        RECT 280.990 135.130 281.220 156.860 ;
        RECT 275.750 134.460 275.920 135.020 ;
        RECT 275.650 133.410 276.060 134.460 ;
        RECT 281.040 133.880 281.210 135.130 ;
        RECT 286.330 135.050 286.560 156.860 ;
        RECT 291.490 156.840 291.910 158.240 ;
        RECT 291.590 135.270 291.820 156.840 ;
        RECT 296.750 156.820 297.230 162.100 ;
        RECT 286.330 134.320 286.500 135.050 ;
        RECT 286.280 133.410 286.690 134.320 ;
        RECT 291.620 133.880 291.790 135.270 ;
        RECT 296.870 135.130 297.100 156.820 ;
        RECT 297.930 140.670 300.150 150.450 ;
        RECT 296.910 134.430 297.080 135.130 ;
        RECT 296.790 134.420 297.200 134.430 ;
        RECT 296.780 133.410 297.260 134.420 ;
        RECT 275.650 132.960 297.900 133.410 ;
        RECT 275.710 132.930 297.900 132.960 ;
        RECT 286.280 132.820 286.690 132.930 ;
        RECT 280.910 129.510 281.250 129.590 ;
        RECT 291.530 129.510 291.870 129.670 ;
        RECT 270.390 129.460 291.870 129.510 ;
        RECT 269.700 129.240 291.870 129.460 ;
        RECT 269.700 129.060 291.910 129.240 ;
        RECT 269.700 129.010 291.150 129.060 ;
        RECT 270.390 128.840 270.870 129.010 ;
        RECT 270.390 127.610 270.730 128.840 ;
        RECT 275.750 127.650 275.920 128.200 ;
        RECT 280.910 127.940 281.250 129.010 ;
        RECT 280.910 127.680 281.280 127.940 ;
        RECT 286.330 127.680 286.500 128.200 ;
        RECT 270.390 126.580 270.630 127.610 ;
        RECT 270.390 122.730 270.620 126.580 ;
        RECT 270.390 121.110 270.630 122.730 ;
        RECT 270.390 117.260 270.620 121.110 ;
        RECT 270.390 115.640 270.630 117.260 ;
        RECT 270.390 111.790 270.620 115.640 ;
        RECT 270.390 110.170 270.630 111.790 ;
        RECT 270.390 106.320 270.620 110.170 ;
        RECT 270.390 105.950 270.630 106.320 ;
        RECT 270.460 105.350 270.630 105.950 ;
        RECT 275.730 105.840 275.960 127.650 ;
        RECT 280.990 105.950 281.220 127.680 ;
        RECT 270.120 100.190 270.750 105.350 ;
        RECT 275.750 105.280 275.920 105.840 ;
        RECT 275.650 104.230 276.060 105.280 ;
        RECT 281.040 104.700 281.210 105.950 ;
        RECT 286.330 105.870 286.560 127.680 ;
        RECT 291.490 127.660 291.910 129.060 ;
        RECT 296.780 127.730 297.260 132.930 ;
        RECT 337.730 130.800 341.560 131.740 ;
        RECT 331.630 129.320 331.970 129.390 ;
        RECT 339.300 129.320 340.390 130.800 ;
        RECT 469.740 130.670 472.390 131.580 ;
        RECT 310.490 129.230 310.830 129.280 ;
        RECT 321.010 129.230 321.350 129.310 ;
        RECT 331.530 129.230 344.620 129.320 ;
        RECT 310.490 129.220 344.620 129.230 ;
        RECT 353.320 129.220 353.660 129.300 ;
        RECT 363.940 129.220 364.280 129.380 ;
        RECT 310.490 129.180 364.280 129.220 ;
        RECT 309.800 129.140 364.280 129.180 ;
        RECT 369.260 129.140 369.630 129.170 ;
        RECT 463.580 129.140 463.920 129.210 ;
        RECT 470.710 129.140 471.850 130.670 ;
        RECT 495.890 129.190 496.230 129.200 ;
        RECT 309.800 128.780 369.630 129.140 ;
        RECT 442.440 129.050 442.780 129.100 ;
        RECT 452.960 129.050 453.300 129.130 ;
        RECT 463.480 129.050 476.570 129.140 ;
        RECT 495.690 129.130 501.670 129.190 ;
        RECT 442.440 129.040 476.570 129.050 ;
        RECT 485.270 129.040 485.610 129.120 ;
        RECT 495.690 129.040 501.780 129.130 ;
        RECT 442.440 129.000 501.780 129.040 ;
        RECT 309.800 128.730 331.250 128.780 ;
        RECT 331.530 128.770 369.630 128.780 ;
        RECT 291.590 106.090 291.820 127.660 ;
        RECT 286.330 105.140 286.500 105.870 ;
        RECT 286.280 104.230 286.690 105.140 ;
        RECT 291.620 104.700 291.790 106.090 ;
        RECT 296.870 105.950 297.100 127.730 ;
        RECT 310.490 127.330 310.830 128.730 ;
        RECT 315.850 127.370 316.020 127.920 ;
        RECT 321.010 127.660 321.350 128.730 ;
        RECT 331.530 128.720 363.560 128.770 ;
        RECT 331.530 128.550 344.620 128.720 ;
        RECT 321.010 127.400 321.380 127.660 ;
        RECT 326.430 127.400 326.600 127.920 ;
        RECT 310.490 126.300 310.730 127.330 ;
        RECT 297.860 112.090 299.670 122.570 ;
        RECT 310.490 122.450 310.720 126.300 ;
        RECT 310.490 120.830 310.730 122.450 ;
        RECT 307.290 112.570 308.040 120.800 ;
        RECT 310.490 116.980 310.720 120.830 ;
        RECT 310.490 115.360 310.730 116.980 ;
        RECT 310.490 111.510 310.720 115.360 ;
        RECT 310.490 109.890 310.730 111.510 ;
        RECT 310.490 106.040 310.720 109.890 ;
        RECT 296.910 105.250 297.080 105.950 ;
        RECT 310.490 105.670 310.730 106.040 ;
        RECT 296.790 105.070 297.200 105.250 ;
        RECT 296.790 104.230 297.300 105.070 ;
        RECT 310.560 104.420 310.730 105.670 ;
        RECT 315.830 105.560 316.060 127.370 ;
        RECT 321.090 105.670 321.320 127.400 ;
        RECT 315.850 105.000 316.020 105.560 ;
        RECT 275.650 103.780 297.900 104.230 ;
        RECT 275.710 103.750 297.900 103.780 ;
        RECT 315.750 103.950 316.160 105.000 ;
        RECT 321.140 104.420 321.310 105.670 ;
        RECT 326.430 105.590 326.660 127.400 ;
        RECT 331.590 127.380 332.010 128.550 ;
        RECT 339.300 128.510 340.390 128.550 ;
        RECT 337.010 127.480 337.180 127.920 ;
        RECT 331.690 105.810 331.920 127.380 ;
        RECT 326.430 104.860 326.600 105.590 ;
        RECT 326.380 103.950 326.790 104.860 ;
        RECT 331.720 104.420 331.890 105.810 ;
        RECT 336.970 105.670 337.200 127.480 ;
        RECT 342.800 127.320 343.140 128.550 ;
        RECT 348.160 127.360 348.330 127.910 ;
        RECT 353.320 127.650 353.660 128.720 ;
        RECT 363.900 128.630 369.630 128.770 ;
        RECT 353.320 127.390 353.690 127.650 ;
        RECT 358.740 127.390 358.910 127.910 ;
        RECT 337.010 104.970 337.180 105.670 ;
        RECT 336.890 103.950 337.300 104.970 ;
        RECT 286.280 103.640 286.690 103.750 ;
        RECT 280.910 100.190 281.250 100.270 ;
        RECT 291.530 100.190 291.870 100.350 ;
        RECT 270.120 100.140 291.870 100.190 ;
        RECT 269.700 99.920 291.870 100.140 ;
        RECT 269.700 99.740 291.910 99.920 ;
        RECT 269.700 99.690 291.150 99.740 ;
        RECT 270.120 98.430 270.750 99.690 ;
        RECT 270.390 98.290 270.730 98.430 ;
        RECT 275.750 98.330 275.920 98.880 ;
        RECT 280.910 98.620 281.250 99.690 ;
        RECT 280.910 98.360 281.280 98.620 ;
        RECT 286.330 98.360 286.500 98.880 ;
        RECT 270.390 97.260 270.630 98.290 ;
        RECT 270.390 93.410 270.620 97.260 ;
        RECT 270.390 91.790 270.630 93.410 ;
        RECT 270.390 87.940 270.620 91.790 ;
        RECT 270.390 86.320 270.630 87.940 ;
        RECT 270.390 82.470 270.620 86.320 ;
        RECT 270.390 80.850 270.630 82.470 ;
        RECT 270.390 77.000 270.620 80.850 ;
        RECT 270.390 76.800 270.630 77.000 ;
        RECT 270.190 70.910 270.820 76.800 ;
        RECT 275.730 76.520 275.960 98.330 ;
        RECT 280.990 76.630 281.220 98.360 ;
        RECT 275.750 75.960 275.920 76.520 ;
        RECT 275.650 74.910 276.060 75.960 ;
        RECT 281.040 75.380 281.210 76.630 ;
        RECT 286.330 76.550 286.560 98.360 ;
        RECT 291.490 98.340 291.910 99.740 ;
        RECT 296.820 98.380 297.300 103.750 ;
        RECT 315.750 103.500 338.000 103.950 ;
        RECT 315.810 103.470 338.000 103.500 ;
        RECT 326.380 103.360 326.790 103.470 ;
        RECT 310.520 100.040 310.860 100.090 ;
        RECT 321.040 100.040 321.380 100.120 ;
        RECT 331.660 100.040 332.000 100.200 ;
        RECT 310.520 99.990 332.000 100.040 ;
        RECT 309.830 99.770 332.000 99.990 ;
        RECT 309.830 99.590 332.040 99.770 ;
        RECT 309.830 99.540 331.280 99.590 ;
        RECT 291.590 76.770 291.820 98.340 ;
        RECT 286.330 75.820 286.500 76.550 ;
        RECT 286.280 74.910 286.690 75.820 ;
        RECT 291.620 75.380 291.790 76.770 ;
        RECT 296.870 76.630 297.100 98.380 ;
        RECT 310.520 98.140 310.860 99.540 ;
        RECT 315.880 98.180 316.050 98.730 ;
        RECT 321.040 98.470 321.380 99.540 ;
        RECT 321.040 98.210 321.410 98.470 ;
        RECT 326.460 98.210 326.630 98.730 ;
        RECT 310.520 97.110 310.760 98.140 ;
        RECT 298.140 83.510 300.010 93.430 ;
        RECT 310.520 93.260 310.750 97.110 ;
        RECT 310.520 91.640 310.760 93.260 ;
        RECT 307.320 83.380 308.070 91.610 ;
        RECT 310.520 87.790 310.750 91.640 ;
        RECT 310.520 86.170 310.760 87.790 ;
        RECT 310.520 82.320 310.750 86.170 ;
        RECT 310.520 80.700 310.760 82.320 ;
        RECT 310.520 76.850 310.750 80.700 ;
        RECT 296.910 75.960 297.080 76.630 ;
        RECT 310.520 76.480 310.760 76.850 ;
        RECT 296.910 75.930 297.540 75.960 ;
        RECT 296.790 74.910 297.540 75.930 ;
        RECT 310.590 75.230 310.760 76.480 ;
        RECT 315.860 76.370 316.090 98.180 ;
        RECT 321.120 76.480 321.350 98.210 ;
        RECT 315.880 75.810 316.050 76.370 ;
        RECT 275.650 74.460 297.900 74.910 ;
        RECT 275.710 74.430 297.900 74.460 ;
        RECT 315.780 74.760 316.190 75.810 ;
        RECT 321.170 75.230 321.340 76.480 ;
        RECT 326.460 76.400 326.690 98.210 ;
        RECT 331.620 98.190 332.040 99.590 ;
        RECT 337.040 98.290 337.210 98.730 ;
        RECT 331.720 76.620 331.950 98.190 ;
        RECT 326.460 75.670 326.630 76.400 ;
        RECT 326.410 74.760 326.820 75.670 ;
        RECT 331.750 75.230 331.920 76.620 ;
        RECT 337.000 76.480 337.230 98.290 ;
        RECT 337.040 75.780 337.210 76.480 ;
        RECT 336.920 74.760 337.330 75.780 ;
        RECT 286.280 74.320 286.690 74.430 ;
        RECT 280.960 70.910 281.300 70.990 ;
        RECT 291.580 70.910 291.920 71.070 ;
        RECT 270.190 70.860 291.920 70.910 ;
        RECT 269.750 70.640 291.920 70.860 ;
        RECT 269.750 70.460 291.960 70.640 ;
        RECT 269.750 70.410 291.200 70.460 ;
        RECT 270.190 69.880 270.820 70.410 ;
        RECT 270.440 69.010 270.780 69.880 ;
        RECT 275.800 69.050 275.970 69.600 ;
        RECT 280.960 69.340 281.300 70.410 ;
        RECT 280.960 69.080 281.330 69.340 ;
        RECT 286.380 69.080 286.550 69.600 ;
        RECT 270.440 67.980 270.680 69.010 ;
        RECT 270.440 64.130 270.670 67.980 ;
        RECT 270.440 62.510 270.680 64.130 ;
        RECT 270.440 58.660 270.670 62.510 ;
        RECT 270.440 57.040 270.680 58.660 ;
        RECT 270.440 53.190 270.670 57.040 ;
        RECT 270.440 51.570 270.680 53.190 ;
        RECT 270.440 47.720 270.670 51.570 ;
        RECT 270.440 47.440 270.680 47.720 ;
        RECT 270.260 47.270 270.880 47.440 ;
        RECT 270.260 41.370 270.890 47.270 ;
        RECT 275.780 47.240 276.010 69.050 ;
        RECT 281.040 47.350 281.270 69.080 ;
        RECT 275.800 46.680 275.970 47.240 ;
        RECT 275.700 45.630 276.110 46.680 ;
        RECT 281.090 46.100 281.260 47.350 ;
        RECT 286.380 47.270 286.610 69.080 ;
        RECT 291.540 69.060 291.960 70.460 ;
        RECT 291.640 47.490 291.870 69.060 ;
        RECT 296.910 69.040 297.540 74.430 ;
        RECT 315.780 74.310 338.030 74.760 ;
        RECT 315.840 74.280 338.030 74.310 ;
        RECT 326.410 74.170 326.820 74.280 ;
        RECT 310.520 70.750 310.860 70.800 ;
        RECT 321.040 70.750 321.380 70.830 ;
        RECT 331.660 70.750 332.000 70.910 ;
        RECT 310.520 70.700 332.000 70.750 ;
        RECT 309.830 70.480 332.000 70.700 ;
        RECT 309.830 70.300 332.040 70.480 ;
        RECT 309.830 70.250 331.280 70.300 ;
        RECT 286.380 46.540 286.550 47.270 ;
        RECT 286.330 45.630 286.740 46.540 ;
        RECT 291.670 46.100 291.840 47.490 ;
        RECT 296.920 47.350 297.150 69.040 ;
        RECT 310.520 68.850 310.860 70.250 ;
        RECT 315.880 68.890 316.050 69.440 ;
        RECT 321.040 69.180 321.380 70.250 ;
        RECT 321.040 68.920 321.410 69.180 ;
        RECT 326.460 68.920 326.630 69.440 ;
        RECT 310.520 67.820 310.760 68.850 ;
        RECT 310.520 63.970 310.750 67.820 ;
        RECT 298.210 55.010 300.010 63.470 ;
        RECT 310.520 62.350 310.760 63.970 ;
        RECT 307.320 54.090 308.070 62.320 ;
        RECT 310.520 58.500 310.750 62.350 ;
        RECT 310.520 56.880 310.760 58.500 ;
        RECT 310.520 53.030 310.750 56.880 ;
        RECT 310.520 51.410 310.760 53.030 ;
        RECT 310.520 47.560 310.750 51.410 ;
        RECT 296.960 46.650 297.130 47.350 ;
        RECT 310.520 47.190 310.760 47.560 ;
        RECT 296.840 46.080 297.250 46.650 ;
        RECT 296.840 45.630 297.470 46.080 ;
        RECT 310.590 45.940 310.760 47.190 ;
        RECT 315.860 47.080 316.090 68.890 ;
        RECT 321.120 47.190 321.350 68.920 ;
        RECT 315.880 46.520 316.050 47.080 ;
        RECT 275.700 45.180 297.950 45.630 ;
        RECT 275.760 45.150 297.950 45.180 ;
        RECT 315.780 45.470 316.190 46.520 ;
        RECT 321.170 45.940 321.340 47.190 ;
        RECT 326.460 47.110 326.690 68.920 ;
        RECT 331.620 68.900 332.040 70.300 ;
        RECT 337.040 69.000 337.210 69.440 ;
        RECT 331.720 47.330 331.950 68.900 ;
        RECT 326.460 46.380 326.630 47.110 ;
        RECT 326.410 45.470 326.820 46.380 ;
        RECT 331.750 45.940 331.920 47.330 ;
        RECT 337.000 47.190 337.230 69.000 ;
        RECT 337.040 46.490 337.210 47.190 ;
        RECT 336.920 45.470 337.330 46.490 ;
        RECT 286.330 45.040 286.740 45.150 ;
        RECT 281.050 41.370 281.390 41.450 ;
        RECT 291.670 41.370 292.010 41.530 ;
        RECT 270.260 41.320 292.010 41.370 ;
        RECT 269.840 41.100 292.010 41.320 ;
        RECT 269.840 40.920 292.050 41.100 ;
        RECT 269.840 40.870 291.290 40.920 ;
        RECT 270.260 40.350 270.890 40.870 ;
        RECT 270.530 39.470 270.870 40.350 ;
        RECT 275.890 39.510 276.060 40.060 ;
        RECT 281.050 39.800 281.390 40.870 ;
        RECT 281.050 39.540 281.420 39.800 ;
        RECT 286.470 39.540 286.640 40.060 ;
        RECT 270.530 38.440 270.770 39.470 ;
        RECT 270.530 34.590 270.760 38.440 ;
        RECT 270.530 32.970 270.770 34.590 ;
        RECT 270.530 29.120 270.760 32.970 ;
        RECT 270.530 27.500 270.770 29.120 ;
        RECT 267.330 24.710 268.080 26.880 ;
        RECT 270.530 23.650 270.760 27.500 ;
        RECT 270.530 22.030 270.770 23.650 ;
        RECT 270.530 18.180 270.760 22.030 ;
        RECT 270.530 17.810 270.770 18.180 ;
        RECT 264.480 17.040 264.650 17.740 ;
        RECT 264.360 16.240 264.770 17.040 ;
        RECT 270.600 16.560 270.770 17.810 ;
        RECT 275.870 17.700 276.100 39.510 ;
        RECT 281.130 17.810 281.360 39.540 ;
        RECT 275.890 17.140 276.060 17.700 ;
        RECT 275.790 16.240 276.200 17.140 ;
        RECT 281.180 16.560 281.350 17.810 ;
        RECT 286.470 17.730 286.700 39.540 ;
        RECT 291.630 39.520 292.050 40.920 ;
        RECT 291.730 17.950 291.960 39.520 ;
        RECT 296.840 39.160 297.470 45.150 ;
        RECT 315.780 45.020 338.030 45.470 ;
        RECT 315.840 44.990 338.030 45.020 ;
        RECT 326.410 44.880 326.820 44.990 ;
        RECT 310.520 41.460 310.860 41.510 ;
        RECT 321.040 41.460 321.380 41.540 ;
        RECT 331.660 41.460 332.000 41.620 ;
        RECT 310.520 41.410 332.000 41.460 ;
        RECT 309.830 41.190 332.000 41.410 ;
        RECT 309.830 41.010 332.040 41.190 ;
        RECT 309.830 40.960 331.280 41.010 ;
        RECT 310.520 39.560 310.860 40.960 ;
        RECT 315.880 39.600 316.050 40.150 ;
        RECT 321.040 39.890 321.380 40.960 ;
        RECT 321.040 39.630 321.410 39.890 ;
        RECT 326.460 39.630 326.630 40.150 ;
        RECT 286.470 17.000 286.640 17.730 ;
        RECT 231.420 16.090 283.600 16.240 ;
        RECT 286.420 16.090 286.830 17.000 ;
        RECT 291.760 16.560 291.930 17.950 ;
        RECT 297.010 17.810 297.240 39.160 ;
        RECT 310.520 38.530 310.760 39.560 ;
        RECT 310.520 34.680 310.750 38.530 ;
        RECT 298.000 29.680 299.740 34.060 ;
        RECT 310.520 33.060 310.760 34.680 ;
        RECT 298.000 25.870 300.800 29.680 ;
        RECT 297.050 17.110 297.220 17.810 ;
        RECT 296.930 16.090 297.340 17.110 ;
        RECT 231.420 15.910 298.040 16.090 ;
        RECT 210.280 15.610 298.040 15.910 ;
        RECT 210.280 15.460 283.600 15.610 ;
        RECT 286.420 15.500 286.830 15.610 ;
        RECT 210.340 15.430 283.600 15.460 ;
        RECT 220.910 15.320 221.320 15.430 ;
        RECT 231.770 15.210 283.600 15.430 ;
        RECT 298.590 -0.920 300.800 25.870 ;
        RECT 307.320 24.800 308.070 33.030 ;
        RECT 310.520 29.210 310.750 33.060 ;
        RECT 310.520 27.590 310.760 29.210 ;
        RECT 310.520 23.740 310.750 27.590 ;
        RECT 310.520 22.120 310.760 23.740 ;
        RECT 310.520 18.270 310.750 22.120 ;
        RECT 310.520 17.900 310.760 18.270 ;
        RECT 310.590 16.650 310.760 17.900 ;
        RECT 315.860 17.790 316.090 39.600 ;
        RECT 321.120 17.900 321.350 39.630 ;
        RECT 315.880 17.230 316.050 17.790 ;
        RECT 315.780 16.180 316.190 17.230 ;
        RECT 321.170 16.650 321.340 17.900 ;
        RECT 326.460 17.820 326.690 39.630 ;
        RECT 331.620 39.610 332.040 41.010 ;
        RECT 337.040 39.710 337.210 40.150 ;
        RECT 331.720 18.040 331.950 39.610 ;
        RECT 326.460 17.090 326.630 17.820 ;
        RECT 326.410 16.180 326.820 17.090 ;
        RECT 331.750 16.650 331.920 18.040 ;
        RECT 337.000 17.900 337.230 39.710 ;
        RECT 338.460 23.960 341.620 126.810 ;
        RECT 342.800 126.290 343.040 127.320 ;
        RECT 342.800 122.440 343.030 126.290 ;
        RECT 342.800 120.820 343.040 122.440 ;
        RECT 342.800 116.970 343.030 120.820 ;
        RECT 342.800 115.350 343.040 116.970 ;
        RECT 342.800 111.500 343.030 115.350 ;
        RECT 342.800 109.880 343.040 111.500 ;
        RECT 342.800 106.030 343.030 109.880 ;
        RECT 342.800 105.660 343.040 106.030 ;
        RECT 342.870 104.410 343.040 105.660 ;
        RECT 348.140 105.550 348.370 127.360 ;
        RECT 353.400 105.660 353.630 127.390 ;
        RECT 348.160 104.990 348.330 105.550 ;
        RECT 348.060 103.940 348.470 104.990 ;
        RECT 353.450 104.410 353.620 105.660 ;
        RECT 358.740 105.580 358.970 127.390 ;
        RECT 363.900 127.370 364.320 128.630 ;
        RECT 364.000 105.800 364.230 127.370 ;
        RECT 369.260 127.260 369.630 128.630 ;
        RECT 441.750 128.600 501.780 129.000 ;
        RECT 441.750 128.550 463.200 128.600 ;
        RECT 463.480 128.590 501.780 128.600 ;
        RECT 358.740 104.850 358.910 105.580 ;
        RECT 358.690 103.940 359.100 104.850 ;
        RECT 364.030 104.410 364.200 105.800 ;
        RECT 369.280 105.660 369.510 127.260 ;
        RECT 381.630 127.230 381.800 127.780 ;
        RECT 392.210 127.260 392.380 127.780 ;
        RECT 402.790 127.340 402.960 127.780 ;
        RECT 369.320 104.960 369.490 105.660 ;
        RECT 369.200 103.940 369.610 104.960 ;
        RECT 348.060 103.490 370.310 103.940 ;
        RECT 348.120 103.460 370.310 103.490 ;
        RECT 358.690 103.350 359.100 103.460 ;
        RECT 342.840 100.100 343.180 100.150 ;
        RECT 353.360 100.100 353.700 100.180 ;
        RECT 363.980 100.100 364.320 100.260 ;
        RECT 342.840 100.050 364.320 100.100 ;
        RECT 342.150 99.830 364.320 100.050 ;
        RECT 342.150 99.650 364.360 99.830 ;
        RECT 342.150 99.600 363.600 99.650 ;
        RECT 342.840 98.200 343.180 99.600 ;
        RECT 348.200 98.240 348.370 98.790 ;
        RECT 353.360 98.530 353.700 99.600 ;
        RECT 353.360 98.270 353.730 98.530 ;
        RECT 358.780 98.270 358.950 98.790 ;
        RECT 342.840 97.170 343.080 98.200 ;
        RECT 342.840 93.320 343.070 97.170 ;
        RECT 342.840 91.700 343.080 93.320 ;
        RECT 342.840 87.850 343.070 91.700 ;
        RECT 342.840 86.230 343.080 87.850 ;
        RECT 342.840 82.380 343.070 86.230 ;
        RECT 342.840 80.760 343.080 82.380 ;
        RECT 342.840 76.910 343.070 80.760 ;
        RECT 342.840 76.540 343.080 76.910 ;
        RECT 342.910 75.290 343.080 76.540 ;
        RECT 348.180 76.430 348.410 98.240 ;
        RECT 353.440 76.540 353.670 98.270 ;
        RECT 348.200 75.870 348.370 76.430 ;
        RECT 348.100 74.820 348.510 75.870 ;
        RECT 353.490 75.290 353.660 76.540 ;
        RECT 358.780 76.460 359.010 98.270 ;
        RECT 363.940 98.250 364.360 99.650 ;
        RECT 369.360 98.350 369.530 98.790 ;
        RECT 364.040 76.680 364.270 98.250 ;
        RECT 358.780 75.730 358.950 76.460 ;
        RECT 358.730 74.820 359.140 75.730 ;
        RECT 364.070 75.290 364.240 76.680 ;
        RECT 369.320 76.540 369.550 98.350 ;
        RECT 369.360 75.840 369.530 76.540 ;
        RECT 369.240 74.820 369.650 75.840 ;
        RECT 348.100 74.370 370.350 74.820 ;
        RECT 348.160 74.340 370.350 74.370 ;
        RECT 358.730 74.230 359.140 74.340 ;
        RECT 342.860 70.740 343.200 70.790 ;
        RECT 353.380 70.740 353.720 70.820 ;
        RECT 364.000 70.740 364.340 70.900 ;
        RECT 342.860 70.690 364.340 70.740 ;
        RECT 342.170 70.470 364.340 70.690 ;
        RECT 342.170 70.290 364.380 70.470 ;
        RECT 342.170 70.240 363.620 70.290 ;
        RECT 342.860 68.840 343.200 70.240 ;
        RECT 348.220 68.880 348.390 69.430 ;
        RECT 353.380 69.170 353.720 70.240 ;
        RECT 353.380 68.910 353.750 69.170 ;
        RECT 358.800 68.910 358.970 69.430 ;
        RECT 342.860 67.810 343.100 68.840 ;
        RECT 342.860 63.960 343.090 67.810 ;
        RECT 342.860 62.340 343.100 63.960 ;
        RECT 342.860 58.490 343.090 62.340 ;
        RECT 342.860 56.870 343.100 58.490 ;
        RECT 342.860 53.020 343.090 56.870 ;
        RECT 342.860 51.400 343.100 53.020 ;
        RECT 342.860 47.550 343.090 51.400 ;
        RECT 342.860 47.180 343.100 47.550 ;
        RECT 342.930 45.930 343.100 47.180 ;
        RECT 348.200 47.070 348.430 68.880 ;
        RECT 353.460 47.180 353.690 68.910 ;
        RECT 348.220 46.510 348.390 47.070 ;
        RECT 348.120 45.460 348.530 46.510 ;
        RECT 353.510 45.930 353.680 47.180 ;
        RECT 358.800 47.100 359.030 68.910 ;
        RECT 363.960 68.890 364.380 70.290 ;
        RECT 369.380 68.990 369.550 69.430 ;
        RECT 364.060 47.320 364.290 68.890 ;
        RECT 358.800 46.370 358.970 47.100 ;
        RECT 358.750 45.460 359.160 46.370 ;
        RECT 364.090 45.930 364.260 47.320 ;
        RECT 369.340 47.180 369.570 68.990 ;
        RECT 369.380 46.480 369.550 47.180 ;
        RECT 369.260 45.460 369.670 46.480 ;
        RECT 348.120 45.010 370.370 45.460 ;
        RECT 348.180 44.980 370.370 45.010 ;
        RECT 358.750 44.870 359.160 44.980 ;
        RECT 342.880 41.450 343.220 41.500 ;
        RECT 353.400 41.450 353.740 41.530 ;
        RECT 364.020 41.450 364.360 41.610 ;
        RECT 342.880 41.400 364.360 41.450 ;
        RECT 342.190 41.180 364.360 41.400 ;
        RECT 342.190 41.000 364.400 41.180 ;
        RECT 342.190 40.950 363.640 41.000 ;
        RECT 342.880 39.550 343.220 40.950 ;
        RECT 348.240 39.590 348.410 40.140 ;
        RECT 353.400 39.880 353.740 40.950 ;
        RECT 353.400 39.620 353.770 39.880 ;
        RECT 358.820 39.620 358.990 40.140 ;
        RECT 342.880 38.520 343.120 39.550 ;
        RECT 342.880 34.670 343.110 38.520 ;
        RECT 342.880 33.050 343.120 34.670 ;
        RECT 342.880 29.200 343.110 33.050 ;
        RECT 342.880 27.580 343.120 29.200 ;
        RECT 337.040 17.200 337.210 17.900 ;
        RECT 336.920 16.210 337.330 17.200 ;
        RECT 338.530 16.210 341.290 23.960 ;
        RECT 342.880 23.730 343.110 27.580 ;
        RECT 342.880 22.110 343.120 23.730 ;
        RECT 342.880 18.260 343.110 22.110 ;
        RECT 342.880 17.890 343.120 18.260 ;
        RECT 342.950 16.640 343.120 17.890 ;
        RECT 348.220 17.780 348.450 39.590 ;
        RECT 353.480 17.890 353.710 39.620 ;
        RECT 348.240 17.220 348.410 17.780 ;
        RECT 348.140 16.210 348.550 17.220 ;
        RECT 353.530 16.640 353.700 17.890 ;
        RECT 358.820 17.810 359.050 39.620 ;
        RECT 363.980 39.600 364.400 41.000 ;
        RECT 369.400 39.700 369.570 40.140 ;
        RECT 364.080 18.030 364.310 39.600 ;
        RECT 358.820 17.080 358.990 17.810 ;
        RECT 336.920 16.180 348.700 16.210 ;
        RECT 315.780 16.170 348.700 16.180 ;
        RECT 358.770 16.170 359.180 17.080 ;
        RECT 364.110 16.640 364.280 18.030 ;
        RECT 369.360 17.890 369.590 39.700 ;
        RECT 369.400 17.190 369.570 17.890 ;
        RECT 369.280 16.170 369.690 17.190 ;
        RECT 371.400 17.060 375.330 124.410 ;
        RECT 381.610 105.420 381.840 127.230 ;
        RECT 392.210 105.450 392.440 127.260 ;
        RECT 402.750 105.530 402.980 127.340 ;
        RECT 413.940 127.220 414.110 127.770 ;
        RECT 424.520 127.250 424.690 127.770 ;
        RECT 435.100 127.330 435.270 127.770 ;
        RECT 381.630 104.860 381.800 105.420 ;
        RECT 381.530 103.810 381.940 104.860 ;
        RECT 392.210 104.720 392.380 105.450 ;
        RECT 402.790 104.830 402.960 105.530 ;
        RECT 392.160 103.810 392.570 104.720 ;
        RECT 402.670 103.810 403.080 104.830 ;
        RECT 403.590 103.850 407.520 124.750 ;
        RECT 413.920 105.410 414.150 127.220 ;
        RECT 424.520 105.440 424.750 127.250 ;
        RECT 435.060 105.520 435.290 127.330 ;
        RECT 442.440 127.150 442.780 128.550 ;
        RECT 447.800 127.190 447.970 127.740 ;
        RECT 452.960 127.480 453.300 128.550 ;
        RECT 463.480 128.540 495.510 128.590 ;
        RECT 463.480 128.370 476.570 128.540 ;
        RECT 452.960 127.220 453.330 127.480 ;
        RECT 458.380 127.220 458.550 127.740 ;
        RECT 442.440 126.120 442.680 127.150 ;
        RECT 438.100 125.520 441.120 125.530 ;
        RECT 413.940 104.850 414.110 105.410 ;
        RECT 381.530 103.360 403.310 103.810 ;
        RECT 381.590 103.330 403.310 103.360 ;
        RECT 392.160 103.220 392.570 103.330 ;
        RECT 403.600 103.180 407.520 103.850 ;
        RECT 413.840 103.800 414.250 104.850 ;
        RECT 424.520 104.710 424.690 105.440 ;
        RECT 435.100 104.820 435.270 105.520 ;
        RECT 424.470 103.800 424.880 104.710 ;
        RECT 434.980 103.800 435.390 104.820 ;
        RECT 413.840 103.350 436.090 103.800 ;
        RECT 413.900 103.320 436.090 103.350 ;
        RECT 424.470 103.210 424.880 103.320 ;
        RECT 381.660 98.040 381.830 98.590 ;
        RECT 392.240 98.070 392.410 98.590 ;
        RECT 402.820 98.150 402.990 98.590 ;
        RECT 381.640 76.230 381.870 98.040 ;
        RECT 392.240 76.260 392.470 98.070 ;
        RECT 402.780 76.340 403.010 98.150 ;
        RECT 381.660 75.670 381.830 76.230 ;
        RECT 381.560 74.620 381.970 75.670 ;
        RECT 392.240 75.530 392.410 76.260 ;
        RECT 402.820 75.640 402.990 76.340 ;
        RECT 392.190 74.620 392.600 75.530 ;
        RECT 402.700 74.620 403.110 75.640 ;
        RECT 403.590 74.620 407.520 103.180 ;
        RECT 413.980 98.100 414.150 98.650 ;
        RECT 424.560 98.130 424.730 98.650 ;
        RECT 435.140 98.210 435.310 98.650 ;
        RECT 413.960 76.290 414.190 98.100 ;
        RECT 424.560 76.320 424.790 98.130 ;
        RECT 435.100 76.400 435.330 98.210 ;
        RECT 413.980 75.730 414.150 76.290 ;
        RECT 381.560 74.170 403.280 74.620 ;
        RECT 381.620 74.140 403.280 74.170 ;
        RECT 403.570 74.140 407.520 74.620 ;
        RECT 413.880 74.680 414.290 75.730 ;
        RECT 424.560 75.590 424.730 76.320 ;
        RECT 435.140 75.700 435.310 76.400 ;
        RECT 424.510 74.680 424.920 75.590 ;
        RECT 435.020 74.680 435.430 75.700 ;
        RECT 413.880 74.230 436.130 74.680 ;
        RECT 413.940 74.200 436.130 74.230 ;
        RECT 392.190 74.030 392.600 74.140 ;
        RECT 381.660 68.750 381.830 69.300 ;
        RECT 392.240 68.780 392.410 69.300 ;
        RECT 402.820 68.860 402.990 69.300 ;
        RECT 381.640 46.940 381.870 68.750 ;
        RECT 392.240 46.970 392.470 68.780 ;
        RECT 402.780 47.050 403.010 68.860 ;
        RECT 381.660 46.380 381.830 46.940 ;
        RECT 381.560 45.330 381.970 46.380 ;
        RECT 392.240 46.240 392.410 46.970 ;
        RECT 402.820 46.350 402.990 47.050 ;
        RECT 392.190 45.330 392.600 46.240 ;
        RECT 402.700 45.330 403.110 46.350 ;
        RECT 403.590 45.440 407.520 74.140 ;
        RECT 424.510 74.090 424.920 74.200 ;
        RECT 414.000 68.740 414.170 69.290 ;
        RECT 424.580 68.770 424.750 69.290 ;
        RECT 435.160 68.850 435.330 69.290 ;
        RECT 413.980 46.930 414.210 68.740 ;
        RECT 424.580 46.960 424.810 68.770 ;
        RECT 435.120 47.040 435.350 68.850 ;
        RECT 414.000 46.370 414.170 46.930 ;
        RECT 381.560 44.880 403.310 45.330 ;
        RECT 381.620 44.850 403.310 44.880 ;
        RECT 392.190 44.740 392.600 44.850 ;
        RECT 403.600 44.770 407.520 45.440 ;
        RECT 413.900 45.320 414.310 46.370 ;
        RECT 424.580 46.230 424.750 46.960 ;
        RECT 435.160 46.340 435.330 47.040 ;
        RECT 424.530 45.320 424.940 46.230 ;
        RECT 435.040 45.320 435.450 46.340 ;
        RECT 413.900 44.870 436.150 45.320 ;
        RECT 413.960 44.840 436.150 44.870 ;
        RECT 381.660 39.460 381.830 40.010 ;
        RECT 392.240 39.490 392.410 40.010 ;
        RECT 402.820 39.570 402.990 40.010 ;
        RECT 381.640 17.650 381.870 39.460 ;
        RECT 392.240 17.680 392.470 39.490 ;
        RECT 402.780 17.760 403.010 39.570 ;
        RECT 381.660 17.090 381.830 17.650 ;
        RECT 315.780 15.730 370.390 16.170 ;
        RECT 315.840 15.700 370.390 15.730 ;
        RECT 326.410 15.590 326.820 15.700 ;
        RECT 337.090 15.690 370.390 15.700 ;
        RECT 337.090 15.660 348.700 15.690 ;
        RECT 338.530 4.200 341.290 15.660 ;
        RECT 358.770 15.580 359.180 15.690 ;
        RECT 199.180 -6.230 207.790 -2.480 ;
        RECT 297.600 -3.410 302.970 -0.920 ;
        RECT 335.400 -0.960 346.270 4.200 ;
        RECT 372.060 4.020 374.820 17.060 ;
        RECT 381.560 16.040 381.970 17.090 ;
        RECT 392.240 16.950 392.410 17.680 ;
        RECT 402.820 17.060 402.990 17.760 ;
        RECT 403.590 17.400 407.520 44.770 ;
        RECT 424.530 44.730 424.940 44.840 ;
        RECT 414.020 39.450 414.190 40.000 ;
        RECT 424.600 39.480 424.770 40.000 ;
        RECT 435.180 39.560 435.350 40.000 ;
        RECT 414.000 17.640 414.230 39.450 ;
        RECT 424.600 17.670 424.830 39.480 ;
        RECT 435.140 17.750 435.370 39.560 ;
        RECT 436.820 18.190 441.120 125.520 ;
        RECT 442.440 122.270 442.670 126.120 ;
        RECT 442.440 120.650 442.680 122.270 ;
        RECT 442.440 116.800 442.670 120.650 ;
        RECT 442.440 115.180 442.680 116.800 ;
        RECT 442.440 111.330 442.670 115.180 ;
        RECT 442.440 109.710 442.680 111.330 ;
        RECT 442.440 105.860 442.670 109.710 ;
        RECT 442.440 105.490 442.680 105.860 ;
        RECT 442.510 104.240 442.680 105.490 ;
        RECT 447.780 105.380 448.010 127.190 ;
        RECT 453.040 105.490 453.270 127.220 ;
        RECT 447.800 104.820 447.970 105.380 ;
        RECT 447.700 103.770 448.110 104.820 ;
        RECT 453.090 104.240 453.260 105.490 ;
        RECT 458.380 105.410 458.610 127.220 ;
        RECT 463.540 127.200 463.960 128.370 ;
        RECT 468.960 127.300 469.130 127.740 ;
        RECT 463.640 105.630 463.870 127.200 ;
        RECT 458.380 104.680 458.550 105.410 ;
        RECT 458.330 103.770 458.740 104.680 ;
        RECT 463.670 104.240 463.840 105.630 ;
        RECT 468.920 105.490 469.150 127.300 ;
        RECT 474.750 127.140 475.090 128.370 ;
        RECT 480.110 127.180 480.280 127.730 ;
        RECT 485.270 127.470 485.610 128.540 ;
        RECT 495.690 128.390 501.780 128.590 ;
        RECT 485.270 127.210 485.640 127.470 ;
        RECT 490.690 127.210 490.860 127.730 ;
        RECT 474.750 126.110 474.990 127.140 ;
        RECT 468.960 104.790 469.130 105.490 ;
        RECT 468.840 103.770 469.250 104.790 ;
        RECT 447.700 103.320 469.950 103.770 ;
        RECT 447.760 103.290 469.950 103.320 ;
        RECT 458.330 103.180 458.740 103.290 ;
        RECT 442.470 99.860 442.810 99.910 ;
        RECT 452.990 99.860 453.330 99.940 ;
        RECT 463.610 99.860 463.950 100.020 ;
        RECT 442.470 99.810 463.950 99.860 ;
        RECT 441.780 99.590 463.950 99.810 ;
        RECT 441.780 99.410 463.990 99.590 ;
        RECT 441.780 99.360 463.230 99.410 ;
        RECT 442.470 97.960 442.810 99.360 ;
        RECT 447.830 98.000 448.000 98.550 ;
        RECT 452.990 98.290 453.330 99.360 ;
        RECT 452.990 98.030 453.360 98.290 ;
        RECT 458.410 98.030 458.580 98.550 ;
        RECT 442.470 96.930 442.710 97.960 ;
        RECT 442.470 93.080 442.700 96.930 ;
        RECT 442.470 91.460 442.710 93.080 ;
        RECT 442.470 87.610 442.700 91.460 ;
        RECT 442.470 85.990 442.710 87.610 ;
        RECT 442.470 82.140 442.700 85.990 ;
        RECT 442.470 80.520 442.710 82.140 ;
        RECT 442.470 76.670 442.700 80.520 ;
        RECT 442.470 76.300 442.710 76.670 ;
        RECT 442.540 75.050 442.710 76.300 ;
        RECT 447.810 76.190 448.040 98.000 ;
        RECT 453.070 76.300 453.300 98.030 ;
        RECT 447.830 75.630 448.000 76.190 ;
        RECT 447.730 74.580 448.140 75.630 ;
        RECT 453.120 75.050 453.290 76.300 ;
        RECT 458.410 76.220 458.640 98.030 ;
        RECT 463.570 98.010 463.990 99.410 ;
        RECT 468.990 98.110 469.160 98.550 ;
        RECT 463.670 76.440 463.900 98.010 ;
        RECT 458.410 75.490 458.580 76.220 ;
        RECT 458.360 74.580 458.770 75.490 ;
        RECT 463.700 75.050 463.870 76.440 ;
        RECT 468.950 76.300 469.180 98.110 ;
        RECT 468.990 75.600 469.160 76.300 ;
        RECT 468.870 74.580 469.280 75.600 ;
        RECT 447.730 74.130 469.980 74.580 ;
        RECT 447.790 74.100 469.980 74.130 ;
        RECT 458.360 73.990 458.770 74.100 ;
        RECT 442.470 70.570 442.810 70.620 ;
        RECT 452.990 70.570 453.330 70.650 ;
        RECT 463.610 70.570 463.950 70.730 ;
        RECT 442.470 70.520 463.950 70.570 ;
        RECT 441.780 70.300 463.950 70.520 ;
        RECT 441.780 70.120 463.990 70.300 ;
        RECT 441.780 70.070 463.230 70.120 ;
        RECT 442.470 68.670 442.810 70.070 ;
        RECT 447.830 68.710 448.000 69.260 ;
        RECT 452.990 69.000 453.330 70.070 ;
        RECT 452.990 68.740 453.360 69.000 ;
        RECT 458.410 68.740 458.580 69.260 ;
        RECT 442.470 67.640 442.710 68.670 ;
        RECT 442.470 63.790 442.700 67.640 ;
        RECT 442.470 62.170 442.710 63.790 ;
        RECT 442.470 58.320 442.700 62.170 ;
        RECT 442.470 56.700 442.710 58.320 ;
        RECT 442.470 52.850 442.700 56.700 ;
        RECT 442.470 51.230 442.710 52.850 ;
        RECT 442.470 47.380 442.700 51.230 ;
        RECT 442.470 47.010 442.710 47.380 ;
        RECT 442.540 45.760 442.710 47.010 ;
        RECT 447.810 46.900 448.040 68.710 ;
        RECT 453.070 47.010 453.300 68.740 ;
        RECT 447.830 46.340 448.000 46.900 ;
        RECT 447.730 45.290 448.140 46.340 ;
        RECT 453.120 45.760 453.290 47.010 ;
        RECT 458.410 46.930 458.640 68.740 ;
        RECT 463.570 68.720 463.990 70.120 ;
        RECT 468.990 68.820 469.160 69.260 ;
        RECT 463.670 47.150 463.900 68.720 ;
        RECT 458.410 46.200 458.580 46.930 ;
        RECT 458.360 45.290 458.770 46.200 ;
        RECT 463.700 45.760 463.870 47.150 ;
        RECT 468.950 47.010 469.180 68.820 ;
        RECT 468.990 46.310 469.160 47.010 ;
        RECT 468.870 45.290 469.280 46.310 ;
        RECT 447.730 44.840 469.980 45.290 ;
        RECT 447.790 44.810 469.980 44.840 ;
        RECT 458.360 44.700 458.770 44.810 ;
        RECT 442.470 41.280 442.810 41.330 ;
        RECT 452.990 41.280 453.330 41.360 ;
        RECT 463.610 41.280 463.950 41.440 ;
        RECT 442.470 41.230 463.950 41.280 ;
        RECT 441.780 41.010 463.950 41.230 ;
        RECT 441.780 40.830 463.990 41.010 ;
        RECT 441.780 40.780 463.230 40.830 ;
        RECT 442.470 39.380 442.810 40.780 ;
        RECT 447.830 39.420 448.000 39.970 ;
        RECT 452.990 39.710 453.330 40.780 ;
        RECT 452.990 39.450 453.360 39.710 ;
        RECT 458.410 39.450 458.580 39.970 ;
        RECT 442.470 38.350 442.710 39.380 ;
        RECT 442.470 34.500 442.700 38.350 ;
        RECT 442.470 32.880 442.710 34.500 ;
        RECT 442.470 29.030 442.700 32.880 ;
        RECT 442.470 27.410 442.710 29.030 ;
        RECT 442.470 23.560 442.700 27.410 ;
        RECT 442.470 21.940 442.710 23.560 ;
        RECT 436.820 17.840 439.360 18.190 ;
        RECT 442.470 18.090 442.700 21.940 ;
        RECT 414.020 17.080 414.190 17.640 ;
        RECT 392.190 16.040 392.600 16.950 ;
        RECT 402.700 16.070 403.110 17.060 ;
        RECT 413.920 16.070 414.330 17.080 ;
        RECT 424.600 16.940 424.770 17.670 ;
        RECT 435.180 17.050 435.350 17.750 ;
        RECT 442.470 17.720 442.710 18.090 ;
        RECT 402.700 16.040 414.480 16.070 ;
        RECT 381.560 16.030 414.480 16.040 ;
        RECT 424.550 16.030 424.960 16.940 ;
        RECT 435.060 16.030 435.470 17.050 ;
        RECT 442.540 16.470 442.710 17.720 ;
        RECT 447.810 17.610 448.040 39.420 ;
        RECT 453.070 17.720 453.300 39.450 ;
        RECT 447.830 17.050 448.000 17.610 ;
        RECT 381.560 15.590 436.170 16.030 ;
        RECT 381.620 15.560 436.170 15.590 ;
        RECT 392.190 15.450 392.600 15.560 ;
        RECT 402.870 15.550 436.170 15.560 ;
        RECT 447.730 16.000 448.140 17.050 ;
        RECT 453.120 16.470 453.290 17.720 ;
        RECT 458.410 17.640 458.640 39.450 ;
        RECT 463.570 39.430 463.990 40.830 ;
        RECT 468.990 39.530 469.160 39.970 ;
        RECT 463.670 17.860 463.900 39.430 ;
        RECT 458.410 16.910 458.580 17.640 ;
        RECT 458.360 16.000 458.770 16.910 ;
        RECT 463.700 16.470 463.870 17.860 ;
        RECT 468.950 17.720 469.180 39.530 ;
        RECT 470.380 21.210 473.400 125.010 ;
        RECT 474.750 122.260 474.980 126.110 ;
        RECT 474.750 120.640 474.990 122.260 ;
        RECT 474.750 116.790 474.980 120.640 ;
        RECT 474.750 115.170 474.990 116.790 ;
        RECT 474.750 111.320 474.980 115.170 ;
        RECT 474.750 109.700 474.990 111.320 ;
        RECT 474.750 105.850 474.980 109.700 ;
        RECT 474.750 105.480 474.990 105.850 ;
        RECT 474.820 104.230 474.990 105.480 ;
        RECT 480.090 105.370 480.320 127.180 ;
        RECT 485.350 105.480 485.580 127.210 ;
        RECT 480.110 104.810 480.280 105.370 ;
        RECT 480.010 103.760 480.420 104.810 ;
        RECT 485.400 104.230 485.570 105.480 ;
        RECT 490.690 105.400 490.920 127.210 ;
        RECT 495.850 127.190 496.270 128.390 ;
        RECT 495.950 105.620 496.180 127.190 ;
        RECT 500.990 126.850 501.780 128.390 ;
        RECT 490.690 104.670 490.860 105.400 ;
        RECT 490.640 103.760 491.050 104.670 ;
        RECT 495.980 104.230 496.150 105.620 ;
        RECT 501.230 105.480 501.460 126.850 ;
        RECT 501.270 104.780 501.440 105.480 ;
        RECT 503.380 105.230 506.600 127.830 ;
        RECT 501.150 103.760 501.560 104.780 ;
        RECT 480.010 103.310 502.260 103.760 ;
        RECT 480.070 103.280 502.260 103.310 ;
        RECT 490.640 103.170 491.050 103.280 ;
        RECT 474.790 99.920 475.130 99.970 ;
        RECT 485.310 99.920 485.650 100.000 ;
        RECT 495.930 99.920 496.270 100.080 ;
        RECT 474.790 99.870 496.270 99.920 ;
        RECT 474.100 99.650 496.270 99.870 ;
        RECT 474.100 99.470 496.310 99.650 ;
        RECT 474.100 99.420 495.550 99.470 ;
        RECT 474.790 98.020 475.130 99.420 ;
        RECT 480.150 98.060 480.320 98.610 ;
        RECT 485.310 98.350 485.650 99.420 ;
        RECT 485.310 98.090 485.680 98.350 ;
        RECT 490.730 98.090 490.900 98.610 ;
        RECT 474.790 96.990 475.030 98.020 ;
        RECT 474.790 93.140 475.020 96.990 ;
        RECT 474.790 91.520 475.030 93.140 ;
        RECT 474.790 87.670 475.020 91.520 ;
        RECT 474.790 86.050 475.030 87.670 ;
        RECT 474.790 82.200 475.020 86.050 ;
        RECT 474.790 80.580 475.030 82.200 ;
        RECT 474.790 76.730 475.020 80.580 ;
        RECT 474.790 76.360 475.030 76.730 ;
        RECT 474.860 75.110 475.030 76.360 ;
        RECT 480.130 76.250 480.360 98.060 ;
        RECT 485.390 76.360 485.620 98.090 ;
        RECT 480.150 75.690 480.320 76.250 ;
        RECT 480.050 74.640 480.460 75.690 ;
        RECT 485.440 75.110 485.610 76.360 ;
        RECT 490.730 76.280 490.960 98.090 ;
        RECT 495.890 98.070 496.310 99.470 ;
        RECT 501.310 98.170 501.480 98.610 ;
        RECT 495.990 76.500 496.220 98.070 ;
        RECT 490.730 75.550 490.900 76.280 ;
        RECT 490.680 74.640 491.090 75.550 ;
        RECT 496.020 75.110 496.190 76.500 ;
        RECT 501.270 76.360 501.500 98.170 ;
        RECT 501.310 75.660 501.480 76.360 ;
        RECT 501.190 74.640 501.600 75.660 ;
        RECT 480.050 74.190 502.300 74.640 ;
        RECT 503.150 74.400 506.380 96.330 ;
        RECT 480.110 74.160 502.300 74.190 ;
        RECT 490.680 74.050 491.090 74.160 ;
        RECT 474.810 70.560 475.150 70.610 ;
        RECT 485.330 70.560 485.670 70.640 ;
        RECT 495.950 70.560 496.290 70.720 ;
        RECT 474.810 70.510 496.290 70.560 ;
        RECT 474.120 70.290 496.290 70.510 ;
        RECT 474.120 70.110 496.330 70.290 ;
        RECT 474.120 70.060 495.570 70.110 ;
        RECT 474.810 68.660 475.150 70.060 ;
        RECT 480.170 68.700 480.340 69.250 ;
        RECT 485.330 68.990 485.670 70.060 ;
        RECT 485.330 68.730 485.700 68.990 ;
        RECT 490.750 68.730 490.920 69.250 ;
        RECT 474.810 67.630 475.050 68.660 ;
        RECT 474.810 63.780 475.040 67.630 ;
        RECT 474.810 62.160 475.050 63.780 ;
        RECT 474.810 58.310 475.040 62.160 ;
        RECT 474.810 56.690 475.050 58.310 ;
        RECT 474.810 52.840 475.040 56.690 ;
        RECT 474.810 51.220 475.050 52.840 ;
        RECT 474.810 47.370 475.040 51.220 ;
        RECT 474.810 47.000 475.050 47.370 ;
        RECT 474.880 45.750 475.050 47.000 ;
        RECT 480.150 46.890 480.380 68.700 ;
        RECT 485.410 47.000 485.640 68.730 ;
        RECT 480.170 46.330 480.340 46.890 ;
        RECT 480.070 45.280 480.480 46.330 ;
        RECT 485.460 45.750 485.630 47.000 ;
        RECT 490.750 46.920 490.980 68.730 ;
        RECT 495.910 68.710 496.330 70.110 ;
        RECT 501.330 68.810 501.500 69.250 ;
        RECT 496.010 47.140 496.240 68.710 ;
        RECT 490.750 46.190 490.920 46.920 ;
        RECT 490.700 45.280 491.110 46.190 ;
        RECT 496.040 45.750 496.210 47.140 ;
        RECT 501.290 47.000 501.520 68.810 ;
        RECT 501.330 46.300 501.500 47.000 ;
        RECT 503.150 46.470 506.490 69.510 ;
        RECT 501.210 45.280 501.620 46.300 ;
        RECT 480.070 44.830 502.320 45.280 ;
        RECT 480.130 44.800 502.320 44.830 ;
        RECT 490.700 44.690 491.110 44.800 ;
        RECT 474.830 41.270 475.170 41.320 ;
        RECT 485.350 41.270 485.690 41.350 ;
        RECT 495.970 41.270 496.310 41.430 ;
        RECT 474.830 41.220 496.310 41.270 ;
        RECT 474.140 41.000 496.310 41.220 ;
        RECT 474.140 40.820 496.350 41.000 ;
        RECT 474.140 40.770 495.590 40.820 ;
        RECT 474.830 39.370 475.170 40.770 ;
        RECT 480.190 39.410 480.360 39.960 ;
        RECT 485.350 39.700 485.690 40.770 ;
        RECT 485.350 39.440 485.720 39.700 ;
        RECT 490.770 39.440 490.940 39.960 ;
        RECT 474.830 38.340 475.070 39.370 ;
        RECT 474.830 34.490 475.060 38.340 ;
        RECT 474.830 32.870 475.070 34.490 ;
        RECT 474.830 29.020 475.060 32.870 ;
        RECT 474.830 27.400 475.070 29.020 ;
        RECT 474.830 23.550 475.060 27.400 ;
        RECT 474.830 21.930 475.070 23.550 ;
        RECT 474.830 18.080 475.060 21.930 ;
        RECT 468.990 17.020 469.160 17.720 ;
        RECT 474.830 17.710 475.070 18.080 ;
        RECT 468.870 16.030 469.280 17.020 ;
        RECT 474.900 16.460 475.070 17.710 ;
        RECT 480.170 17.600 480.400 39.410 ;
        RECT 485.430 17.710 485.660 39.440 ;
        RECT 480.190 17.040 480.360 17.600 ;
        RECT 480.090 16.030 480.500 17.040 ;
        RECT 485.480 16.460 485.650 17.710 ;
        RECT 490.770 17.630 491.000 39.440 ;
        RECT 495.930 39.420 496.350 40.820 ;
        RECT 501.350 39.520 501.520 39.960 ;
        RECT 496.030 17.850 496.260 39.420 ;
        RECT 490.770 16.900 490.940 17.630 ;
        RECT 468.870 16.000 480.650 16.030 ;
        RECT 447.730 15.990 480.650 16.000 ;
        RECT 490.720 15.990 491.130 16.900 ;
        RECT 496.060 16.460 496.230 17.850 ;
        RECT 501.310 17.710 501.540 39.520 ;
        RECT 501.350 17.010 501.520 17.710 ;
        RECT 501.230 15.990 501.640 17.010 ;
        RECT 447.730 15.550 502.340 15.990 ;
        RECT 503.040 15.860 506.490 38.560 ;
        RECT 402.870 15.520 414.480 15.550 ;
        RECT 424.550 15.440 424.960 15.550 ;
        RECT 447.790 15.520 502.340 15.550 ;
        RECT 458.360 15.410 458.770 15.520 ;
        RECT 469.040 15.510 502.340 15.520 ;
        RECT 469.040 15.480 480.650 15.510 ;
        RECT 490.720 15.400 491.130 15.510 ;
        RECT 368.370 -1.140 379.240 4.020 ;
      LAYER mcon ;
        RECT -97.360 355.395 -97.190 355.565 ;
        RECT -97.360 355.035 -97.190 355.205 ;
        RECT -97.360 354.675 -97.190 354.845 ;
        RECT -97.360 354.315 -97.190 354.485 ;
        RECT -94.780 355.395 -94.610 355.565 ;
        RECT -94.780 355.035 -94.610 355.205 ;
        RECT -94.780 354.675 -94.610 354.845 ;
        RECT -94.780 354.315 -94.610 354.485 ;
        RECT -92.200 355.395 -92.030 355.565 ;
        RECT -92.200 355.035 -92.030 355.205 ;
        RECT -92.200 354.675 -92.030 354.845 ;
        RECT -92.200 354.315 -92.030 354.485 ;
        RECT -89.620 355.395 -89.450 355.565 ;
        RECT -89.620 355.035 -89.450 355.205 ;
        RECT -89.620 354.675 -89.450 354.845 ;
        RECT -89.620 354.315 -89.450 354.485 ;
        RECT -87.040 355.395 -86.870 355.565 ;
        RECT -87.040 355.035 -86.870 355.205 ;
        RECT -87.040 354.675 -86.870 354.845 ;
        RECT -87.040 354.315 -86.870 354.485 ;
        RECT -84.460 355.395 -84.290 355.565 ;
        RECT -84.460 355.035 -84.290 355.205 ;
        RECT -84.460 354.675 -84.290 354.845 ;
        RECT -84.460 354.315 -84.290 354.485 ;
        RECT -81.880 355.395 -81.710 355.565 ;
        RECT -81.880 355.035 -81.710 355.205 ;
        RECT -81.880 354.675 -81.710 354.845 ;
        RECT -81.880 354.315 -81.710 354.485 ;
        RECT -79.300 355.395 -79.130 355.565 ;
        RECT -79.300 355.035 -79.130 355.205 ;
        RECT -79.300 354.675 -79.130 354.845 ;
        RECT -79.300 354.315 -79.130 354.485 ;
        RECT -76.720 355.395 -76.550 355.565 ;
        RECT -76.720 355.035 -76.550 355.205 ;
        RECT -76.720 354.675 -76.550 354.845 ;
        RECT -76.720 354.315 -76.550 354.485 ;
        RECT -74.140 355.395 -73.970 355.565 ;
        RECT -74.140 355.035 -73.970 355.205 ;
        RECT -74.140 354.675 -73.970 354.845 ;
        RECT -74.140 354.315 -73.970 354.485 ;
        RECT -71.560 355.395 -71.390 355.565 ;
        RECT -71.560 355.035 -71.390 355.205 ;
        RECT -71.560 354.675 -71.390 354.845 ;
        RECT -71.560 354.315 -71.390 354.485 ;
        RECT -96.715 352.080 -96.545 352.250 ;
        RECT -95.425 352.080 -95.255 352.250 ;
        RECT -94.135 352.080 -93.965 352.250 ;
        RECT -92.845 352.080 -92.675 352.250 ;
        RECT -91.555 352.080 -91.385 352.250 ;
        RECT -90.265 352.080 -90.095 352.250 ;
        RECT -88.975 352.080 -88.805 352.250 ;
        RECT -87.685 352.080 -87.515 352.250 ;
        RECT -86.395 352.080 -86.225 352.250 ;
        RECT -85.105 352.080 -84.935 352.250 ;
        RECT -83.815 352.080 -83.645 352.250 ;
        RECT -82.525 352.080 -82.355 352.250 ;
        RECT -81.235 352.080 -81.065 352.250 ;
        RECT -79.945 352.080 -79.775 352.250 ;
        RECT -78.655 352.080 -78.485 352.250 ;
        RECT -77.365 352.080 -77.195 352.250 ;
        RECT -76.075 352.080 -75.905 352.250 ;
        RECT -74.785 352.080 -74.615 352.250 ;
        RECT -73.495 352.080 -73.325 352.250 ;
        RECT -72.205 352.080 -72.035 352.250 ;
        RECT -90.810 349.705 -77.680 351.675 ;
        RECT 654.760 351.255 654.930 351.425 ;
        RECT 655.120 351.255 655.290 351.425 ;
        RECT 658.255 351.245 658.425 351.415 ;
        RECT 658.615 351.245 658.785 351.415 ;
        RECT 658.975 351.245 659.145 351.415 ;
        RECT 660.860 351.245 661.030 351.415 ;
        RECT 661.220 351.245 661.390 351.415 ;
        RECT 661.580 351.245 661.750 351.415 ;
        RECT 664.830 351.245 665.000 351.415 ;
        RECT 665.190 351.245 665.360 351.415 ;
        RECT 665.550 351.245 665.720 351.415 ;
        RECT 670.150 351.245 670.320 351.415 ;
        RECT 670.510 351.245 670.680 351.415 ;
        RECT 671.430 351.245 671.600 351.415 ;
        RECT 671.790 351.245 671.960 351.415 ;
        RECT 672.150 351.245 672.320 351.415 ;
        RECT 676.305 351.205 676.475 351.375 ;
        RECT 676.665 351.205 676.835 351.375 ;
        RECT 677.025 351.205 677.195 351.375 ;
        RECT 678.910 351.205 679.080 351.375 ;
        RECT 679.270 351.205 679.440 351.375 ;
        RECT 679.630 351.205 679.800 351.375 ;
        RECT 682.880 351.205 683.050 351.375 ;
        RECT 683.240 351.205 683.410 351.375 ;
        RECT 683.600 351.205 683.770 351.375 ;
        RECT 688.200 351.205 688.370 351.375 ;
        RECT 688.560 351.205 688.730 351.375 ;
        RECT 689.480 351.205 689.650 351.375 ;
        RECT 689.840 351.205 690.010 351.375 ;
        RECT 690.200 351.205 690.370 351.375 ;
        RECT 693.895 351.225 694.065 351.395 ;
        RECT 694.255 351.225 694.425 351.395 ;
        RECT 694.615 351.225 694.785 351.395 ;
        RECT 696.500 351.225 696.670 351.395 ;
        RECT 696.860 351.225 697.030 351.395 ;
        RECT 697.220 351.225 697.390 351.395 ;
        RECT 700.470 351.225 700.640 351.395 ;
        RECT 700.830 351.225 701.000 351.395 ;
        RECT 701.190 351.225 701.360 351.395 ;
        RECT 705.790 351.225 705.960 351.395 ;
        RECT 706.150 351.225 706.320 351.395 ;
        RECT 707.070 351.225 707.240 351.395 ;
        RECT 707.430 351.225 707.600 351.395 ;
        RECT 707.790 351.225 707.960 351.395 ;
        RECT 711.745 351.225 711.915 351.395 ;
        RECT 712.105 351.225 712.275 351.395 ;
        RECT 712.465 351.225 712.635 351.395 ;
        RECT 714.350 351.225 714.520 351.395 ;
        RECT 714.710 351.225 714.880 351.395 ;
        RECT 715.070 351.225 715.240 351.395 ;
        RECT 718.320 351.225 718.490 351.395 ;
        RECT 718.680 351.225 718.850 351.395 ;
        RECT 719.040 351.225 719.210 351.395 ;
        RECT 723.640 351.225 723.810 351.395 ;
        RECT 724.000 351.225 724.170 351.395 ;
        RECT 724.920 351.225 725.090 351.395 ;
        RECT 725.280 351.225 725.450 351.395 ;
        RECT 725.640 351.225 725.810 351.395 ;
        RECT 730.005 351.225 730.175 351.395 ;
        RECT 730.365 351.225 730.535 351.395 ;
        RECT 730.725 351.225 730.895 351.395 ;
        RECT 732.610 351.225 732.780 351.395 ;
        RECT 732.970 351.225 733.140 351.395 ;
        RECT 733.330 351.225 733.500 351.395 ;
        RECT 736.580 351.225 736.750 351.395 ;
        RECT 736.940 351.225 737.110 351.395 ;
        RECT 737.300 351.225 737.470 351.395 ;
        RECT 741.900 351.225 742.070 351.395 ;
        RECT 742.260 351.225 742.430 351.395 ;
        RECT 743.180 351.225 743.350 351.395 ;
        RECT 743.540 351.225 743.710 351.395 ;
        RECT 743.900 351.225 744.070 351.395 ;
        RECT 747.775 351.195 747.945 351.365 ;
        RECT 748.135 351.195 748.305 351.365 ;
        RECT 748.495 351.195 748.665 351.365 ;
        RECT 750.380 351.195 750.550 351.365 ;
        RECT 750.740 351.195 750.910 351.365 ;
        RECT 751.100 351.195 751.270 351.365 ;
        RECT 754.350 351.195 754.520 351.365 ;
        RECT 754.710 351.195 754.880 351.365 ;
        RECT 755.070 351.195 755.240 351.365 ;
        RECT 759.670 351.195 759.840 351.365 ;
        RECT 760.030 351.195 760.200 351.365 ;
        RECT 760.950 351.195 761.120 351.365 ;
        RECT 761.310 351.195 761.480 351.365 ;
        RECT 761.670 351.195 761.840 351.365 ;
        RECT 765.815 351.115 765.985 351.285 ;
        RECT 766.175 351.115 766.345 351.285 ;
        RECT 766.535 351.115 766.705 351.285 ;
        RECT 768.420 351.115 768.590 351.285 ;
        RECT 768.780 351.115 768.950 351.285 ;
        RECT 769.140 351.115 769.310 351.285 ;
        RECT 772.390 351.115 772.560 351.285 ;
        RECT 772.750 351.115 772.920 351.285 ;
        RECT 773.110 351.115 773.280 351.285 ;
        RECT 777.710 351.115 777.880 351.285 ;
        RECT 778.070 351.115 778.240 351.285 ;
        RECT 778.990 351.115 779.160 351.285 ;
        RECT 779.350 351.115 779.520 351.285 ;
        RECT 779.710 351.115 779.880 351.285 ;
        RECT 783.975 351.155 784.145 351.325 ;
        RECT 784.335 351.155 784.505 351.325 ;
        RECT 784.695 351.155 784.865 351.325 ;
        RECT 786.580 351.155 786.750 351.325 ;
        RECT 786.940 351.155 787.110 351.325 ;
        RECT 787.300 351.155 787.470 351.325 ;
        RECT 790.550 351.155 790.720 351.325 ;
        RECT 790.910 351.155 791.080 351.325 ;
        RECT 791.270 351.155 791.440 351.325 ;
        RECT 795.870 351.155 796.040 351.325 ;
        RECT 796.230 351.155 796.400 351.325 ;
        RECT 797.150 351.155 797.320 351.325 ;
        RECT 797.510 351.155 797.680 351.325 ;
        RECT 797.870 351.155 798.040 351.325 ;
        RECT 802.355 351.165 802.525 351.335 ;
        RECT 802.715 351.165 802.885 351.335 ;
        RECT 803.075 351.165 803.245 351.335 ;
        RECT 804.960 351.165 805.130 351.335 ;
        RECT 805.320 351.165 805.490 351.335 ;
        RECT 805.680 351.165 805.850 351.335 ;
        RECT 808.930 351.165 809.100 351.335 ;
        RECT 809.290 351.165 809.460 351.335 ;
        RECT 809.650 351.165 809.820 351.335 ;
        RECT 814.250 351.165 814.420 351.335 ;
        RECT 814.610 351.165 814.780 351.335 ;
        RECT 815.530 351.165 815.700 351.335 ;
        RECT 815.890 351.165 816.060 351.335 ;
        RECT 816.250 351.165 816.420 351.335 ;
        RECT 821.155 351.145 821.325 351.315 ;
        RECT 821.515 351.145 821.685 351.315 ;
        RECT 821.875 351.145 822.045 351.315 ;
        RECT 823.760 351.145 823.930 351.315 ;
        RECT 824.120 351.145 824.290 351.315 ;
        RECT 824.480 351.145 824.650 351.315 ;
        RECT 827.730 351.145 827.900 351.315 ;
        RECT 828.090 351.145 828.260 351.315 ;
        RECT 828.450 351.145 828.620 351.315 ;
        RECT 833.050 351.145 833.220 351.315 ;
        RECT 833.410 351.145 833.580 351.315 ;
        RECT 834.330 351.145 834.500 351.315 ;
        RECT 834.690 351.145 834.860 351.315 ;
        RECT 835.050 351.145 835.220 351.315 ;
        RECT 839.710 351.125 839.880 351.295 ;
        RECT 840.070 351.125 840.240 351.295 ;
        RECT 654.125 350.775 654.295 350.945 ;
        RECT 654.605 350.775 654.775 350.945 ;
        RECT 655.085 350.775 655.255 350.945 ;
        RECT 657.705 350.765 657.875 350.935 ;
        RECT 658.185 350.765 658.355 350.935 ;
        RECT 658.665 350.765 658.835 350.935 ;
        RECT 659.145 350.765 659.315 350.935 ;
        RECT 659.625 350.765 659.795 350.935 ;
        RECT 660.105 350.765 660.275 350.935 ;
        RECT 660.585 350.765 660.755 350.935 ;
        RECT 661.065 350.765 661.235 350.935 ;
        RECT 661.545 350.765 661.715 350.935 ;
        RECT 662.025 350.765 662.195 350.935 ;
        RECT 662.505 350.765 662.675 350.935 ;
        RECT 662.985 350.765 663.155 350.935 ;
        RECT 663.465 350.765 663.635 350.935 ;
        RECT 663.945 350.765 664.115 350.935 ;
        RECT 664.425 350.765 664.595 350.935 ;
        RECT 664.905 350.765 665.075 350.935 ;
        RECT 665.385 350.765 665.555 350.935 ;
        RECT 665.865 350.765 666.035 350.935 ;
        RECT 666.345 350.765 666.515 350.935 ;
        RECT 666.825 350.765 666.995 350.935 ;
        RECT 667.305 350.765 667.475 350.935 ;
        RECT 667.785 350.765 667.955 350.935 ;
        RECT 668.265 350.765 668.435 350.935 ;
        RECT 668.745 350.765 668.915 350.935 ;
        RECT 669.225 350.765 669.395 350.935 ;
        RECT 669.705 350.765 669.875 350.935 ;
        RECT 670.185 350.765 670.355 350.935 ;
        RECT 670.665 350.765 670.835 350.935 ;
        RECT 671.145 350.765 671.315 350.935 ;
        RECT 671.625 350.765 671.795 350.935 ;
        RECT 672.105 350.765 672.275 350.935 ;
        RECT 672.585 350.765 672.755 350.935 ;
        RECT 675.755 350.725 675.925 350.895 ;
        RECT 676.235 350.725 676.405 350.895 ;
        RECT 676.715 350.725 676.885 350.895 ;
        RECT 677.195 350.725 677.365 350.895 ;
        RECT 677.675 350.725 677.845 350.895 ;
        RECT 678.155 350.725 678.325 350.895 ;
        RECT 678.635 350.725 678.805 350.895 ;
        RECT 679.115 350.725 679.285 350.895 ;
        RECT 679.595 350.725 679.765 350.895 ;
        RECT 680.075 350.725 680.245 350.895 ;
        RECT 680.555 350.725 680.725 350.895 ;
        RECT 681.035 350.725 681.205 350.895 ;
        RECT 681.515 350.725 681.685 350.895 ;
        RECT 681.995 350.725 682.165 350.895 ;
        RECT 682.475 350.725 682.645 350.895 ;
        RECT 682.955 350.725 683.125 350.895 ;
        RECT 683.435 350.725 683.605 350.895 ;
        RECT 683.915 350.725 684.085 350.895 ;
        RECT 684.395 350.725 684.565 350.895 ;
        RECT 684.875 350.725 685.045 350.895 ;
        RECT 685.355 350.725 685.525 350.895 ;
        RECT 685.835 350.725 686.005 350.895 ;
        RECT 686.315 350.725 686.485 350.895 ;
        RECT 686.795 350.725 686.965 350.895 ;
        RECT 687.275 350.725 687.445 350.895 ;
        RECT 687.755 350.725 687.925 350.895 ;
        RECT 688.235 350.725 688.405 350.895 ;
        RECT 688.715 350.725 688.885 350.895 ;
        RECT 689.195 350.725 689.365 350.895 ;
        RECT 689.675 350.725 689.845 350.895 ;
        RECT 690.155 350.725 690.325 350.895 ;
        RECT 690.635 350.725 690.805 350.895 ;
        RECT 693.345 350.745 693.515 350.915 ;
        RECT 693.825 350.745 693.995 350.915 ;
        RECT 694.305 350.745 694.475 350.915 ;
        RECT 694.785 350.745 694.955 350.915 ;
        RECT 695.265 350.745 695.435 350.915 ;
        RECT 695.745 350.745 695.915 350.915 ;
        RECT 696.225 350.745 696.395 350.915 ;
        RECT 696.705 350.745 696.875 350.915 ;
        RECT 697.185 350.745 697.355 350.915 ;
        RECT 697.665 350.745 697.835 350.915 ;
        RECT 698.145 350.745 698.315 350.915 ;
        RECT 698.625 350.745 698.795 350.915 ;
        RECT 699.105 350.745 699.275 350.915 ;
        RECT 699.585 350.745 699.755 350.915 ;
        RECT 700.065 350.745 700.235 350.915 ;
        RECT 700.545 350.745 700.715 350.915 ;
        RECT 701.025 350.745 701.195 350.915 ;
        RECT 701.505 350.745 701.675 350.915 ;
        RECT 701.985 350.745 702.155 350.915 ;
        RECT 702.465 350.745 702.635 350.915 ;
        RECT 702.945 350.745 703.115 350.915 ;
        RECT 703.425 350.745 703.595 350.915 ;
        RECT 703.905 350.745 704.075 350.915 ;
        RECT 704.385 350.745 704.555 350.915 ;
        RECT 704.865 350.745 705.035 350.915 ;
        RECT 705.345 350.745 705.515 350.915 ;
        RECT 705.825 350.745 705.995 350.915 ;
        RECT 706.305 350.745 706.475 350.915 ;
        RECT 706.785 350.745 706.955 350.915 ;
        RECT 707.265 350.745 707.435 350.915 ;
        RECT 707.745 350.745 707.915 350.915 ;
        RECT 708.225 350.745 708.395 350.915 ;
        RECT 711.195 350.745 711.365 350.915 ;
        RECT 711.675 350.745 711.845 350.915 ;
        RECT 712.155 350.745 712.325 350.915 ;
        RECT 712.635 350.745 712.805 350.915 ;
        RECT 713.115 350.745 713.285 350.915 ;
        RECT 713.595 350.745 713.765 350.915 ;
        RECT 714.075 350.745 714.245 350.915 ;
        RECT 714.555 350.745 714.725 350.915 ;
        RECT 715.035 350.745 715.205 350.915 ;
        RECT 715.515 350.745 715.685 350.915 ;
        RECT 715.995 350.745 716.165 350.915 ;
        RECT 716.475 350.745 716.645 350.915 ;
        RECT 716.955 350.745 717.125 350.915 ;
        RECT 717.435 350.745 717.605 350.915 ;
        RECT 717.915 350.745 718.085 350.915 ;
        RECT 718.395 350.745 718.565 350.915 ;
        RECT 718.875 350.745 719.045 350.915 ;
        RECT 719.355 350.745 719.525 350.915 ;
        RECT 719.835 350.745 720.005 350.915 ;
        RECT 720.315 350.745 720.485 350.915 ;
        RECT 720.795 350.745 720.965 350.915 ;
        RECT 721.275 350.745 721.445 350.915 ;
        RECT 721.755 350.745 721.925 350.915 ;
        RECT 722.235 350.745 722.405 350.915 ;
        RECT 722.715 350.745 722.885 350.915 ;
        RECT 723.195 350.745 723.365 350.915 ;
        RECT 723.675 350.745 723.845 350.915 ;
        RECT 724.155 350.745 724.325 350.915 ;
        RECT 724.635 350.745 724.805 350.915 ;
        RECT 725.115 350.745 725.285 350.915 ;
        RECT 725.595 350.745 725.765 350.915 ;
        RECT 726.075 350.745 726.245 350.915 ;
        RECT 729.455 350.745 729.625 350.915 ;
        RECT 729.935 350.745 730.105 350.915 ;
        RECT 730.415 350.745 730.585 350.915 ;
        RECT 730.895 350.745 731.065 350.915 ;
        RECT 731.375 350.745 731.545 350.915 ;
        RECT 731.855 350.745 732.025 350.915 ;
        RECT 732.335 350.745 732.505 350.915 ;
        RECT 732.815 350.745 732.985 350.915 ;
        RECT 733.295 350.745 733.465 350.915 ;
        RECT 733.775 350.745 733.945 350.915 ;
        RECT 734.255 350.745 734.425 350.915 ;
        RECT 734.735 350.745 734.905 350.915 ;
        RECT 735.215 350.745 735.385 350.915 ;
        RECT 735.695 350.745 735.865 350.915 ;
        RECT 736.175 350.745 736.345 350.915 ;
        RECT 736.655 350.745 736.825 350.915 ;
        RECT 737.135 350.745 737.305 350.915 ;
        RECT 737.615 350.745 737.785 350.915 ;
        RECT 738.095 350.745 738.265 350.915 ;
        RECT 738.575 350.745 738.745 350.915 ;
        RECT 739.055 350.745 739.225 350.915 ;
        RECT 739.535 350.745 739.705 350.915 ;
        RECT 740.015 350.745 740.185 350.915 ;
        RECT 740.495 350.745 740.665 350.915 ;
        RECT 740.975 350.745 741.145 350.915 ;
        RECT 741.455 350.745 741.625 350.915 ;
        RECT 741.935 350.745 742.105 350.915 ;
        RECT 742.415 350.745 742.585 350.915 ;
        RECT 742.895 350.745 743.065 350.915 ;
        RECT 743.375 350.745 743.545 350.915 ;
        RECT 743.855 350.745 744.025 350.915 ;
        RECT 744.335 350.745 744.505 350.915 ;
        RECT 747.225 350.715 747.395 350.885 ;
        RECT 747.705 350.715 747.875 350.885 ;
        RECT 748.185 350.715 748.355 350.885 ;
        RECT 748.665 350.715 748.835 350.885 ;
        RECT 749.145 350.715 749.315 350.885 ;
        RECT 749.625 350.715 749.795 350.885 ;
        RECT 750.105 350.715 750.275 350.885 ;
        RECT 750.585 350.715 750.755 350.885 ;
        RECT 751.065 350.715 751.235 350.885 ;
        RECT 751.545 350.715 751.715 350.885 ;
        RECT 752.025 350.715 752.195 350.885 ;
        RECT 752.505 350.715 752.675 350.885 ;
        RECT 752.985 350.715 753.155 350.885 ;
        RECT 753.465 350.715 753.635 350.885 ;
        RECT 753.945 350.715 754.115 350.885 ;
        RECT 754.425 350.715 754.595 350.885 ;
        RECT 754.905 350.715 755.075 350.885 ;
        RECT 755.385 350.715 755.555 350.885 ;
        RECT 755.865 350.715 756.035 350.885 ;
        RECT 756.345 350.715 756.515 350.885 ;
        RECT 756.825 350.715 756.995 350.885 ;
        RECT 757.305 350.715 757.475 350.885 ;
        RECT 757.785 350.715 757.955 350.885 ;
        RECT 758.265 350.715 758.435 350.885 ;
        RECT 758.745 350.715 758.915 350.885 ;
        RECT 759.225 350.715 759.395 350.885 ;
        RECT 759.705 350.715 759.875 350.885 ;
        RECT 760.185 350.715 760.355 350.885 ;
        RECT 760.665 350.715 760.835 350.885 ;
        RECT 761.145 350.715 761.315 350.885 ;
        RECT 761.625 350.715 761.795 350.885 ;
        RECT 762.105 350.715 762.275 350.885 ;
        RECT 765.265 350.635 765.435 350.805 ;
        RECT 765.745 350.635 765.915 350.805 ;
        RECT 766.225 350.635 766.395 350.805 ;
        RECT 766.705 350.635 766.875 350.805 ;
        RECT 767.185 350.635 767.355 350.805 ;
        RECT 767.665 350.635 767.835 350.805 ;
        RECT 768.145 350.635 768.315 350.805 ;
        RECT 768.625 350.635 768.795 350.805 ;
        RECT 769.105 350.635 769.275 350.805 ;
        RECT 769.585 350.635 769.755 350.805 ;
        RECT 770.065 350.635 770.235 350.805 ;
        RECT 770.545 350.635 770.715 350.805 ;
        RECT 771.025 350.635 771.195 350.805 ;
        RECT 771.505 350.635 771.675 350.805 ;
        RECT 771.985 350.635 772.155 350.805 ;
        RECT 772.465 350.635 772.635 350.805 ;
        RECT 772.945 350.635 773.115 350.805 ;
        RECT 773.425 350.635 773.595 350.805 ;
        RECT 773.905 350.635 774.075 350.805 ;
        RECT 774.385 350.635 774.555 350.805 ;
        RECT 774.865 350.635 775.035 350.805 ;
        RECT 775.345 350.635 775.515 350.805 ;
        RECT 775.825 350.635 775.995 350.805 ;
        RECT 776.305 350.635 776.475 350.805 ;
        RECT 776.785 350.635 776.955 350.805 ;
        RECT 777.265 350.635 777.435 350.805 ;
        RECT 777.745 350.635 777.915 350.805 ;
        RECT 778.225 350.635 778.395 350.805 ;
        RECT 778.705 350.635 778.875 350.805 ;
        RECT 779.185 350.635 779.355 350.805 ;
        RECT 779.665 350.635 779.835 350.805 ;
        RECT 780.145 350.635 780.315 350.805 ;
        RECT 783.425 350.675 783.595 350.845 ;
        RECT 783.905 350.675 784.075 350.845 ;
        RECT 784.385 350.675 784.555 350.845 ;
        RECT 784.865 350.675 785.035 350.845 ;
        RECT 785.345 350.675 785.515 350.845 ;
        RECT 785.825 350.675 785.995 350.845 ;
        RECT 786.305 350.675 786.475 350.845 ;
        RECT 786.785 350.675 786.955 350.845 ;
        RECT 787.265 350.675 787.435 350.845 ;
        RECT 787.745 350.675 787.915 350.845 ;
        RECT 788.225 350.675 788.395 350.845 ;
        RECT 788.705 350.675 788.875 350.845 ;
        RECT 789.185 350.675 789.355 350.845 ;
        RECT 789.665 350.675 789.835 350.845 ;
        RECT 790.145 350.675 790.315 350.845 ;
        RECT 790.625 350.675 790.795 350.845 ;
        RECT 791.105 350.675 791.275 350.845 ;
        RECT 791.585 350.675 791.755 350.845 ;
        RECT 792.065 350.675 792.235 350.845 ;
        RECT 792.545 350.675 792.715 350.845 ;
        RECT 793.025 350.675 793.195 350.845 ;
        RECT 793.505 350.675 793.675 350.845 ;
        RECT 793.985 350.675 794.155 350.845 ;
        RECT 794.465 350.675 794.635 350.845 ;
        RECT 794.945 350.675 795.115 350.845 ;
        RECT 795.425 350.675 795.595 350.845 ;
        RECT 795.905 350.675 796.075 350.845 ;
        RECT 796.385 350.675 796.555 350.845 ;
        RECT 796.865 350.675 797.035 350.845 ;
        RECT 797.345 350.675 797.515 350.845 ;
        RECT 797.825 350.675 797.995 350.845 ;
        RECT 798.305 350.675 798.475 350.845 ;
        RECT 801.805 350.685 801.975 350.855 ;
        RECT 802.285 350.685 802.455 350.855 ;
        RECT 802.765 350.685 802.935 350.855 ;
        RECT 803.245 350.685 803.415 350.855 ;
        RECT 803.725 350.685 803.895 350.855 ;
        RECT 804.205 350.685 804.375 350.855 ;
        RECT 804.685 350.685 804.855 350.855 ;
        RECT 805.165 350.685 805.335 350.855 ;
        RECT 805.645 350.685 805.815 350.855 ;
        RECT 806.125 350.685 806.295 350.855 ;
        RECT 806.605 350.685 806.775 350.855 ;
        RECT 807.085 350.685 807.255 350.855 ;
        RECT 807.565 350.685 807.735 350.855 ;
        RECT 808.045 350.685 808.215 350.855 ;
        RECT 808.525 350.685 808.695 350.855 ;
        RECT 809.005 350.685 809.175 350.855 ;
        RECT 809.485 350.685 809.655 350.855 ;
        RECT 809.965 350.685 810.135 350.855 ;
        RECT 810.445 350.685 810.615 350.855 ;
        RECT 810.925 350.685 811.095 350.855 ;
        RECT 811.405 350.685 811.575 350.855 ;
        RECT 811.885 350.685 812.055 350.855 ;
        RECT 812.365 350.685 812.535 350.855 ;
        RECT 812.845 350.685 813.015 350.855 ;
        RECT 813.325 350.685 813.495 350.855 ;
        RECT 813.805 350.685 813.975 350.855 ;
        RECT 814.285 350.685 814.455 350.855 ;
        RECT 814.765 350.685 814.935 350.855 ;
        RECT 815.245 350.685 815.415 350.855 ;
        RECT 815.725 350.685 815.895 350.855 ;
        RECT 816.205 350.685 816.375 350.855 ;
        RECT 816.685 350.685 816.855 350.855 ;
        RECT 820.605 350.665 820.775 350.835 ;
        RECT 821.085 350.665 821.255 350.835 ;
        RECT 821.565 350.665 821.735 350.835 ;
        RECT 822.045 350.665 822.215 350.835 ;
        RECT 822.525 350.665 822.695 350.835 ;
        RECT 823.005 350.665 823.175 350.835 ;
        RECT 823.485 350.665 823.655 350.835 ;
        RECT 823.965 350.665 824.135 350.835 ;
        RECT 824.445 350.665 824.615 350.835 ;
        RECT 824.925 350.665 825.095 350.835 ;
        RECT 825.405 350.665 825.575 350.835 ;
        RECT 825.885 350.665 826.055 350.835 ;
        RECT 826.365 350.665 826.535 350.835 ;
        RECT 826.845 350.665 827.015 350.835 ;
        RECT 827.325 350.665 827.495 350.835 ;
        RECT 827.805 350.665 827.975 350.835 ;
        RECT 828.285 350.665 828.455 350.835 ;
        RECT 828.765 350.665 828.935 350.835 ;
        RECT 829.245 350.665 829.415 350.835 ;
        RECT 829.725 350.665 829.895 350.835 ;
        RECT 830.205 350.665 830.375 350.835 ;
        RECT 830.685 350.665 830.855 350.835 ;
        RECT 831.165 350.665 831.335 350.835 ;
        RECT 831.645 350.665 831.815 350.835 ;
        RECT 832.125 350.665 832.295 350.835 ;
        RECT 832.605 350.665 832.775 350.835 ;
        RECT 833.085 350.665 833.255 350.835 ;
        RECT 833.565 350.665 833.735 350.835 ;
        RECT 834.045 350.665 834.215 350.835 ;
        RECT 834.525 350.665 834.695 350.835 ;
        RECT 835.005 350.665 835.175 350.835 ;
        RECT 835.485 350.665 835.655 350.835 ;
        RECT 839.075 350.645 839.245 350.815 ;
        RECT 839.555 350.645 839.725 350.815 ;
        RECT 840.035 350.645 840.205 350.815 ;
        RECT 784.615 342.985 784.785 343.155 ;
        RECT 784.975 342.985 785.145 343.155 ;
        RECT 785.335 342.985 785.505 343.155 ;
        RECT 791.180 343.015 791.350 343.185 ;
        RECT 791.540 343.015 791.710 343.185 ;
        RECT 794.555 343.075 794.725 343.245 ;
        RECT 794.915 343.075 795.085 343.245 ;
        RECT 795.275 343.075 795.445 343.245 ;
        RECT 797.160 343.075 797.330 343.245 ;
        RECT 797.520 343.075 797.690 343.245 ;
        RECT 797.880 343.075 798.050 343.245 ;
        RECT 801.130 343.075 801.300 343.245 ;
        RECT 801.490 343.075 801.660 343.245 ;
        RECT 801.850 343.075 802.020 343.245 ;
        RECT 806.450 343.075 806.620 343.245 ;
        RECT 806.810 343.075 806.980 343.245 ;
        RECT 807.730 343.075 807.900 343.245 ;
        RECT 808.090 343.075 808.260 343.245 ;
        RECT 808.450 343.075 808.620 343.245 ;
        RECT 813.915 342.985 814.085 343.155 ;
        RECT 814.275 342.985 814.445 343.155 ;
        RECT 814.635 342.985 814.805 343.155 ;
        RECT 816.520 342.985 816.690 343.155 ;
        RECT 816.880 342.985 817.050 343.155 ;
        RECT 817.240 342.985 817.410 343.155 ;
        RECT 820.490 342.985 820.660 343.155 ;
        RECT 820.850 342.985 821.020 343.155 ;
        RECT 821.210 342.985 821.380 343.155 ;
        RECT 825.810 342.985 825.980 343.155 ;
        RECT 826.170 342.985 826.340 343.155 ;
        RECT 827.090 342.985 827.260 343.155 ;
        RECT 827.450 342.985 827.620 343.155 ;
        RECT 827.810 342.985 827.980 343.155 ;
        RECT 783.985 342.505 784.155 342.675 ;
        RECT 784.465 342.505 784.635 342.675 ;
        RECT 784.945 342.505 785.115 342.675 ;
        RECT 785.425 342.505 785.595 342.675 ;
        RECT 785.905 342.505 786.075 342.675 ;
        RECT 786.385 342.505 786.555 342.675 ;
        RECT 786.865 342.505 787.035 342.675 ;
        RECT 790.545 342.535 790.715 342.705 ;
        RECT 791.025 342.535 791.195 342.705 ;
        RECT 791.505 342.535 791.675 342.705 ;
        RECT 794.005 342.595 794.175 342.765 ;
        RECT 794.485 342.595 794.655 342.765 ;
        RECT 794.965 342.595 795.135 342.765 ;
        RECT 795.445 342.595 795.615 342.765 ;
        RECT 795.925 342.595 796.095 342.765 ;
        RECT 796.405 342.595 796.575 342.765 ;
        RECT 796.885 342.595 797.055 342.765 ;
        RECT 797.365 342.595 797.535 342.765 ;
        RECT 797.845 342.595 798.015 342.765 ;
        RECT 798.325 342.595 798.495 342.765 ;
        RECT 798.805 342.595 798.975 342.765 ;
        RECT 799.285 342.595 799.455 342.765 ;
        RECT 799.765 342.595 799.935 342.765 ;
        RECT 800.245 342.595 800.415 342.765 ;
        RECT 800.725 342.595 800.895 342.765 ;
        RECT 801.205 342.595 801.375 342.765 ;
        RECT 801.685 342.595 801.855 342.765 ;
        RECT 802.165 342.595 802.335 342.765 ;
        RECT 802.645 342.595 802.815 342.765 ;
        RECT 803.125 342.595 803.295 342.765 ;
        RECT 803.605 342.595 803.775 342.765 ;
        RECT 804.085 342.595 804.255 342.765 ;
        RECT 804.565 342.595 804.735 342.765 ;
        RECT 805.045 342.595 805.215 342.765 ;
        RECT 805.525 342.595 805.695 342.765 ;
        RECT 806.005 342.595 806.175 342.765 ;
        RECT 806.485 342.595 806.655 342.765 ;
        RECT 806.965 342.595 807.135 342.765 ;
        RECT 807.445 342.595 807.615 342.765 ;
        RECT 807.925 342.595 808.095 342.765 ;
        RECT 808.405 342.595 808.575 342.765 ;
        RECT 808.885 342.595 809.055 342.765 ;
        RECT 813.365 342.505 813.535 342.675 ;
        RECT 813.845 342.505 814.015 342.675 ;
        RECT 814.325 342.505 814.495 342.675 ;
        RECT 814.805 342.505 814.975 342.675 ;
        RECT 815.285 342.505 815.455 342.675 ;
        RECT 815.765 342.505 815.935 342.675 ;
        RECT 816.245 342.505 816.415 342.675 ;
        RECT 816.725 342.505 816.895 342.675 ;
        RECT 817.205 342.505 817.375 342.675 ;
        RECT 817.685 342.505 817.855 342.675 ;
        RECT 818.165 342.505 818.335 342.675 ;
        RECT 818.645 342.505 818.815 342.675 ;
        RECT 819.125 342.505 819.295 342.675 ;
        RECT 819.605 342.505 819.775 342.675 ;
        RECT 820.085 342.505 820.255 342.675 ;
        RECT 820.565 342.505 820.735 342.675 ;
        RECT 821.045 342.505 821.215 342.675 ;
        RECT 821.525 342.505 821.695 342.675 ;
        RECT 822.005 342.505 822.175 342.675 ;
        RECT 822.485 342.505 822.655 342.675 ;
        RECT 822.965 342.505 823.135 342.675 ;
        RECT 823.445 342.505 823.615 342.675 ;
        RECT 823.925 342.505 824.095 342.675 ;
        RECT 824.405 342.505 824.575 342.675 ;
        RECT 824.885 342.505 825.055 342.675 ;
        RECT 825.365 342.505 825.535 342.675 ;
        RECT 825.845 342.505 826.015 342.675 ;
        RECT 826.325 342.505 826.495 342.675 ;
        RECT 826.805 342.505 826.975 342.675 ;
        RECT 827.285 342.505 827.455 342.675 ;
        RECT 827.765 342.505 827.935 342.675 ;
        RECT 828.245 342.505 828.415 342.675 ;
        RECT 853.910 337.645 854.080 337.815 ;
        RECT 853.910 336.175 854.080 336.345 ;
        RECT 853.910 334.705 854.080 334.875 ;
        RECT 853.910 333.235 854.080 333.405 ;
        RECT 853.910 331.765 854.080 331.935 ;
        RECT 853.910 330.295 854.080 330.465 ;
        RECT 664.875 328.895 665.045 329.065 ;
        RECT 665.235 328.895 665.405 329.065 ;
        RECT 665.595 328.895 665.765 329.065 ;
        RECT 670.505 328.895 670.675 329.065 ;
        RECT 670.865 328.895 671.035 329.065 ;
        RECT 671.225 328.895 671.395 329.065 ;
        RECT 674.680 328.795 674.850 328.965 ;
        RECT 675.040 328.795 675.210 328.965 ;
        RECT 675.400 328.795 675.570 328.965 ;
        RECT 676.650 328.795 676.820 328.965 ;
        RECT 677.010 328.795 677.180 328.965 ;
        RECT 684.095 328.835 684.265 329.005 ;
        RECT 684.625 328.835 684.795 329.005 ;
        RECT 689.155 328.845 689.325 329.015 ;
        RECT 689.515 328.845 689.685 329.015 ;
        RECT 689.875 328.845 690.045 329.015 ;
        RECT 853.910 328.825 854.080 328.995 ;
        RECT 635.380 327.555 635.550 327.725 ;
        RECT 635.740 327.555 635.910 327.725 ;
        RECT 639.570 327.645 639.740 327.815 ;
        RECT 639.930 327.645 640.100 327.815 ;
        RECT 643.670 327.625 643.840 327.795 ;
        RECT 644.030 327.625 644.200 327.795 ;
        RECT 596.160 327.105 596.330 327.275 ;
        RECT 596.520 327.105 596.690 327.275 ;
        RECT 595.525 326.625 595.695 326.795 ;
        RECT 596.005 326.625 596.175 326.795 ;
        RECT 596.485 326.625 596.655 326.795 ;
        RECT 596.630 325.905 596.800 326.075 ;
        RECT 596.990 325.905 597.160 326.075 ;
        RECT 605.495 322.895 606.025 326.305 ;
        RECT 635.415 327.075 635.585 327.245 ;
        RECT 635.895 327.075 636.065 327.245 ;
        RECT 636.375 327.075 636.545 327.245 ;
        RECT 639.605 327.165 639.775 327.335 ;
        RECT 640.085 327.165 640.255 327.335 ;
        RECT 640.565 327.165 640.735 327.335 ;
        RECT 643.705 327.145 643.875 327.315 ;
        RECT 644.185 327.145 644.355 327.315 ;
        RECT 644.665 327.145 644.835 327.315 ;
        RECT 663.345 328.415 663.515 328.585 ;
        RECT 663.825 328.415 663.995 328.585 ;
        RECT 664.305 328.415 664.475 328.585 ;
        RECT 664.785 328.415 664.955 328.585 ;
        RECT 665.265 328.415 665.435 328.585 ;
        RECT 665.745 328.415 665.915 328.585 ;
        RECT 666.225 328.415 666.395 328.585 ;
        RECT 668.975 328.415 669.145 328.585 ;
        RECT 669.455 328.415 669.625 328.585 ;
        RECT 669.935 328.415 670.105 328.585 ;
        RECT 670.415 328.415 670.585 328.585 ;
        RECT 670.895 328.415 671.065 328.585 ;
        RECT 671.375 328.415 671.545 328.585 ;
        RECT 671.855 328.415 672.025 328.585 ;
        RECT 674.735 328.315 674.905 328.485 ;
        RECT 675.215 328.315 675.385 328.485 ;
        RECT 675.695 328.315 675.865 328.485 ;
        RECT 676.175 328.315 676.345 328.485 ;
        RECT 676.655 328.315 676.825 328.485 ;
        RECT 677.135 328.315 677.305 328.485 ;
        RECT 677.615 328.315 677.785 328.485 ;
        RECT 681.765 328.355 681.935 328.525 ;
        RECT 682.245 328.355 682.415 328.525 ;
        RECT 682.725 328.355 682.895 328.525 ;
        RECT 683.205 328.355 683.375 328.525 ;
        RECT 683.685 328.355 683.855 328.525 ;
        RECT 684.165 328.355 684.335 328.525 ;
        RECT 684.645 328.355 684.815 328.525 ;
        RECT 685.125 328.355 685.295 328.525 ;
        RECT 687.625 328.365 687.795 328.535 ;
        RECT 688.105 328.365 688.275 328.535 ;
        RECT 688.585 328.365 688.755 328.535 ;
        RECT 689.065 328.365 689.235 328.535 ;
        RECT 689.545 328.365 689.715 328.535 ;
        RECT 690.025 328.365 690.195 328.535 ;
        RECT 690.505 328.365 690.675 328.535 ;
        RECT 625.900 326.235 626.070 326.405 ;
        RECT 625.900 325.875 626.070 326.045 ;
        RECT 625.900 325.515 626.070 325.685 ;
        RECT 625.900 325.155 626.070 325.325 ;
        RECT 625.900 324.795 626.070 324.965 ;
        RECT 615.020 324.425 615.190 324.595 ;
        RECT 616.600 324.425 616.770 324.595 ;
        RECT 625.900 324.435 626.070 324.605 ;
        RECT 625.900 324.075 626.070 324.245 ;
        RECT 625.900 323.715 626.070 323.885 ;
        RECT 853.910 327.355 854.080 327.525 ;
        RECT 851.745 326.540 851.915 326.710 ;
        RECT 851.745 326.180 851.915 326.350 ;
        RECT 851.745 325.820 851.915 325.990 ;
        RECT 853.910 325.885 854.080 326.055 ;
        RECT 851.745 325.460 851.915 325.630 ;
        RECT 851.745 325.100 851.915 325.270 ;
        RECT 851.745 324.740 851.915 324.910 ;
        RECT 851.745 324.380 851.915 324.550 ;
        RECT 853.910 324.415 854.080 324.585 ;
        RECT 851.745 324.020 851.915 324.190 ;
        RECT 625.900 323.355 626.070 323.525 ;
        RECT 640.370 323.535 640.540 323.705 ;
        RECT 644.420 323.585 644.590 323.755 ;
        RECT 851.745 323.660 851.915 323.830 ;
        RECT 615.020 322.955 615.190 323.125 ;
        RECT 616.600 322.955 616.770 323.125 ;
        RECT 658.880 322.595 659.050 322.765 ;
        RECT 659.240 322.595 659.410 322.765 ;
        RECT 663.780 322.555 663.950 322.725 ;
        RECT 664.140 322.555 664.310 322.725 ;
        RECT 668.370 322.585 668.540 322.755 ;
        RECT 668.730 322.585 668.900 322.755 ;
        RECT 672.910 322.565 673.080 322.735 ;
        RECT 673.270 322.565 673.440 322.735 ;
        RECT 678.705 322.575 678.875 322.745 ;
        RECT 679.235 322.575 679.405 322.745 ;
        RECT 683.675 322.575 683.845 322.745 ;
        RECT 684.035 322.575 684.205 322.745 ;
        RECT 684.395 322.575 684.565 322.745 ;
        RECT 689.125 322.575 689.295 322.745 ;
        RECT 689.485 322.575 689.655 322.745 ;
        RECT 689.845 322.575 690.015 322.745 ;
        RECT 692.850 322.595 693.020 322.765 ;
        RECT 693.210 322.595 693.380 322.765 ;
        RECT 693.570 322.595 693.740 322.765 ;
        RECT 694.820 322.595 694.990 322.765 ;
        RECT 695.180 322.595 695.350 322.765 ;
        RECT 851.745 323.300 851.915 323.470 ;
        RECT 851.745 322.940 851.915 323.110 ;
        RECT 853.910 322.945 854.080 323.115 ;
        RECT 851.745 322.580 851.915 322.750 ;
        RECT 658.915 322.115 659.085 322.285 ;
        RECT 659.395 322.115 659.565 322.285 ;
        RECT 659.875 322.115 660.045 322.285 ;
        RECT 663.815 322.075 663.985 322.245 ;
        RECT 664.295 322.075 664.465 322.245 ;
        RECT 664.775 322.075 664.945 322.245 ;
        RECT 668.405 322.105 668.575 322.275 ;
        RECT 668.885 322.105 669.055 322.275 ;
        RECT 669.365 322.105 669.535 322.275 ;
        RECT 672.945 322.085 673.115 322.255 ;
        RECT 673.425 322.085 673.595 322.255 ;
        RECT 673.905 322.085 674.075 322.255 ;
        RECT 676.375 322.095 676.545 322.265 ;
        RECT 676.855 322.095 677.025 322.265 ;
        RECT 677.335 322.095 677.505 322.265 ;
        RECT 677.815 322.095 677.985 322.265 ;
        RECT 678.295 322.095 678.465 322.265 ;
        RECT 678.775 322.095 678.945 322.265 ;
        RECT 679.255 322.095 679.425 322.265 ;
        RECT 679.735 322.095 679.905 322.265 ;
        RECT 682.145 322.095 682.315 322.265 ;
        RECT 682.625 322.095 682.795 322.265 ;
        RECT 683.105 322.095 683.275 322.265 ;
        RECT 683.585 322.095 683.755 322.265 ;
        RECT 684.065 322.095 684.235 322.265 ;
        RECT 684.545 322.095 684.715 322.265 ;
        RECT 685.025 322.095 685.195 322.265 ;
        RECT 687.595 322.095 687.765 322.265 ;
        RECT 688.075 322.095 688.245 322.265 ;
        RECT 688.555 322.095 688.725 322.265 ;
        RECT 689.035 322.095 689.205 322.265 ;
        RECT 689.515 322.095 689.685 322.265 ;
        RECT 689.995 322.095 690.165 322.265 ;
        RECT 690.475 322.095 690.645 322.265 ;
        RECT 692.905 322.115 693.075 322.285 ;
        RECT 693.385 322.115 693.555 322.285 ;
        RECT 693.865 322.115 694.035 322.285 ;
        RECT 694.345 322.115 694.515 322.285 ;
        RECT 694.825 322.115 694.995 322.285 ;
        RECT 695.305 322.115 695.475 322.285 ;
        RECT 695.785 322.115 695.955 322.285 ;
        RECT 851.745 322.220 851.915 322.390 ;
        RECT 851.745 321.860 851.915 322.030 ;
        RECT 851.745 321.500 851.915 321.670 ;
        RECT 853.910 321.475 854.080 321.645 ;
        RECT 851.745 321.140 851.915 321.310 ;
        RECT 851.745 320.780 851.915 320.950 ;
        RECT 851.745 320.420 851.915 320.590 ;
        RECT 874.510 320.505 874.680 320.675 ;
        RECT 851.745 320.060 851.915 320.230 ;
        RECT 853.910 320.005 854.080 320.175 ;
        RECT 851.745 319.700 851.915 319.870 ;
        RECT 851.745 319.340 851.915 319.510 ;
        RECT 876.870 319.825 877.040 319.995 ;
        RECT 876.870 319.465 877.040 319.635 ;
        RECT 851.745 318.980 851.915 319.150 ;
        RECT 874.510 319.035 874.680 319.205 ;
        RECT 876.870 319.105 877.040 319.275 ;
        RECT 851.745 318.620 851.915 318.790 ;
        RECT 851.745 318.260 851.915 318.430 ;
        RECT 853.910 318.535 854.080 318.705 ;
        RECT 876.870 318.745 877.040 318.915 ;
        RECT 851.745 317.900 851.915 318.070 ;
        RECT 876.870 318.385 877.040 318.555 ;
        RECT 876.870 318.025 877.040 318.195 ;
        RECT 663.885 316.715 664.055 316.885 ;
        RECT 664.415 316.715 664.585 316.885 ;
        RECT 668.905 316.725 669.075 316.895 ;
        RECT 669.265 316.725 669.435 316.895 ;
        RECT 669.625 316.725 669.795 316.895 ;
        RECT 674.345 316.735 674.515 316.905 ;
        RECT 674.705 316.735 674.875 316.905 ;
        RECT 675.065 316.735 675.235 316.905 ;
        RECT 678.080 316.735 678.250 316.905 ;
        RECT 678.440 316.735 678.610 316.905 ;
        RECT 678.800 316.735 678.970 316.905 ;
        RECT 680.050 316.735 680.220 316.905 ;
        RECT 680.410 316.735 680.580 316.905 ;
        RECT 851.745 317.540 851.915 317.710 ;
        RECT 874.510 317.565 874.680 317.735 ;
        RECT 876.870 317.665 877.040 317.835 ;
        RECT 685.015 316.735 685.185 316.905 ;
        RECT 685.375 316.735 685.545 316.905 ;
        RECT 685.735 316.735 685.905 316.905 ;
        RECT 689.755 316.715 689.925 316.885 ;
        RECT 690.115 316.715 690.285 316.885 ;
        RECT 690.475 316.715 690.645 316.885 ;
        RECT 690.835 316.715 691.005 316.885 ;
        RECT 694.155 316.715 694.325 316.885 ;
        RECT 694.515 316.715 694.685 316.885 ;
        RECT 694.875 316.715 695.045 316.885 ;
        RECT 695.235 316.715 695.405 316.885 ;
        RECT 851.745 317.180 851.915 317.350 ;
        RECT 851.745 316.820 851.915 316.990 ;
        RECT 853.910 317.065 854.080 317.235 ;
        RECT 876.870 317.305 877.040 317.475 ;
        RECT 876.870 316.945 877.040 317.115 ;
        RECT 661.555 316.235 661.725 316.405 ;
        RECT 662.035 316.235 662.205 316.405 ;
        RECT 662.515 316.235 662.685 316.405 ;
        RECT 662.995 316.235 663.165 316.405 ;
        RECT 663.475 316.235 663.645 316.405 ;
        RECT 663.955 316.235 664.125 316.405 ;
        RECT 664.435 316.235 664.605 316.405 ;
        RECT 664.915 316.235 665.085 316.405 ;
        RECT 667.375 316.245 667.545 316.415 ;
        RECT 667.855 316.245 668.025 316.415 ;
        RECT 668.335 316.245 668.505 316.415 ;
        RECT 668.815 316.245 668.985 316.415 ;
        RECT 669.295 316.245 669.465 316.415 ;
        RECT 669.775 316.245 669.945 316.415 ;
        RECT 670.255 316.245 670.425 316.415 ;
        RECT 672.815 316.255 672.985 316.425 ;
        RECT 673.295 316.255 673.465 316.425 ;
        RECT 673.775 316.255 673.945 316.425 ;
        RECT 674.255 316.255 674.425 316.425 ;
        RECT 674.735 316.255 674.905 316.425 ;
        RECT 675.215 316.255 675.385 316.425 ;
        RECT 675.695 316.255 675.865 316.425 ;
        RECT 678.135 316.255 678.305 316.425 ;
        RECT 678.615 316.255 678.785 316.425 ;
        RECT 679.095 316.255 679.265 316.425 ;
        RECT 679.575 316.255 679.745 316.425 ;
        RECT 680.055 316.255 680.225 316.425 ;
        RECT 680.535 316.255 680.705 316.425 ;
        RECT 681.015 316.255 681.185 316.425 ;
        RECT 683.485 316.255 683.655 316.425 ;
        RECT 683.965 316.255 684.135 316.425 ;
        RECT 684.445 316.255 684.615 316.425 ;
        RECT 684.925 316.255 685.095 316.425 ;
        RECT 685.405 316.255 685.575 316.425 ;
        RECT 685.885 316.255 686.055 316.425 ;
        RECT 686.365 316.255 686.535 316.425 ;
        RECT 689.305 316.235 689.475 316.405 ;
        RECT 689.785 316.235 689.955 316.405 ;
        RECT 690.265 316.235 690.435 316.405 ;
        RECT 690.745 316.235 690.915 316.405 ;
        RECT 691.225 316.235 691.395 316.405 ;
        RECT 693.705 316.235 693.875 316.405 ;
        RECT 694.185 316.235 694.355 316.405 ;
        RECT 694.665 316.235 694.835 316.405 ;
        RECT 695.145 316.235 695.315 316.405 ;
        RECT 695.625 316.235 695.795 316.405 ;
        RECT 876.870 316.585 877.040 316.755 ;
        RECT 874.510 316.095 874.680 316.265 ;
        RECT 876.870 316.225 877.040 316.395 ;
        RECT 853.910 315.595 854.080 315.765 ;
        RECT 876.870 315.865 877.040 316.035 ;
        RECT 876.870 315.505 877.040 315.675 ;
        RECT 876.870 315.145 877.040 315.315 ;
        RECT 874.510 314.625 874.680 314.795 ;
        RECT 853.910 314.125 854.080 314.295 ;
        RECT 635.230 309.385 635.400 309.555 ;
        RECT 635.590 309.385 635.760 309.555 ;
        RECT 639.420 309.475 639.590 309.645 ;
        RECT 639.780 309.475 639.950 309.645 ;
        RECT 643.520 309.455 643.690 309.625 ;
        RECT 643.880 309.455 644.050 309.625 ;
        RECT 596.010 308.935 596.180 309.105 ;
        RECT 596.370 308.935 596.540 309.105 ;
        RECT 595.375 308.455 595.545 308.625 ;
        RECT 595.855 308.455 596.025 308.625 ;
        RECT 596.335 308.455 596.505 308.625 ;
        RECT 596.480 307.735 596.650 307.905 ;
        RECT 596.840 307.735 597.010 307.905 ;
        RECT 605.345 304.725 605.875 308.135 ;
        RECT 635.265 308.905 635.435 309.075 ;
        RECT 635.745 308.905 635.915 309.075 ;
        RECT 636.225 308.905 636.395 309.075 ;
        RECT 639.455 308.995 639.625 309.165 ;
        RECT 639.935 308.995 640.105 309.165 ;
        RECT 640.415 308.995 640.585 309.165 ;
        RECT 643.555 308.975 643.725 309.145 ;
        RECT 644.035 308.975 644.205 309.145 ;
        RECT 644.515 308.975 644.685 309.145 ;
        RECT 625.750 308.065 625.920 308.235 ;
        RECT 625.750 307.705 625.920 307.875 ;
        RECT 625.750 307.345 625.920 307.515 ;
        RECT 625.750 306.985 625.920 307.155 ;
        RECT 625.750 306.625 625.920 306.795 ;
        RECT 614.870 306.255 615.040 306.425 ;
        RECT 616.450 306.255 616.620 306.425 ;
        RECT 625.750 306.265 625.920 306.435 ;
        RECT 625.750 305.905 625.920 306.075 ;
        RECT 625.750 305.545 625.920 305.715 ;
        RECT 625.750 305.185 625.920 305.355 ;
        RECT 640.220 305.365 640.390 305.535 ;
        RECT 644.270 305.415 644.440 305.585 ;
        RECT 614.870 304.785 615.040 304.955 ;
        RECT 616.450 304.785 616.620 304.955 ;
        RECT 797.070 304.425 797.240 304.595 ;
        RECT 797.430 304.425 797.600 304.595 ;
        RECT 797.790 304.425 797.960 304.595 ;
        RECT 798.710 304.425 798.880 304.595 ;
        RECT 799.070 304.425 799.240 304.595 ;
        RECT 803.670 304.425 803.840 304.595 ;
        RECT 804.030 304.425 804.200 304.595 ;
        RECT 804.390 304.425 804.560 304.595 ;
        RECT 807.640 304.425 807.810 304.595 ;
        RECT 808.000 304.425 808.170 304.595 ;
        RECT 808.360 304.425 808.530 304.595 ;
        RECT 810.245 304.425 810.415 304.595 ;
        RECT 810.605 304.425 810.775 304.595 ;
        RECT 810.965 304.425 811.135 304.595 ;
        RECT 814.830 304.425 815.000 304.595 ;
        RECT 815.190 304.425 815.360 304.595 ;
        RECT 815.550 304.425 815.720 304.595 ;
        RECT 816.470 304.425 816.640 304.595 ;
        RECT 816.830 304.425 817.000 304.595 ;
        RECT 821.430 304.425 821.600 304.595 ;
        RECT 821.790 304.425 821.960 304.595 ;
        RECT 822.150 304.425 822.320 304.595 ;
        RECT 825.400 304.425 825.570 304.595 ;
        RECT 825.760 304.425 825.930 304.595 ;
        RECT 826.120 304.425 826.290 304.595 ;
        RECT 828.005 304.425 828.175 304.595 ;
        RECT 828.365 304.425 828.535 304.595 ;
        RECT 828.725 304.425 828.895 304.595 ;
        RECT 831.900 304.395 832.070 304.565 ;
        RECT 832.260 304.395 832.430 304.565 ;
        RECT 835.540 304.455 835.710 304.625 ;
        RECT 835.900 304.455 836.070 304.625 ;
        RECT 836.760 304.455 836.930 304.625 ;
        RECT 837.120 304.455 837.290 304.625 ;
        RECT 837.480 304.455 837.650 304.625 ;
        RECT 837.840 304.455 838.010 304.625 ;
        RECT 838.200 304.455 838.370 304.625 ;
        RECT 838.560 304.455 838.730 304.625 ;
        RECT 838.920 304.455 839.090 304.625 ;
        RECT 840.000 304.455 840.170 304.625 ;
        RECT 840.360 304.455 840.530 304.625 ;
        RECT 842.810 304.455 842.980 304.625 ;
        RECT 843.170 304.455 843.340 304.625 ;
        RECT 796.635 303.945 796.805 304.115 ;
        RECT 797.115 303.945 797.285 304.115 ;
        RECT 797.595 303.945 797.765 304.115 ;
        RECT 798.075 303.945 798.245 304.115 ;
        RECT 798.555 303.945 798.725 304.115 ;
        RECT 799.035 303.945 799.205 304.115 ;
        RECT 799.515 303.945 799.685 304.115 ;
        RECT 799.995 303.945 800.165 304.115 ;
        RECT 800.475 303.945 800.645 304.115 ;
        RECT 800.955 303.945 801.125 304.115 ;
        RECT 801.435 303.945 801.605 304.115 ;
        RECT 801.915 303.945 802.085 304.115 ;
        RECT 802.395 303.945 802.565 304.115 ;
        RECT 802.875 303.945 803.045 304.115 ;
        RECT 803.355 303.945 803.525 304.115 ;
        RECT 803.835 303.945 804.005 304.115 ;
        RECT 804.315 303.945 804.485 304.115 ;
        RECT 804.795 303.945 804.965 304.115 ;
        RECT 805.275 303.945 805.445 304.115 ;
        RECT 805.755 303.945 805.925 304.115 ;
        RECT 806.235 303.945 806.405 304.115 ;
        RECT 806.715 303.945 806.885 304.115 ;
        RECT 807.195 303.945 807.365 304.115 ;
        RECT 807.675 303.945 807.845 304.115 ;
        RECT 808.155 303.945 808.325 304.115 ;
        RECT 808.635 303.945 808.805 304.115 ;
        RECT 809.115 303.945 809.285 304.115 ;
        RECT 809.595 303.945 809.765 304.115 ;
        RECT 810.075 303.945 810.245 304.115 ;
        RECT 810.555 303.945 810.725 304.115 ;
        RECT 811.035 303.945 811.205 304.115 ;
        RECT 811.515 303.945 811.685 304.115 ;
        RECT 814.395 303.945 814.565 304.115 ;
        RECT 814.875 303.945 815.045 304.115 ;
        RECT 815.355 303.945 815.525 304.115 ;
        RECT 815.835 303.945 816.005 304.115 ;
        RECT 816.315 303.945 816.485 304.115 ;
        RECT 816.795 303.945 816.965 304.115 ;
        RECT 817.275 303.945 817.445 304.115 ;
        RECT 817.755 303.945 817.925 304.115 ;
        RECT 818.235 303.945 818.405 304.115 ;
        RECT 818.715 303.945 818.885 304.115 ;
        RECT 819.195 303.945 819.365 304.115 ;
        RECT 819.675 303.945 819.845 304.115 ;
        RECT 820.155 303.945 820.325 304.115 ;
        RECT 820.635 303.945 820.805 304.115 ;
        RECT 821.115 303.945 821.285 304.115 ;
        RECT 821.595 303.945 821.765 304.115 ;
        RECT 822.075 303.945 822.245 304.115 ;
        RECT 822.555 303.945 822.725 304.115 ;
        RECT 823.035 303.945 823.205 304.115 ;
        RECT 823.515 303.945 823.685 304.115 ;
        RECT 823.995 303.945 824.165 304.115 ;
        RECT 824.475 303.945 824.645 304.115 ;
        RECT 824.955 303.945 825.125 304.115 ;
        RECT 825.435 303.945 825.605 304.115 ;
        RECT 825.915 303.945 826.085 304.115 ;
        RECT 826.395 303.945 826.565 304.115 ;
        RECT 826.875 303.945 827.045 304.115 ;
        RECT 827.355 303.945 827.525 304.115 ;
        RECT 827.835 303.945 828.005 304.115 ;
        RECT 828.315 303.945 828.485 304.115 ;
        RECT 828.795 303.945 828.965 304.115 ;
        RECT 829.275 303.945 829.445 304.115 ;
        RECT 831.935 303.915 832.105 304.085 ;
        RECT 832.415 303.915 832.585 304.085 ;
        RECT 832.895 303.915 833.065 304.085 ;
        RECT 835.575 303.975 835.745 304.145 ;
        RECT 836.055 303.975 836.225 304.145 ;
        RECT 836.535 303.975 836.705 304.145 ;
        RECT 837.015 303.975 837.185 304.145 ;
        RECT 837.495 303.975 837.665 304.145 ;
        RECT 837.975 303.975 838.145 304.145 ;
        RECT 838.455 303.975 838.625 304.145 ;
        RECT 838.935 303.975 839.105 304.145 ;
        RECT 839.415 303.975 839.585 304.145 ;
        RECT 839.895 303.975 840.065 304.145 ;
        RECT 840.375 303.975 840.545 304.145 ;
        RECT 842.845 303.975 843.015 304.145 ;
        RECT 843.325 303.975 843.495 304.145 ;
        RECT 843.805 303.975 843.975 304.145 ;
        RECT 680.650 295.365 680.820 295.535 ;
        RECT 681.010 295.365 681.180 295.535 ;
        RECT 681.370 295.365 681.540 295.535 ;
        RECT 682.290 295.365 682.460 295.535 ;
        RECT 682.650 295.365 682.820 295.535 ;
        RECT 687.250 295.365 687.420 295.535 ;
        RECT 687.610 295.365 687.780 295.535 ;
        RECT 687.970 295.365 688.140 295.535 ;
        RECT 691.220 295.365 691.390 295.535 ;
        RECT 691.580 295.365 691.750 295.535 ;
        RECT 691.940 295.365 692.110 295.535 ;
        RECT 693.825 295.365 693.995 295.535 ;
        RECT 694.185 295.365 694.355 295.535 ;
        RECT 694.545 295.365 694.715 295.535 ;
        RECT 698.140 295.325 698.310 295.495 ;
        RECT 698.500 295.325 698.670 295.495 ;
        RECT 698.860 295.325 699.030 295.495 ;
        RECT 699.780 295.325 699.950 295.495 ;
        RECT 700.140 295.325 700.310 295.495 ;
        RECT 704.740 295.325 704.910 295.495 ;
        RECT 705.100 295.325 705.270 295.495 ;
        RECT 705.460 295.325 705.630 295.495 ;
        RECT 708.710 295.325 708.880 295.495 ;
        RECT 709.070 295.325 709.240 295.495 ;
        RECT 709.430 295.325 709.600 295.495 ;
        RECT 711.315 295.325 711.485 295.495 ;
        RECT 711.675 295.325 711.845 295.495 ;
        RECT 712.035 295.325 712.205 295.495 ;
        RECT 715.750 295.385 715.920 295.555 ;
        RECT 716.110 295.385 716.280 295.555 ;
        RECT 716.470 295.385 716.640 295.555 ;
        RECT 717.390 295.385 717.560 295.555 ;
        RECT 717.750 295.385 717.920 295.555 ;
        RECT 722.350 295.385 722.520 295.555 ;
        RECT 722.710 295.385 722.880 295.555 ;
        RECT 723.070 295.385 723.240 295.555 ;
        RECT 726.320 295.385 726.490 295.555 ;
        RECT 726.680 295.385 726.850 295.555 ;
        RECT 727.040 295.385 727.210 295.555 ;
        RECT 728.925 295.385 729.095 295.555 ;
        RECT 729.285 295.385 729.455 295.555 ;
        RECT 729.645 295.385 729.815 295.555 ;
        RECT 733.450 295.335 733.620 295.505 ;
        RECT 733.810 295.335 733.980 295.505 ;
        RECT 734.170 295.335 734.340 295.505 ;
        RECT 735.090 295.335 735.260 295.505 ;
        RECT 735.450 295.335 735.620 295.505 ;
        RECT 740.050 295.335 740.220 295.505 ;
        RECT 740.410 295.335 740.580 295.505 ;
        RECT 740.770 295.335 740.940 295.505 ;
        RECT 744.020 295.335 744.190 295.505 ;
        RECT 744.380 295.335 744.550 295.505 ;
        RECT 744.740 295.335 744.910 295.505 ;
        RECT 746.625 295.335 746.795 295.505 ;
        RECT 746.985 295.335 747.155 295.505 ;
        RECT 747.345 295.335 747.515 295.505 ;
        RECT 751.190 295.325 751.360 295.495 ;
        RECT 751.550 295.325 751.720 295.495 ;
        RECT 751.910 295.325 752.080 295.495 ;
        RECT 752.830 295.325 753.000 295.495 ;
        RECT 753.190 295.325 753.360 295.495 ;
        RECT 757.790 295.325 757.960 295.495 ;
        RECT 758.150 295.325 758.320 295.495 ;
        RECT 758.510 295.325 758.680 295.495 ;
        RECT 761.760 295.325 761.930 295.495 ;
        RECT 762.120 295.325 762.290 295.495 ;
        RECT 762.480 295.325 762.650 295.495 ;
        RECT 764.365 295.325 764.535 295.495 ;
        RECT 764.725 295.325 764.895 295.495 ;
        RECT 765.085 295.325 765.255 295.495 ;
        RECT 680.215 294.885 680.385 295.055 ;
        RECT 680.695 294.885 680.865 295.055 ;
        RECT 681.175 294.885 681.345 295.055 ;
        RECT 681.655 294.885 681.825 295.055 ;
        RECT 682.135 294.885 682.305 295.055 ;
        RECT 682.615 294.885 682.785 295.055 ;
        RECT 683.095 294.885 683.265 295.055 ;
        RECT 683.575 294.885 683.745 295.055 ;
        RECT 684.055 294.885 684.225 295.055 ;
        RECT 684.535 294.885 684.705 295.055 ;
        RECT 685.015 294.885 685.185 295.055 ;
        RECT 685.495 294.885 685.665 295.055 ;
        RECT 685.975 294.885 686.145 295.055 ;
        RECT 686.455 294.885 686.625 295.055 ;
        RECT 686.935 294.885 687.105 295.055 ;
        RECT 687.415 294.885 687.585 295.055 ;
        RECT 687.895 294.885 688.065 295.055 ;
        RECT 688.375 294.885 688.545 295.055 ;
        RECT 688.855 294.885 689.025 295.055 ;
        RECT 689.335 294.885 689.505 295.055 ;
        RECT 689.815 294.885 689.985 295.055 ;
        RECT 690.295 294.885 690.465 295.055 ;
        RECT 690.775 294.885 690.945 295.055 ;
        RECT 691.255 294.885 691.425 295.055 ;
        RECT 691.735 294.885 691.905 295.055 ;
        RECT 692.215 294.885 692.385 295.055 ;
        RECT 692.695 294.885 692.865 295.055 ;
        RECT 693.175 294.885 693.345 295.055 ;
        RECT 693.655 294.885 693.825 295.055 ;
        RECT 694.135 294.885 694.305 295.055 ;
        RECT 694.615 294.885 694.785 295.055 ;
        RECT 695.095 294.885 695.265 295.055 ;
        RECT 697.705 294.845 697.875 295.015 ;
        RECT 698.185 294.845 698.355 295.015 ;
        RECT 698.665 294.845 698.835 295.015 ;
        RECT 699.145 294.845 699.315 295.015 ;
        RECT 699.625 294.845 699.795 295.015 ;
        RECT 700.105 294.845 700.275 295.015 ;
        RECT 700.585 294.845 700.755 295.015 ;
        RECT 701.065 294.845 701.235 295.015 ;
        RECT 701.545 294.845 701.715 295.015 ;
        RECT 702.025 294.845 702.195 295.015 ;
        RECT 702.505 294.845 702.675 295.015 ;
        RECT 702.985 294.845 703.155 295.015 ;
        RECT 703.465 294.845 703.635 295.015 ;
        RECT 703.945 294.845 704.115 295.015 ;
        RECT 704.425 294.845 704.595 295.015 ;
        RECT 704.905 294.845 705.075 295.015 ;
        RECT 705.385 294.845 705.555 295.015 ;
        RECT 705.865 294.845 706.035 295.015 ;
        RECT 706.345 294.845 706.515 295.015 ;
        RECT 706.825 294.845 706.995 295.015 ;
        RECT 707.305 294.845 707.475 295.015 ;
        RECT 707.785 294.845 707.955 295.015 ;
        RECT 708.265 294.845 708.435 295.015 ;
        RECT 708.745 294.845 708.915 295.015 ;
        RECT 709.225 294.845 709.395 295.015 ;
        RECT 709.705 294.845 709.875 295.015 ;
        RECT 710.185 294.845 710.355 295.015 ;
        RECT 710.665 294.845 710.835 295.015 ;
        RECT 711.145 294.845 711.315 295.015 ;
        RECT 711.625 294.845 711.795 295.015 ;
        RECT 712.105 294.845 712.275 295.015 ;
        RECT 712.585 294.845 712.755 295.015 ;
        RECT 715.315 294.905 715.485 295.075 ;
        RECT 715.795 294.905 715.965 295.075 ;
        RECT 716.275 294.905 716.445 295.075 ;
        RECT 716.755 294.905 716.925 295.075 ;
        RECT 717.235 294.905 717.405 295.075 ;
        RECT 717.715 294.905 717.885 295.075 ;
        RECT 718.195 294.905 718.365 295.075 ;
        RECT 718.675 294.905 718.845 295.075 ;
        RECT 719.155 294.905 719.325 295.075 ;
        RECT 719.635 294.905 719.805 295.075 ;
        RECT 720.115 294.905 720.285 295.075 ;
        RECT 720.595 294.905 720.765 295.075 ;
        RECT 721.075 294.905 721.245 295.075 ;
        RECT 721.555 294.905 721.725 295.075 ;
        RECT 722.035 294.905 722.205 295.075 ;
        RECT 722.515 294.905 722.685 295.075 ;
        RECT 722.995 294.905 723.165 295.075 ;
        RECT 723.475 294.905 723.645 295.075 ;
        RECT 723.955 294.905 724.125 295.075 ;
        RECT 724.435 294.905 724.605 295.075 ;
        RECT 724.915 294.905 725.085 295.075 ;
        RECT 725.395 294.905 725.565 295.075 ;
        RECT 725.875 294.905 726.045 295.075 ;
        RECT 726.355 294.905 726.525 295.075 ;
        RECT 726.835 294.905 727.005 295.075 ;
        RECT 727.315 294.905 727.485 295.075 ;
        RECT 727.795 294.905 727.965 295.075 ;
        RECT 728.275 294.905 728.445 295.075 ;
        RECT 728.755 294.905 728.925 295.075 ;
        RECT 729.235 294.905 729.405 295.075 ;
        RECT 729.715 294.905 729.885 295.075 ;
        RECT 730.195 294.905 730.365 295.075 ;
        RECT 733.015 294.855 733.185 295.025 ;
        RECT 733.495 294.855 733.665 295.025 ;
        RECT 733.975 294.855 734.145 295.025 ;
        RECT 734.455 294.855 734.625 295.025 ;
        RECT 734.935 294.855 735.105 295.025 ;
        RECT 735.415 294.855 735.585 295.025 ;
        RECT 735.895 294.855 736.065 295.025 ;
        RECT 736.375 294.855 736.545 295.025 ;
        RECT 736.855 294.855 737.025 295.025 ;
        RECT 737.335 294.855 737.505 295.025 ;
        RECT 737.815 294.855 737.985 295.025 ;
        RECT 738.295 294.855 738.465 295.025 ;
        RECT 738.775 294.855 738.945 295.025 ;
        RECT 739.255 294.855 739.425 295.025 ;
        RECT 739.735 294.855 739.905 295.025 ;
        RECT 740.215 294.855 740.385 295.025 ;
        RECT 740.695 294.855 740.865 295.025 ;
        RECT 741.175 294.855 741.345 295.025 ;
        RECT 741.655 294.855 741.825 295.025 ;
        RECT 742.135 294.855 742.305 295.025 ;
        RECT 742.615 294.855 742.785 295.025 ;
        RECT 743.095 294.855 743.265 295.025 ;
        RECT 743.575 294.855 743.745 295.025 ;
        RECT 744.055 294.855 744.225 295.025 ;
        RECT 744.535 294.855 744.705 295.025 ;
        RECT 745.015 294.855 745.185 295.025 ;
        RECT 745.495 294.855 745.665 295.025 ;
        RECT 745.975 294.855 746.145 295.025 ;
        RECT 746.455 294.855 746.625 295.025 ;
        RECT 746.935 294.855 747.105 295.025 ;
        RECT 747.415 294.855 747.585 295.025 ;
        RECT 747.895 294.855 748.065 295.025 ;
        RECT 750.755 294.845 750.925 295.015 ;
        RECT 751.235 294.845 751.405 295.015 ;
        RECT 751.715 294.845 751.885 295.015 ;
        RECT 752.195 294.845 752.365 295.015 ;
        RECT 752.675 294.845 752.845 295.015 ;
        RECT 753.155 294.845 753.325 295.015 ;
        RECT 753.635 294.845 753.805 295.015 ;
        RECT 754.115 294.845 754.285 295.015 ;
        RECT 754.595 294.845 754.765 295.015 ;
        RECT 755.075 294.845 755.245 295.015 ;
        RECT 755.555 294.845 755.725 295.015 ;
        RECT 756.035 294.845 756.205 295.015 ;
        RECT 756.515 294.845 756.685 295.015 ;
        RECT 756.995 294.845 757.165 295.015 ;
        RECT 757.475 294.845 757.645 295.015 ;
        RECT 757.955 294.845 758.125 295.015 ;
        RECT 758.435 294.845 758.605 295.015 ;
        RECT 758.915 294.845 759.085 295.015 ;
        RECT 759.395 294.845 759.565 295.015 ;
        RECT 759.875 294.845 760.045 295.015 ;
        RECT 760.355 294.845 760.525 295.015 ;
        RECT 760.835 294.845 761.005 295.015 ;
        RECT 761.315 294.845 761.485 295.015 ;
        RECT 761.795 294.845 761.965 295.015 ;
        RECT 762.275 294.845 762.445 295.015 ;
        RECT 762.755 294.845 762.925 295.015 ;
        RECT 763.235 294.845 763.405 295.015 ;
        RECT 763.715 294.845 763.885 295.015 ;
        RECT 764.195 294.845 764.365 295.015 ;
        RECT 764.675 294.845 764.845 295.015 ;
        RECT 765.155 294.845 765.325 295.015 ;
        RECT 765.635 294.845 765.805 295.015 ;
        RECT 857.485 294.685 857.655 294.855 ;
        RECT 857.845 294.685 858.015 294.855 ;
        RECT 858.205 294.685 858.375 294.855 ;
        RECT 855.955 294.205 856.125 294.375 ;
        RECT 856.435 294.205 856.605 294.375 ;
        RECT 856.915 294.205 857.085 294.375 ;
        RECT 857.395 294.205 857.565 294.375 ;
        RECT 857.875 294.205 858.045 294.375 ;
        RECT 858.355 294.205 858.525 294.375 ;
        RECT 858.835 294.205 859.005 294.375 ;
        RECT 841.075 292.705 841.245 292.875 ;
        RECT 841.435 292.705 841.605 292.875 ;
        RECT 841.795 292.705 841.965 292.875 ;
        RECT 839.545 292.225 839.715 292.395 ;
        RECT 840.025 292.225 840.195 292.395 ;
        RECT 840.505 292.225 840.675 292.395 ;
        RECT 840.985 292.225 841.155 292.395 ;
        RECT 841.465 292.225 841.635 292.395 ;
        RECT 841.945 292.225 842.115 292.395 ;
        RECT 842.425 292.225 842.595 292.395 ;
        RECT 635.180 290.205 635.350 290.375 ;
        RECT 635.540 290.205 635.710 290.375 ;
        RECT 639.370 290.295 639.540 290.465 ;
        RECT 639.730 290.295 639.900 290.465 ;
        RECT 643.470 290.275 643.640 290.445 ;
        RECT 643.830 290.275 644.000 290.445 ;
        RECT 595.960 289.755 596.130 289.925 ;
        RECT 596.320 289.755 596.490 289.925 ;
        RECT 595.325 289.275 595.495 289.445 ;
        RECT 595.805 289.275 595.975 289.445 ;
        RECT 596.285 289.275 596.455 289.445 ;
        RECT 596.430 288.555 596.600 288.725 ;
        RECT 596.790 288.555 596.960 288.725 ;
        RECT 118.335 287.230 118.505 287.400 ;
        RECT 118.695 287.230 118.865 287.400 ;
        RECT 121.805 287.230 121.975 287.400 ;
        RECT 122.165 287.230 122.335 287.400 ;
        RECT 125.275 287.230 125.445 287.400 ;
        RECT 125.635 287.230 125.805 287.400 ;
        RECT 128.745 287.230 128.915 287.400 ;
        RECT 129.105 287.230 129.275 287.400 ;
        RECT 132.215 287.230 132.385 287.400 ;
        RECT 132.575 287.230 132.745 287.400 ;
        RECT 135.685 287.230 135.855 287.400 ;
        RECT 136.045 287.230 136.215 287.400 ;
        RECT 139.155 287.230 139.325 287.400 ;
        RECT 139.515 287.230 139.685 287.400 ;
        RECT 142.625 287.230 142.795 287.400 ;
        RECT 142.985 287.230 143.155 287.400 ;
        RECT 146.095 287.230 146.265 287.400 ;
        RECT 146.455 287.230 146.625 287.400 ;
        RECT 149.565 287.230 149.735 287.400 ;
        RECT 149.925 287.230 150.095 287.400 ;
        RECT 605.295 285.545 605.825 288.955 ;
        RECT 635.215 289.725 635.385 289.895 ;
        RECT 635.695 289.725 635.865 289.895 ;
        RECT 636.175 289.725 636.345 289.895 ;
        RECT 639.405 289.815 639.575 289.985 ;
        RECT 639.885 289.815 640.055 289.985 ;
        RECT 640.365 289.815 640.535 289.985 ;
        RECT 643.505 289.795 643.675 289.965 ;
        RECT 643.985 289.795 644.155 289.965 ;
        RECT 644.465 289.795 644.635 289.965 ;
        RECT 845.190 291.055 845.360 291.225 ;
        RECT 845.550 291.055 845.720 291.225 ;
        RECT 845.910 291.055 846.080 291.225 ;
        RECT 847.160 291.055 847.330 291.225 ;
        RECT 847.520 291.055 847.690 291.225 ;
        RECT 861.280 290.785 861.450 290.955 ;
        RECT 861.640 290.785 861.810 290.955 ;
        RECT 862.000 290.785 862.170 290.955 ;
        RECT 863.250 290.785 863.420 290.955 ;
        RECT 863.610 290.785 863.780 290.955 ;
        RECT 845.245 290.575 845.415 290.745 ;
        RECT 845.725 290.575 845.895 290.745 ;
        RECT 846.205 290.575 846.375 290.745 ;
        RECT 846.685 290.575 846.855 290.745 ;
        RECT 847.165 290.575 847.335 290.745 ;
        RECT 847.645 290.575 847.815 290.745 ;
        RECT 848.125 290.575 848.295 290.745 ;
        RECT 861.335 290.305 861.505 290.475 ;
        RECT 861.815 290.305 861.985 290.475 ;
        RECT 862.295 290.305 862.465 290.475 ;
        RECT 862.775 290.305 862.945 290.475 ;
        RECT 863.255 290.305 863.425 290.475 ;
        RECT 863.735 290.305 863.905 290.475 ;
        RECT 864.215 290.305 864.385 290.475 ;
        RECT 820.625 289.695 820.795 289.865 ;
        RECT 820.985 289.695 821.155 289.865 ;
        RECT 821.345 289.695 821.515 289.865 ;
        RECT 819.095 289.215 819.265 289.385 ;
        RECT 819.575 289.215 819.745 289.385 ;
        RECT 820.055 289.215 820.225 289.385 ;
        RECT 820.535 289.215 820.705 289.385 ;
        RECT 821.015 289.215 821.185 289.385 ;
        RECT 821.495 289.215 821.665 289.385 ;
        RECT 821.975 289.215 822.145 289.385 ;
        RECT 857.525 289.155 857.695 289.325 ;
        RECT 857.885 289.155 858.055 289.325 ;
        RECT 858.245 289.155 858.415 289.325 ;
        RECT 625.700 288.885 625.870 289.055 ;
        RECT 625.700 288.525 625.870 288.695 ;
        RECT 855.995 288.675 856.165 288.845 ;
        RECT 856.475 288.675 856.645 288.845 ;
        RECT 856.955 288.675 857.125 288.845 ;
        RECT 857.435 288.675 857.605 288.845 ;
        RECT 857.915 288.675 858.085 288.845 ;
        RECT 858.395 288.675 858.565 288.845 ;
        RECT 858.875 288.675 859.045 288.845 ;
        RECT 625.700 288.165 625.870 288.335 ;
        RECT 625.700 287.805 625.870 287.975 ;
        RECT 625.700 287.445 625.870 287.615 ;
        RECT 826.075 287.525 826.245 287.695 ;
        RECT 826.435 287.525 826.605 287.695 ;
        RECT 826.795 287.525 826.965 287.695 ;
        RECT 830.050 287.545 830.220 287.715 ;
        RECT 830.410 287.545 830.580 287.715 ;
        RECT 831.270 287.545 831.440 287.715 ;
        RECT 831.630 287.545 831.800 287.715 ;
        RECT 831.990 287.545 832.160 287.715 ;
        RECT 832.350 287.545 832.520 287.715 ;
        RECT 832.710 287.545 832.880 287.715 ;
        RECT 833.070 287.545 833.240 287.715 ;
        RECT 833.430 287.545 833.600 287.715 ;
        RECT 834.510 287.545 834.680 287.715 ;
        RECT 834.870 287.545 835.040 287.715 ;
        RECT 841.085 287.585 841.255 287.755 ;
        RECT 841.445 287.585 841.615 287.755 ;
        RECT 841.805 287.585 841.975 287.755 ;
        RECT 614.820 287.075 614.990 287.245 ;
        RECT 616.400 287.075 616.570 287.245 ;
        RECT 625.700 287.085 625.870 287.255 ;
        RECT 824.545 287.045 824.715 287.215 ;
        RECT 825.025 287.045 825.195 287.215 ;
        RECT 825.505 287.045 825.675 287.215 ;
        RECT 825.985 287.045 826.155 287.215 ;
        RECT 826.465 287.045 826.635 287.215 ;
        RECT 826.945 287.045 827.115 287.215 ;
        RECT 827.425 287.045 827.595 287.215 ;
        RECT 830.085 287.065 830.255 287.235 ;
        RECT 830.565 287.065 830.735 287.235 ;
        RECT 831.045 287.065 831.215 287.235 ;
        RECT 831.525 287.065 831.695 287.235 ;
        RECT 832.005 287.065 832.175 287.235 ;
        RECT 832.485 287.065 832.655 287.235 ;
        RECT 832.965 287.065 833.135 287.235 ;
        RECT 833.445 287.065 833.615 287.235 ;
        RECT 833.925 287.065 834.095 287.235 ;
        RECT 834.405 287.065 834.575 287.235 ;
        RECT 834.885 287.065 835.055 287.235 ;
        RECT 839.555 287.105 839.725 287.275 ;
        RECT 840.035 287.105 840.205 287.275 ;
        RECT 840.515 287.105 840.685 287.275 ;
        RECT 840.995 287.105 841.165 287.275 ;
        RECT 841.475 287.105 841.645 287.275 ;
        RECT 841.955 287.105 842.125 287.275 ;
        RECT 842.435 287.105 842.605 287.275 ;
        RECT 625.700 286.725 625.870 286.895 ;
        RECT 625.700 286.365 625.870 286.535 ;
        RECT 625.700 286.005 625.870 286.175 ;
        RECT 640.170 286.185 640.340 286.355 ;
        RECT 644.220 286.235 644.390 286.405 ;
        RECT 614.820 285.605 614.990 285.775 ;
        RECT 616.400 285.605 616.570 285.775 ;
        RECT 820.595 284.535 820.765 284.705 ;
        RECT 820.955 284.535 821.125 284.705 ;
        RECT 821.315 284.535 821.485 284.705 ;
        RECT 118.335 283.940 118.505 284.110 ;
        RECT 118.695 283.940 118.865 284.110 ;
        RECT 121.805 283.940 121.975 284.110 ;
        RECT 122.165 283.940 122.335 284.110 ;
        RECT 125.275 283.940 125.445 284.110 ;
        RECT 125.635 283.940 125.805 284.110 ;
        RECT 128.745 283.940 128.915 284.110 ;
        RECT 129.105 283.940 129.275 284.110 ;
        RECT 132.215 283.940 132.385 284.110 ;
        RECT 132.575 283.940 132.745 284.110 ;
        RECT 135.685 283.940 135.855 284.110 ;
        RECT 136.045 283.940 136.215 284.110 ;
        RECT 139.155 283.940 139.325 284.110 ;
        RECT 139.515 283.940 139.685 284.110 ;
        RECT 142.625 283.940 142.795 284.110 ;
        RECT 142.985 283.940 143.155 284.110 ;
        RECT 146.095 283.940 146.265 284.110 ;
        RECT 146.455 283.940 146.625 284.110 ;
        RECT 149.565 283.940 149.735 284.110 ;
        RECT 149.925 283.940 150.095 284.110 ;
        RECT 151.750 283.970 151.920 284.140 ;
        RECT 819.065 284.055 819.235 284.225 ;
        RECT 819.545 284.055 819.715 284.225 ;
        RECT 820.025 284.055 820.195 284.225 ;
        RECT 820.505 284.055 820.675 284.225 ;
        RECT 820.985 284.055 821.155 284.225 ;
        RECT 821.465 284.055 821.635 284.225 ;
        RECT 821.945 284.055 822.115 284.225 ;
        RECT 857.595 283.755 857.765 283.925 ;
        RECT 857.955 283.755 858.125 283.925 ;
        RECT 858.315 283.755 858.485 283.925 ;
        RECT 856.065 283.275 856.235 283.445 ;
        RECT 856.545 283.275 856.715 283.445 ;
        RECT 857.025 283.275 857.195 283.445 ;
        RECT 857.505 283.275 857.675 283.445 ;
        RECT 857.985 283.275 858.155 283.445 ;
        RECT 858.465 283.275 858.635 283.445 ;
        RECT 858.945 283.275 859.115 283.445 ;
        RECT 861.360 281.735 861.530 281.905 ;
        RECT 861.720 281.735 861.890 281.905 ;
        RECT 862.080 281.735 862.250 281.905 ;
        RECT 863.330 281.735 863.500 281.905 ;
        RECT 863.690 281.735 863.860 281.905 ;
        RECT 861.415 281.255 861.585 281.425 ;
        RECT 861.895 281.255 862.065 281.425 ;
        RECT 862.375 281.255 862.545 281.425 ;
        RECT 862.855 281.255 863.025 281.425 ;
        RECT 863.335 281.255 863.505 281.425 ;
        RECT 863.815 281.255 863.985 281.425 ;
        RECT 864.295 281.255 864.465 281.425 ;
        RECT 118.335 280.650 118.505 280.820 ;
        RECT 118.695 280.650 118.865 280.820 ;
        RECT 121.805 280.650 121.975 280.820 ;
        RECT 122.165 280.650 122.335 280.820 ;
        RECT 125.275 280.650 125.445 280.820 ;
        RECT 125.635 280.650 125.805 280.820 ;
        RECT 128.745 280.650 128.915 280.820 ;
        RECT 129.105 280.650 129.275 280.820 ;
        RECT 132.215 280.650 132.385 280.820 ;
        RECT 132.575 280.650 132.745 280.820 ;
        RECT 135.685 280.650 135.855 280.820 ;
        RECT 136.045 280.650 136.215 280.820 ;
        RECT 139.155 280.650 139.325 280.820 ;
        RECT 139.515 280.650 139.685 280.820 ;
        RECT 142.625 280.650 142.795 280.820 ;
        RECT 142.985 280.650 143.155 280.820 ;
        RECT 146.095 280.650 146.265 280.820 ;
        RECT 146.455 280.650 146.625 280.820 ;
        RECT 149.565 280.650 149.735 280.820 ;
        RECT 149.925 280.650 150.095 280.820 ;
        RECT 799.650 279.845 799.820 280.015 ;
        RECT 800.010 279.845 800.180 280.015 ;
        RECT 144.205 279.535 144.375 279.705 ;
        RECT 144.565 279.535 144.735 279.705 ;
        RECT 144.925 279.535 145.095 279.705 ;
        RECT 145.285 279.535 145.455 279.705 ;
        RECT 145.645 279.535 145.815 279.705 ;
        RECT 146.005 279.535 146.175 279.705 ;
        RECT 146.365 279.535 146.535 279.705 ;
        RECT 146.725 279.535 146.895 279.705 ;
        RECT 147.085 279.535 147.255 279.705 ;
        RECT 122.125 278.995 122.295 279.165 ;
        RECT 122.485 278.995 122.655 279.165 ;
        RECT 122.845 278.995 123.015 279.165 ;
        RECT 123.205 278.995 123.375 279.165 ;
        RECT 123.565 278.995 123.735 279.165 ;
        RECT 123.925 278.995 124.095 279.165 ;
        RECT 124.285 278.995 124.455 279.165 ;
        RECT 124.645 278.995 124.815 279.165 ;
        RECT 125.005 278.995 125.175 279.165 ;
        RECT 679.510 278.625 679.680 278.795 ;
        RECT 679.870 278.625 680.040 278.795 ;
        RECT 680.730 278.625 680.900 278.795 ;
        RECT 681.090 278.625 681.260 278.795 ;
        RECT 681.450 278.625 681.620 278.795 ;
        RECT 681.810 278.625 681.980 278.795 ;
        RECT 682.170 278.625 682.340 278.795 ;
        RECT 682.530 278.625 682.700 278.795 ;
        RECT 682.890 278.625 683.060 278.795 ;
        RECT 683.970 278.625 684.140 278.795 ;
        RECT 684.330 278.625 684.500 278.795 ;
        RECT 696.790 278.635 696.960 278.805 ;
        RECT 697.150 278.635 697.320 278.805 ;
        RECT 698.010 278.635 698.180 278.805 ;
        RECT 698.370 278.635 698.540 278.805 ;
        RECT 698.730 278.635 698.900 278.805 ;
        RECT 699.090 278.635 699.260 278.805 ;
        RECT 699.450 278.635 699.620 278.805 ;
        RECT 699.810 278.635 699.980 278.805 ;
        RECT 700.170 278.635 700.340 278.805 ;
        RECT 701.250 278.635 701.420 278.805 ;
        RECT 701.610 278.635 701.780 278.805 ;
        RECT 714.560 278.635 714.730 278.805 ;
        RECT 714.920 278.635 715.090 278.805 ;
        RECT 715.780 278.635 715.950 278.805 ;
        RECT 716.140 278.635 716.310 278.805 ;
        RECT 716.500 278.635 716.670 278.805 ;
        RECT 716.860 278.635 717.030 278.805 ;
        RECT 717.220 278.635 717.390 278.805 ;
        RECT 717.580 278.635 717.750 278.805 ;
        RECT 717.940 278.635 718.110 278.805 ;
        RECT 719.020 278.635 719.190 278.805 ;
        RECT 719.380 278.635 719.550 278.805 ;
        RECT 731.800 278.635 731.970 278.805 ;
        RECT 732.160 278.635 732.330 278.805 ;
        RECT 733.020 278.635 733.190 278.805 ;
        RECT 733.380 278.635 733.550 278.805 ;
        RECT 733.740 278.635 733.910 278.805 ;
        RECT 734.100 278.635 734.270 278.805 ;
        RECT 734.460 278.635 734.630 278.805 ;
        RECT 734.820 278.635 734.990 278.805 ;
        RECT 735.180 278.635 735.350 278.805 ;
        RECT 736.260 278.635 736.430 278.805 ;
        RECT 736.620 278.635 736.790 278.805 ;
        RECT 749.280 278.645 749.450 278.815 ;
        RECT 749.640 278.645 749.810 278.815 ;
        RECT 750.500 278.645 750.670 278.815 ;
        RECT 750.860 278.645 751.030 278.815 ;
        RECT 751.220 278.645 751.390 278.815 ;
        RECT 751.580 278.645 751.750 278.815 ;
        RECT 751.940 278.645 752.110 278.815 ;
        RECT 752.300 278.645 752.470 278.815 ;
        RECT 752.660 278.645 752.830 278.815 ;
        RECT 799.685 279.365 799.855 279.535 ;
        RECT 800.165 279.365 800.335 279.535 ;
        RECT 800.645 279.365 800.815 279.535 ;
        RECT 819.470 279.505 819.640 279.675 ;
        RECT 819.830 279.505 820.000 279.675 ;
        RECT 820.690 279.505 820.860 279.675 ;
        RECT 821.050 279.505 821.220 279.675 ;
        RECT 821.410 279.505 821.580 279.675 ;
        RECT 821.770 279.505 821.940 279.675 ;
        RECT 822.130 279.505 822.300 279.675 ;
        RECT 822.490 279.505 822.660 279.675 ;
        RECT 822.850 279.505 823.020 279.675 ;
        RECT 823.930 279.505 824.100 279.675 ;
        RECT 824.290 279.505 824.460 279.675 ;
        RECT 829.645 279.415 829.815 279.585 ;
        RECT 830.005 279.415 830.175 279.585 ;
        RECT 830.365 279.415 830.535 279.585 ;
        RECT 833.370 279.415 833.540 279.585 ;
        RECT 833.730 279.415 833.900 279.585 ;
        RECT 834.590 279.415 834.760 279.585 ;
        RECT 834.950 279.415 835.120 279.585 ;
        RECT 835.310 279.415 835.480 279.585 ;
        RECT 835.670 279.415 835.840 279.585 ;
        RECT 836.030 279.415 836.200 279.585 ;
        RECT 836.390 279.415 836.560 279.585 ;
        RECT 836.750 279.415 836.920 279.585 ;
        RECT 837.830 279.415 838.000 279.585 ;
        RECT 838.190 279.415 838.360 279.585 ;
        RECT 842.945 279.415 843.115 279.585 ;
        RECT 843.475 279.415 843.645 279.585 ;
        RECT 846.420 279.415 846.590 279.585 ;
        RECT 846.780 279.415 846.950 279.585 ;
        RECT 847.640 279.415 847.810 279.585 ;
        RECT 848.000 279.415 848.170 279.585 ;
        RECT 848.360 279.415 848.530 279.585 ;
        RECT 848.720 279.415 848.890 279.585 ;
        RECT 849.080 279.415 849.250 279.585 ;
        RECT 849.440 279.415 849.610 279.585 ;
        RECT 849.800 279.415 849.970 279.585 ;
        RECT 850.880 279.415 851.050 279.585 ;
        RECT 851.240 279.415 851.410 279.585 ;
        RECT 819.505 279.025 819.675 279.195 ;
        RECT 819.985 279.025 820.155 279.195 ;
        RECT 820.465 279.025 820.635 279.195 ;
        RECT 820.945 279.025 821.115 279.195 ;
        RECT 821.425 279.025 821.595 279.195 ;
        RECT 821.905 279.025 822.075 279.195 ;
        RECT 822.385 279.025 822.555 279.195 ;
        RECT 822.865 279.025 823.035 279.195 ;
        RECT 823.345 279.025 823.515 279.195 ;
        RECT 823.825 279.025 823.995 279.195 ;
        RECT 824.305 279.025 824.475 279.195 ;
        RECT 828.115 278.935 828.285 279.105 ;
        RECT 828.595 278.935 828.765 279.105 ;
        RECT 829.075 278.935 829.245 279.105 ;
        RECT 829.555 278.935 829.725 279.105 ;
        RECT 830.035 278.935 830.205 279.105 ;
        RECT 830.515 278.935 830.685 279.105 ;
        RECT 830.995 278.935 831.165 279.105 ;
        RECT 833.405 278.935 833.575 279.105 ;
        RECT 833.885 278.935 834.055 279.105 ;
        RECT 834.365 278.935 834.535 279.105 ;
        RECT 834.845 278.935 835.015 279.105 ;
        RECT 835.325 278.935 835.495 279.105 ;
        RECT 835.805 278.935 835.975 279.105 ;
        RECT 836.285 278.935 836.455 279.105 ;
        RECT 836.765 278.935 836.935 279.105 ;
        RECT 837.245 278.935 837.415 279.105 ;
        RECT 837.725 278.935 837.895 279.105 ;
        RECT 838.205 278.935 838.375 279.105 ;
        RECT 840.615 278.935 840.785 279.105 ;
        RECT 841.095 278.935 841.265 279.105 ;
        RECT 841.575 278.935 841.745 279.105 ;
        RECT 842.055 278.935 842.225 279.105 ;
        RECT 842.535 278.935 842.705 279.105 ;
        RECT 843.015 278.935 843.185 279.105 ;
        RECT 843.495 278.935 843.665 279.105 ;
        RECT 843.975 278.935 844.145 279.105 ;
        RECT 846.455 278.935 846.625 279.105 ;
        RECT 846.935 278.935 847.105 279.105 ;
        RECT 847.415 278.935 847.585 279.105 ;
        RECT 847.895 278.935 848.065 279.105 ;
        RECT 848.375 278.935 848.545 279.105 ;
        RECT 848.855 278.935 849.025 279.105 ;
        RECT 849.335 278.935 849.505 279.105 ;
        RECT 849.815 278.935 849.985 279.105 ;
        RECT 850.295 278.935 850.465 279.105 ;
        RECT 850.775 278.935 850.945 279.105 ;
        RECT 851.255 278.935 851.425 279.105 ;
        RECT 753.740 278.645 753.910 278.815 ;
        RECT 754.100 278.645 754.270 278.815 ;
        RECT 679.545 278.145 679.715 278.315 ;
        RECT 680.025 278.145 680.195 278.315 ;
        RECT 680.505 278.145 680.675 278.315 ;
        RECT 680.985 278.145 681.155 278.315 ;
        RECT 681.465 278.145 681.635 278.315 ;
        RECT 681.945 278.145 682.115 278.315 ;
        RECT 682.425 278.145 682.595 278.315 ;
        RECT 682.905 278.145 683.075 278.315 ;
        RECT 683.385 278.145 683.555 278.315 ;
        RECT 683.865 278.145 684.035 278.315 ;
        RECT 684.345 278.145 684.515 278.315 ;
        RECT 696.825 278.155 696.995 278.325 ;
        RECT 697.305 278.155 697.475 278.325 ;
        RECT 697.785 278.155 697.955 278.325 ;
        RECT 698.265 278.155 698.435 278.325 ;
        RECT 698.745 278.155 698.915 278.325 ;
        RECT 699.225 278.155 699.395 278.325 ;
        RECT 699.705 278.155 699.875 278.325 ;
        RECT 700.185 278.155 700.355 278.325 ;
        RECT 700.665 278.155 700.835 278.325 ;
        RECT 701.145 278.155 701.315 278.325 ;
        RECT 701.625 278.155 701.795 278.325 ;
        RECT 714.595 278.155 714.765 278.325 ;
        RECT 715.075 278.155 715.245 278.325 ;
        RECT 715.555 278.155 715.725 278.325 ;
        RECT 716.035 278.155 716.205 278.325 ;
        RECT 716.515 278.155 716.685 278.325 ;
        RECT 716.995 278.155 717.165 278.325 ;
        RECT 717.475 278.155 717.645 278.325 ;
        RECT 717.955 278.155 718.125 278.325 ;
        RECT 718.435 278.155 718.605 278.325 ;
        RECT 718.915 278.155 719.085 278.325 ;
        RECT 719.395 278.155 719.565 278.325 ;
        RECT 731.835 278.155 732.005 278.325 ;
        RECT 732.315 278.155 732.485 278.325 ;
        RECT 732.795 278.155 732.965 278.325 ;
        RECT 733.275 278.155 733.445 278.325 ;
        RECT 733.755 278.155 733.925 278.325 ;
        RECT 734.235 278.155 734.405 278.325 ;
        RECT 734.715 278.155 734.885 278.325 ;
        RECT 735.195 278.155 735.365 278.325 ;
        RECT 735.675 278.155 735.845 278.325 ;
        RECT 736.155 278.155 736.325 278.325 ;
        RECT 736.635 278.155 736.805 278.325 ;
        RECT 749.315 278.165 749.485 278.335 ;
        RECT 749.795 278.165 749.965 278.335 ;
        RECT 750.275 278.165 750.445 278.335 ;
        RECT 750.755 278.165 750.925 278.335 ;
        RECT 751.235 278.165 751.405 278.335 ;
        RECT 751.715 278.165 751.885 278.335 ;
        RECT 752.195 278.165 752.365 278.335 ;
        RECT 752.675 278.165 752.845 278.335 ;
        RECT 753.155 278.165 753.325 278.335 ;
        RECT 753.635 278.165 753.805 278.335 ;
        RECT 754.115 278.165 754.285 278.335 ;
        RECT 857.615 278.295 857.785 278.465 ;
        RECT 857.975 278.295 858.145 278.465 ;
        RECT 858.335 278.295 858.505 278.465 ;
        RECT 856.085 277.815 856.255 277.985 ;
        RECT 856.565 277.815 856.735 277.985 ;
        RECT 857.045 277.815 857.215 277.985 ;
        RECT 857.525 277.815 857.695 277.985 ;
        RECT 858.005 277.815 858.175 277.985 ;
        RECT 858.485 277.815 858.655 277.985 ;
        RECT 858.965 277.815 859.135 277.985 ;
        RECT 115.150 276.500 115.320 276.670 ;
        RECT 115.150 276.140 115.320 276.310 ;
        RECT 115.150 275.780 115.320 275.950 ;
        RECT 115.150 275.420 115.320 275.590 ;
        RECT 115.150 275.060 115.320 275.230 ;
        RECT 751.665 274.720 751.835 274.890 ;
        RECT 118.365 274.490 118.535 274.660 ;
        RECT 118.725 274.490 118.895 274.660 ;
        RECT 121.835 274.490 122.005 274.660 ;
        RECT 122.195 274.490 122.365 274.660 ;
        RECT 125.305 274.490 125.475 274.660 ;
        RECT 125.665 274.490 125.835 274.660 ;
        RECT 128.775 274.490 128.945 274.660 ;
        RECT 129.135 274.490 129.305 274.660 ;
        RECT 132.245 274.490 132.415 274.660 ;
        RECT 132.605 274.490 132.775 274.660 ;
        RECT 135.715 274.490 135.885 274.660 ;
        RECT 136.075 274.490 136.245 274.660 ;
        RECT 139.185 274.490 139.355 274.660 ;
        RECT 139.545 274.490 139.715 274.660 ;
        RECT 142.655 274.490 142.825 274.660 ;
        RECT 143.015 274.490 143.185 274.660 ;
        RECT 146.125 274.490 146.295 274.660 ;
        RECT 146.485 274.490 146.655 274.660 ;
        RECT 149.595 274.490 149.765 274.660 ;
        RECT 149.955 274.490 150.125 274.660 ;
        RECT 679.920 272.965 680.090 273.135 ;
        RECT 680.280 272.965 680.450 273.135 ;
        RECT 681.140 272.965 681.310 273.135 ;
        RECT 681.500 272.965 681.670 273.135 ;
        RECT 681.860 272.965 682.030 273.135 ;
        RECT 682.220 272.965 682.390 273.135 ;
        RECT 682.580 272.965 682.750 273.135 ;
        RECT 682.940 272.965 683.110 273.135 ;
        RECT 683.300 272.965 683.470 273.135 ;
        RECT 684.380 272.965 684.550 273.135 ;
        RECT 684.740 272.965 684.910 273.135 ;
        RECT 687.160 272.925 687.330 273.095 ;
        RECT 687.520 272.925 687.690 273.095 ;
        RECT 688.380 272.925 688.550 273.095 ;
        RECT 688.740 272.925 688.910 273.095 ;
        RECT 689.100 272.925 689.270 273.095 ;
        RECT 689.460 272.925 689.630 273.095 ;
        RECT 689.820 272.925 689.990 273.095 ;
        RECT 690.180 272.925 690.350 273.095 ;
        RECT 690.540 272.925 690.710 273.095 ;
        RECT 691.620 272.925 691.790 273.095 ;
        RECT 691.980 272.925 692.150 273.095 ;
        RECT 697.150 272.985 697.320 273.155 ;
        RECT 697.510 272.985 697.680 273.155 ;
        RECT 698.370 272.985 698.540 273.155 ;
        RECT 698.730 272.985 698.900 273.155 ;
        RECT 699.090 272.985 699.260 273.155 ;
        RECT 699.450 272.985 699.620 273.155 ;
        RECT 699.810 272.985 699.980 273.155 ;
        RECT 700.170 272.985 700.340 273.155 ;
        RECT 700.530 272.985 700.700 273.155 ;
        RECT 701.610 272.985 701.780 273.155 ;
        RECT 701.970 272.985 702.140 273.155 ;
        RECT 704.390 272.945 704.560 273.115 ;
        RECT 704.750 272.945 704.920 273.115 ;
        RECT 705.610 272.945 705.780 273.115 ;
        RECT 705.970 272.945 706.140 273.115 ;
        RECT 706.330 272.945 706.500 273.115 ;
        RECT 706.690 272.945 706.860 273.115 ;
        RECT 707.050 272.945 707.220 273.115 ;
        RECT 707.410 272.945 707.580 273.115 ;
        RECT 707.770 272.945 707.940 273.115 ;
        RECT 708.850 272.945 709.020 273.115 ;
        RECT 709.210 272.945 709.380 273.115 ;
        RECT 714.720 273.085 714.890 273.255 ;
        RECT 715.080 273.085 715.250 273.255 ;
        RECT 715.940 273.085 716.110 273.255 ;
        RECT 716.300 273.085 716.470 273.255 ;
        RECT 716.660 273.085 716.830 273.255 ;
        RECT 717.020 273.085 717.190 273.255 ;
        RECT 717.380 273.085 717.550 273.255 ;
        RECT 717.740 273.085 717.910 273.255 ;
        RECT 718.100 273.085 718.270 273.255 ;
        RECT 719.180 273.085 719.350 273.255 ;
        RECT 719.540 273.085 719.710 273.255 ;
        RECT 721.960 273.045 722.130 273.215 ;
        RECT 722.320 273.045 722.490 273.215 ;
        RECT 723.180 273.045 723.350 273.215 ;
        RECT 723.540 273.045 723.710 273.215 ;
        RECT 723.900 273.045 724.070 273.215 ;
        RECT 724.260 273.045 724.430 273.215 ;
        RECT 724.620 273.045 724.790 273.215 ;
        RECT 724.980 273.045 725.150 273.215 ;
        RECT 725.340 273.045 725.510 273.215 ;
        RECT 726.420 273.045 726.590 273.215 ;
        RECT 726.780 273.045 726.950 273.215 ;
        RECT 731.890 273.115 732.060 273.285 ;
        RECT 732.250 273.115 732.420 273.285 ;
        RECT 733.110 273.115 733.280 273.285 ;
        RECT 733.470 273.115 733.640 273.285 ;
        RECT 733.830 273.115 734.000 273.285 ;
        RECT 734.190 273.115 734.360 273.285 ;
        RECT 734.550 273.115 734.720 273.285 ;
        RECT 734.910 273.115 735.080 273.285 ;
        RECT 735.270 273.115 735.440 273.285 ;
        RECT 736.350 273.115 736.520 273.285 ;
        RECT 736.710 273.115 736.880 273.285 ;
        RECT 739.130 273.075 739.300 273.245 ;
        RECT 739.490 273.075 739.660 273.245 ;
        RECT 740.350 273.075 740.520 273.245 ;
        RECT 740.710 273.075 740.880 273.245 ;
        RECT 741.070 273.075 741.240 273.245 ;
        RECT 741.430 273.075 741.600 273.245 ;
        RECT 741.790 273.075 741.960 273.245 ;
        RECT 742.150 273.075 742.320 273.245 ;
        RECT 742.510 273.075 742.680 273.245 ;
        RECT 743.590 273.075 743.760 273.245 ;
        RECT 743.950 273.075 744.120 273.245 ;
        RECT 749.700 273.175 749.870 273.345 ;
        RECT 750.060 273.175 750.230 273.345 ;
        RECT 750.920 273.175 751.090 273.345 ;
        RECT 751.280 273.175 751.450 273.345 ;
        RECT 751.640 273.175 751.810 273.345 ;
        RECT 752.000 273.175 752.170 273.345 ;
        RECT 752.360 273.175 752.530 273.345 ;
        RECT 752.720 273.175 752.890 273.345 ;
        RECT 753.080 273.175 753.250 273.345 ;
        RECT 754.160 273.175 754.330 273.345 ;
        RECT 754.520 273.175 754.690 273.345 ;
        RECT 756.940 273.135 757.110 273.305 ;
        RECT 757.300 273.135 757.470 273.305 ;
        RECT 758.160 273.135 758.330 273.305 ;
        RECT 758.520 273.135 758.690 273.305 ;
        RECT 758.880 273.135 759.050 273.305 ;
        RECT 759.240 273.135 759.410 273.305 ;
        RECT 759.600 273.135 759.770 273.305 ;
        RECT 759.960 273.135 760.130 273.305 ;
        RECT 760.320 273.135 760.490 273.305 ;
        RECT 761.400 273.135 761.570 273.305 ;
        RECT 761.760 273.135 761.930 273.305 ;
        RECT 635.100 271.735 635.270 271.905 ;
        RECT 635.460 271.735 635.630 271.905 ;
        RECT 639.290 271.825 639.460 271.995 ;
        RECT 639.650 271.825 639.820 271.995 ;
        RECT 679.955 272.485 680.125 272.655 ;
        RECT 680.435 272.485 680.605 272.655 ;
        RECT 680.915 272.485 681.085 272.655 ;
        RECT 681.395 272.485 681.565 272.655 ;
        RECT 681.875 272.485 682.045 272.655 ;
        RECT 682.355 272.485 682.525 272.655 ;
        RECT 682.835 272.485 683.005 272.655 ;
        RECT 683.315 272.485 683.485 272.655 ;
        RECT 683.795 272.485 683.965 272.655 ;
        RECT 684.275 272.485 684.445 272.655 ;
        RECT 684.755 272.485 684.925 272.655 ;
        RECT 687.195 272.445 687.365 272.615 ;
        RECT 687.675 272.445 687.845 272.615 ;
        RECT 688.155 272.445 688.325 272.615 ;
        RECT 688.635 272.445 688.805 272.615 ;
        RECT 689.115 272.445 689.285 272.615 ;
        RECT 689.595 272.445 689.765 272.615 ;
        RECT 690.075 272.445 690.245 272.615 ;
        RECT 690.555 272.445 690.725 272.615 ;
        RECT 691.035 272.445 691.205 272.615 ;
        RECT 691.515 272.445 691.685 272.615 ;
        RECT 691.995 272.445 692.165 272.615 ;
        RECT 697.185 272.505 697.355 272.675 ;
        RECT 697.665 272.505 697.835 272.675 ;
        RECT 698.145 272.505 698.315 272.675 ;
        RECT 698.625 272.505 698.795 272.675 ;
        RECT 699.105 272.505 699.275 272.675 ;
        RECT 699.585 272.505 699.755 272.675 ;
        RECT 700.065 272.505 700.235 272.675 ;
        RECT 700.545 272.505 700.715 272.675 ;
        RECT 701.025 272.505 701.195 272.675 ;
        RECT 701.505 272.505 701.675 272.675 ;
        RECT 701.985 272.505 702.155 272.675 ;
        RECT 704.425 272.465 704.595 272.635 ;
        RECT 704.905 272.465 705.075 272.635 ;
        RECT 705.385 272.465 705.555 272.635 ;
        RECT 705.865 272.465 706.035 272.635 ;
        RECT 706.345 272.465 706.515 272.635 ;
        RECT 706.825 272.465 706.995 272.635 ;
        RECT 707.305 272.465 707.475 272.635 ;
        RECT 707.785 272.465 707.955 272.635 ;
        RECT 708.265 272.465 708.435 272.635 ;
        RECT 708.745 272.465 708.915 272.635 ;
        RECT 709.225 272.465 709.395 272.635 ;
        RECT 714.755 272.605 714.925 272.775 ;
        RECT 715.235 272.605 715.405 272.775 ;
        RECT 715.715 272.605 715.885 272.775 ;
        RECT 716.195 272.605 716.365 272.775 ;
        RECT 716.675 272.605 716.845 272.775 ;
        RECT 717.155 272.605 717.325 272.775 ;
        RECT 717.635 272.605 717.805 272.775 ;
        RECT 718.115 272.605 718.285 272.775 ;
        RECT 718.595 272.605 718.765 272.775 ;
        RECT 719.075 272.605 719.245 272.775 ;
        RECT 719.555 272.605 719.725 272.775 ;
        RECT 721.995 272.565 722.165 272.735 ;
        RECT 722.475 272.565 722.645 272.735 ;
        RECT 722.955 272.565 723.125 272.735 ;
        RECT 723.435 272.565 723.605 272.735 ;
        RECT 723.915 272.565 724.085 272.735 ;
        RECT 724.395 272.565 724.565 272.735 ;
        RECT 724.875 272.565 725.045 272.735 ;
        RECT 725.355 272.565 725.525 272.735 ;
        RECT 725.835 272.565 726.005 272.735 ;
        RECT 726.315 272.565 726.485 272.735 ;
        RECT 726.795 272.565 726.965 272.735 ;
        RECT 731.925 272.635 732.095 272.805 ;
        RECT 732.405 272.635 732.575 272.805 ;
        RECT 732.885 272.635 733.055 272.805 ;
        RECT 733.365 272.635 733.535 272.805 ;
        RECT 733.845 272.635 734.015 272.805 ;
        RECT 734.325 272.635 734.495 272.805 ;
        RECT 734.805 272.635 734.975 272.805 ;
        RECT 735.285 272.635 735.455 272.805 ;
        RECT 735.765 272.635 735.935 272.805 ;
        RECT 736.245 272.635 736.415 272.805 ;
        RECT 736.725 272.635 736.895 272.805 ;
        RECT 739.165 272.595 739.335 272.765 ;
        RECT 739.645 272.595 739.815 272.765 ;
        RECT 740.125 272.595 740.295 272.765 ;
        RECT 740.605 272.595 740.775 272.765 ;
        RECT 741.085 272.595 741.255 272.765 ;
        RECT 741.565 272.595 741.735 272.765 ;
        RECT 742.045 272.595 742.215 272.765 ;
        RECT 742.525 272.595 742.695 272.765 ;
        RECT 743.005 272.595 743.175 272.765 ;
        RECT 743.485 272.595 743.655 272.765 ;
        RECT 743.965 272.595 744.135 272.765 ;
        RECT 749.735 272.695 749.905 272.865 ;
        RECT 750.215 272.695 750.385 272.865 ;
        RECT 750.695 272.695 750.865 272.865 ;
        RECT 751.175 272.695 751.345 272.865 ;
        RECT 751.655 272.695 751.825 272.865 ;
        RECT 752.135 272.695 752.305 272.865 ;
        RECT 752.615 272.695 752.785 272.865 ;
        RECT 753.095 272.695 753.265 272.865 ;
        RECT 753.575 272.695 753.745 272.865 ;
        RECT 754.055 272.695 754.225 272.865 ;
        RECT 754.535 272.695 754.705 272.865 ;
        RECT 756.975 272.655 757.145 272.825 ;
        RECT 757.455 272.655 757.625 272.825 ;
        RECT 757.935 272.655 758.105 272.825 ;
        RECT 758.415 272.655 758.585 272.825 ;
        RECT 758.895 272.655 759.065 272.825 ;
        RECT 759.375 272.655 759.545 272.825 ;
        RECT 759.855 272.655 760.025 272.825 ;
        RECT 760.335 272.655 760.505 272.825 ;
        RECT 760.815 272.655 760.985 272.825 ;
        RECT 761.295 272.655 761.465 272.825 ;
        RECT 761.775 272.655 761.945 272.825 ;
        RECT 643.390 271.805 643.560 271.975 ;
        RECT 643.750 271.805 643.920 271.975 ;
        RECT 781.550 271.805 781.720 271.975 ;
        RECT 781.910 271.805 782.080 271.975 ;
        RECT 782.270 271.805 782.440 271.975 ;
        RECT 783.190 271.805 783.360 271.975 ;
        RECT 783.550 271.805 783.720 271.975 ;
        RECT 788.150 271.805 788.320 271.975 ;
        RECT 788.510 271.805 788.680 271.975 ;
        RECT 788.870 271.805 789.040 271.975 ;
        RECT 792.120 271.805 792.290 271.975 ;
        RECT 792.480 271.805 792.650 271.975 ;
        RECT 792.840 271.805 793.010 271.975 ;
        RECT 794.725 271.805 794.895 271.975 ;
        RECT 795.085 271.805 795.255 271.975 ;
        RECT 795.445 271.805 795.615 271.975 ;
        RECT 800.440 271.795 800.610 271.965 ;
        RECT 800.800 271.795 800.970 271.965 ;
        RECT 801.160 271.795 801.330 271.965 ;
        RECT 802.080 271.795 802.250 271.965 ;
        RECT 802.440 271.795 802.610 271.965 ;
        RECT 807.040 271.795 807.210 271.965 ;
        RECT 807.400 271.795 807.570 271.965 ;
        RECT 807.760 271.795 807.930 271.965 ;
        RECT 811.010 271.795 811.180 271.965 ;
        RECT 811.370 271.795 811.540 271.965 ;
        RECT 811.730 271.795 811.900 271.965 ;
        RECT 813.615 271.795 813.785 271.965 ;
        RECT 813.975 271.795 814.145 271.965 ;
        RECT 814.335 271.795 814.505 271.965 ;
        RECT 819.290 271.765 819.460 271.935 ;
        RECT 819.650 271.765 819.820 271.935 ;
        RECT 820.010 271.765 820.180 271.935 ;
        RECT 820.930 271.765 821.100 271.935 ;
        RECT 821.290 271.765 821.460 271.935 ;
        RECT 825.890 271.765 826.060 271.935 ;
        RECT 826.250 271.765 826.420 271.935 ;
        RECT 826.610 271.765 826.780 271.935 ;
        RECT 829.860 271.765 830.030 271.935 ;
        RECT 830.220 271.765 830.390 271.935 ;
        RECT 830.580 271.765 830.750 271.935 ;
        RECT 832.465 271.765 832.635 271.935 ;
        RECT 832.825 271.765 832.995 271.935 ;
        RECT 833.185 271.765 833.355 271.935 ;
        RECT 840.905 271.805 841.075 271.975 ;
        RECT 841.435 271.805 841.605 271.975 ;
        RECT 857.615 271.755 857.785 271.925 ;
        RECT 857.975 271.755 858.145 271.925 ;
        RECT 858.335 271.755 858.505 271.925 ;
        RECT 595.880 271.285 596.050 271.455 ;
        RECT 596.240 271.285 596.410 271.455 ;
        RECT 595.245 270.805 595.415 270.975 ;
        RECT 595.725 270.805 595.895 270.975 ;
        RECT 596.205 270.805 596.375 270.975 ;
        RECT 144.235 270.085 144.405 270.255 ;
        RECT 144.595 270.085 144.765 270.255 ;
        RECT 144.955 270.085 145.125 270.255 ;
        RECT 145.315 270.085 145.485 270.255 ;
        RECT 145.675 270.085 145.845 270.255 ;
        RECT 146.035 270.085 146.205 270.255 ;
        RECT 146.395 270.085 146.565 270.255 ;
        RECT 146.755 270.085 146.925 270.255 ;
        RECT 147.115 270.085 147.285 270.255 ;
        RECT 596.350 270.085 596.520 270.255 ;
        RECT 596.710 270.085 596.880 270.255 ;
        RECT 122.155 269.545 122.325 269.715 ;
        RECT 122.515 269.545 122.685 269.715 ;
        RECT 122.875 269.545 123.045 269.715 ;
        RECT 123.235 269.545 123.405 269.715 ;
        RECT 123.595 269.545 123.765 269.715 ;
        RECT 123.955 269.545 124.125 269.715 ;
        RECT 124.315 269.545 124.485 269.715 ;
        RECT 124.675 269.545 124.845 269.715 ;
        RECT 125.035 269.545 125.205 269.715 ;
        RECT 118.445 268.070 118.615 268.240 ;
        RECT 118.805 268.070 118.975 268.240 ;
        RECT 121.915 268.070 122.085 268.240 ;
        RECT 122.275 268.070 122.445 268.240 ;
        RECT 125.385 268.070 125.555 268.240 ;
        RECT 125.745 268.070 125.915 268.240 ;
        RECT 128.855 268.070 129.025 268.240 ;
        RECT 129.215 268.070 129.385 268.240 ;
        RECT 132.325 268.070 132.495 268.240 ;
        RECT 132.685 268.070 132.855 268.240 ;
        RECT 135.795 268.070 135.965 268.240 ;
        RECT 136.155 268.070 136.325 268.240 ;
        RECT 139.265 268.070 139.435 268.240 ;
        RECT 139.625 268.070 139.795 268.240 ;
        RECT 142.735 268.070 142.905 268.240 ;
        RECT 143.095 268.070 143.265 268.240 ;
        RECT 146.205 268.070 146.375 268.240 ;
        RECT 146.565 268.070 146.735 268.240 ;
        RECT 149.675 268.070 149.845 268.240 ;
        RECT 150.035 268.070 150.205 268.240 ;
        RECT 605.215 267.075 605.745 270.485 ;
        RECT 635.135 271.255 635.305 271.425 ;
        RECT 635.615 271.255 635.785 271.425 ;
        RECT 636.095 271.255 636.265 271.425 ;
        RECT 639.325 271.345 639.495 271.515 ;
        RECT 639.805 271.345 639.975 271.515 ;
        RECT 640.285 271.345 640.455 271.515 ;
        RECT 643.425 271.325 643.595 271.495 ;
        RECT 643.905 271.325 644.075 271.495 ;
        RECT 644.385 271.325 644.555 271.495 ;
        RECT 781.115 271.325 781.285 271.495 ;
        RECT 781.595 271.325 781.765 271.495 ;
        RECT 782.075 271.325 782.245 271.495 ;
        RECT 782.555 271.325 782.725 271.495 ;
        RECT 783.035 271.325 783.205 271.495 ;
        RECT 783.515 271.325 783.685 271.495 ;
        RECT 783.995 271.325 784.165 271.495 ;
        RECT 784.475 271.325 784.645 271.495 ;
        RECT 784.955 271.325 785.125 271.495 ;
        RECT 785.435 271.325 785.605 271.495 ;
        RECT 785.915 271.325 786.085 271.495 ;
        RECT 786.395 271.325 786.565 271.495 ;
        RECT 786.875 271.325 787.045 271.495 ;
        RECT 787.355 271.325 787.525 271.495 ;
        RECT 787.835 271.325 788.005 271.495 ;
        RECT 788.315 271.325 788.485 271.495 ;
        RECT 788.795 271.325 788.965 271.495 ;
        RECT 789.275 271.325 789.445 271.495 ;
        RECT 789.755 271.325 789.925 271.495 ;
        RECT 790.235 271.325 790.405 271.495 ;
        RECT 790.715 271.325 790.885 271.495 ;
        RECT 791.195 271.325 791.365 271.495 ;
        RECT 791.675 271.325 791.845 271.495 ;
        RECT 792.155 271.325 792.325 271.495 ;
        RECT 792.635 271.325 792.805 271.495 ;
        RECT 793.115 271.325 793.285 271.495 ;
        RECT 793.595 271.325 793.765 271.495 ;
        RECT 794.075 271.325 794.245 271.495 ;
        RECT 794.555 271.325 794.725 271.495 ;
        RECT 795.035 271.325 795.205 271.495 ;
        RECT 795.515 271.325 795.685 271.495 ;
        RECT 795.995 271.325 796.165 271.495 ;
        RECT 800.005 271.315 800.175 271.485 ;
        RECT 800.485 271.315 800.655 271.485 ;
        RECT 800.965 271.315 801.135 271.485 ;
        RECT 801.445 271.315 801.615 271.485 ;
        RECT 801.925 271.315 802.095 271.485 ;
        RECT 802.405 271.315 802.575 271.485 ;
        RECT 802.885 271.315 803.055 271.485 ;
        RECT 803.365 271.315 803.535 271.485 ;
        RECT 803.845 271.315 804.015 271.485 ;
        RECT 804.325 271.315 804.495 271.485 ;
        RECT 804.805 271.315 804.975 271.485 ;
        RECT 805.285 271.315 805.455 271.485 ;
        RECT 805.765 271.315 805.935 271.485 ;
        RECT 806.245 271.315 806.415 271.485 ;
        RECT 806.725 271.315 806.895 271.485 ;
        RECT 807.205 271.315 807.375 271.485 ;
        RECT 807.685 271.315 807.855 271.485 ;
        RECT 808.165 271.315 808.335 271.485 ;
        RECT 808.645 271.315 808.815 271.485 ;
        RECT 809.125 271.315 809.295 271.485 ;
        RECT 809.605 271.315 809.775 271.485 ;
        RECT 810.085 271.315 810.255 271.485 ;
        RECT 810.565 271.315 810.735 271.485 ;
        RECT 811.045 271.315 811.215 271.485 ;
        RECT 811.525 271.315 811.695 271.485 ;
        RECT 812.005 271.315 812.175 271.485 ;
        RECT 812.485 271.315 812.655 271.485 ;
        RECT 812.965 271.315 813.135 271.485 ;
        RECT 813.445 271.315 813.615 271.485 ;
        RECT 813.925 271.315 814.095 271.485 ;
        RECT 814.405 271.315 814.575 271.485 ;
        RECT 814.885 271.315 815.055 271.485 ;
        RECT 818.855 271.285 819.025 271.455 ;
        RECT 819.335 271.285 819.505 271.455 ;
        RECT 819.815 271.285 819.985 271.455 ;
        RECT 820.295 271.285 820.465 271.455 ;
        RECT 820.775 271.285 820.945 271.455 ;
        RECT 821.255 271.285 821.425 271.455 ;
        RECT 821.735 271.285 821.905 271.455 ;
        RECT 822.215 271.285 822.385 271.455 ;
        RECT 822.695 271.285 822.865 271.455 ;
        RECT 823.175 271.285 823.345 271.455 ;
        RECT 823.655 271.285 823.825 271.455 ;
        RECT 824.135 271.285 824.305 271.455 ;
        RECT 824.615 271.285 824.785 271.455 ;
        RECT 825.095 271.285 825.265 271.455 ;
        RECT 825.575 271.285 825.745 271.455 ;
        RECT 826.055 271.285 826.225 271.455 ;
        RECT 826.535 271.285 826.705 271.455 ;
        RECT 827.015 271.285 827.185 271.455 ;
        RECT 827.495 271.285 827.665 271.455 ;
        RECT 827.975 271.285 828.145 271.455 ;
        RECT 828.455 271.285 828.625 271.455 ;
        RECT 828.935 271.285 829.105 271.455 ;
        RECT 829.415 271.285 829.585 271.455 ;
        RECT 829.895 271.285 830.065 271.455 ;
        RECT 830.375 271.285 830.545 271.455 ;
        RECT 830.855 271.285 831.025 271.455 ;
        RECT 831.335 271.285 831.505 271.455 ;
        RECT 831.815 271.285 831.985 271.455 ;
        RECT 832.295 271.285 832.465 271.455 ;
        RECT 832.775 271.285 832.945 271.455 ;
        RECT 833.255 271.285 833.425 271.455 ;
        RECT 833.735 271.285 833.905 271.455 ;
        RECT 838.575 271.325 838.745 271.495 ;
        RECT 839.055 271.325 839.225 271.495 ;
        RECT 839.535 271.325 839.705 271.495 ;
        RECT 840.015 271.325 840.185 271.495 ;
        RECT 840.495 271.325 840.665 271.495 ;
        RECT 840.975 271.325 841.145 271.495 ;
        RECT 841.455 271.325 841.625 271.495 ;
        RECT 841.935 271.325 842.105 271.495 ;
        RECT 856.085 271.275 856.255 271.445 ;
        RECT 856.565 271.275 856.735 271.445 ;
        RECT 857.045 271.275 857.215 271.445 ;
        RECT 857.525 271.275 857.695 271.445 ;
        RECT 858.005 271.275 858.175 271.445 ;
        RECT 858.485 271.275 858.655 271.445 ;
        RECT 858.965 271.275 859.135 271.445 ;
        RECT 625.620 270.415 625.790 270.585 ;
        RECT 625.620 270.055 625.790 270.225 ;
        RECT 625.620 269.695 625.790 269.865 ;
        RECT 846.355 269.545 846.525 269.715 ;
        RECT 846.715 269.545 846.885 269.715 ;
        RECT 847.075 269.545 847.245 269.715 ;
        RECT 850.200 269.555 850.370 269.725 ;
        RECT 850.560 269.555 850.730 269.725 ;
        RECT 625.620 269.335 625.790 269.505 ;
        RECT 625.620 268.975 625.790 269.145 ;
        RECT 844.825 269.065 844.995 269.235 ;
        RECT 845.305 269.065 845.475 269.235 ;
        RECT 845.785 269.065 845.955 269.235 ;
        RECT 846.265 269.065 846.435 269.235 ;
        RECT 846.745 269.065 846.915 269.235 ;
        RECT 847.225 269.065 847.395 269.235 ;
        RECT 847.705 269.065 847.875 269.235 ;
        RECT 850.235 269.075 850.405 269.245 ;
        RECT 850.715 269.075 850.885 269.245 ;
        RECT 851.195 269.075 851.365 269.245 ;
        RECT 614.740 268.605 614.910 268.775 ;
        RECT 616.320 268.605 616.490 268.775 ;
        RECT 625.620 268.615 625.790 268.785 ;
        RECT 625.620 268.255 625.790 268.425 ;
        RECT 749.925 268.550 750.095 268.720 ;
        RECT 625.620 267.895 625.790 268.065 ;
        RECT 625.620 267.535 625.790 267.705 ;
        RECT 640.090 267.715 640.260 267.885 ;
        RECT 644.140 267.765 644.310 267.935 ;
        RECT 614.740 267.135 614.910 267.305 ;
        RECT 616.320 267.135 616.490 267.305 ;
        RECT 681.605 267.285 681.775 267.455 ;
        RECT 681.965 267.285 682.135 267.455 ;
        RECT 682.325 267.285 682.495 267.455 ;
        RECT 687.265 267.295 687.435 267.465 ;
        RECT 687.625 267.295 687.795 267.465 ;
        RECT 687.985 267.295 688.155 267.465 ;
        RECT 691.030 267.315 691.200 267.485 ;
        RECT 691.390 267.315 691.560 267.485 ;
        RECT 691.750 267.315 691.920 267.485 ;
        RECT 693.000 267.315 693.170 267.485 ;
        RECT 693.360 267.315 693.530 267.485 ;
        RECT 698.835 267.305 699.005 267.475 ;
        RECT 699.195 267.305 699.365 267.475 ;
        RECT 699.555 267.305 699.725 267.475 ;
        RECT 704.495 267.315 704.665 267.485 ;
        RECT 704.855 267.315 705.025 267.485 ;
        RECT 705.215 267.315 705.385 267.485 ;
        RECT 708.260 267.335 708.430 267.505 ;
        RECT 708.620 267.335 708.790 267.505 ;
        RECT 708.980 267.335 709.150 267.505 ;
        RECT 710.230 267.335 710.400 267.505 ;
        RECT 710.590 267.335 710.760 267.505 ;
        RECT 716.405 267.405 716.575 267.575 ;
        RECT 716.765 267.405 716.935 267.575 ;
        RECT 717.125 267.405 717.295 267.575 ;
        RECT 722.065 267.415 722.235 267.585 ;
        RECT 722.425 267.415 722.595 267.585 ;
        RECT 722.785 267.415 722.955 267.585 ;
        RECT 725.830 267.435 726.000 267.605 ;
        RECT 726.190 267.435 726.360 267.605 ;
        RECT 726.550 267.435 726.720 267.605 ;
        RECT 727.800 267.435 727.970 267.605 ;
        RECT 728.160 267.435 728.330 267.605 ;
        RECT 733.575 267.435 733.745 267.605 ;
        RECT 733.935 267.435 734.105 267.605 ;
        RECT 734.295 267.435 734.465 267.605 ;
        RECT 739.235 267.445 739.405 267.615 ;
        RECT 739.595 267.445 739.765 267.615 ;
        RECT 739.955 267.445 740.125 267.615 ;
        RECT 743.000 267.465 743.170 267.635 ;
        RECT 743.360 267.465 743.530 267.635 ;
        RECT 743.720 267.465 743.890 267.635 ;
        RECT 744.970 267.465 745.140 267.635 ;
        RECT 745.330 267.465 745.500 267.635 ;
        RECT 751.385 267.495 751.555 267.665 ;
        RECT 751.745 267.495 751.915 267.665 ;
        RECT 752.105 267.495 752.275 267.665 ;
        RECT 757.045 267.505 757.215 267.675 ;
        RECT 757.405 267.505 757.575 267.675 ;
        RECT 757.765 267.505 757.935 267.675 ;
        RECT 760.810 267.525 760.980 267.695 ;
        RECT 761.170 267.525 761.340 267.695 ;
        RECT 761.530 267.525 761.700 267.695 ;
        RECT 861.350 268.365 861.520 268.535 ;
        RECT 861.710 268.365 861.880 268.535 ;
        RECT 862.070 268.365 862.240 268.535 ;
        RECT 863.320 268.365 863.490 268.535 ;
        RECT 863.680 268.365 863.850 268.535 ;
        RECT 861.405 267.885 861.575 268.055 ;
        RECT 861.885 267.885 862.055 268.055 ;
        RECT 862.365 267.885 862.535 268.055 ;
        RECT 862.845 267.885 863.015 268.055 ;
        RECT 863.325 267.885 863.495 268.055 ;
        RECT 863.805 267.885 863.975 268.055 ;
        RECT 864.285 267.885 864.455 268.055 ;
        RECT 762.780 267.525 762.950 267.695 ;
        RECT 763.140 267.525 763.310 267.695 ;
        RECT 680.075 266.805 680.245 266.975 ;
        RECT 680.555 266.805 680.725 266.975 ;
        RECT 681.035 266.805 681.205 266.975 ;
        RECT 681.515 266.805 681.685 266.975 ;
        RECT 681.995 266.805 682.165 266.975 ;
        RECT 682.475 266.805 682.645 266.975 ;
        RECT 682.955 266.805 683.125 266.975 ;
        RECT 685.735 266.815 685.905 266.985 ;
        RECT 686.215 266.815 686.385 266.985 ;
        RECT 686.695 266.815 686.865 266.985 ;
        RECT 687.175 266.815 687.345 266.985 ;
        RECT 687.655 266.815 687.825 266.985 ;
        RECT 688.135 266.815 688.305 266.985 ;
        RECT 688.615 266.815 688.785 266.985 ;
        RECT 691.085 266.835 691.255 267.005 ;
        RECT 691.565 266.835 691.735 267.005 ;
        RECT 692.045 266.835 692.215 267.005 ;
        RECT 692.525 266.835 692.695 267.005 ;
        RECT 693.005 266.835 693.175 267.005 ;
        RECT 693.485 266.835 693.655 267.005 ;
        RECT 693.965 266.835 694.135 267.005 ;
        RECT 697.305 266.825 697.475 266.995 ;
        RECT 697.785 266.825 697.955 266.995 ;
        RECT 698.265 266.825 698.435 266.995 ;
        RECT 698.745 266.825 698.915 266.995 ;
        RECT 699.225 266.825 699.395 266.995 ;
        RECT 699.705 266.825 699.875 266.995 ;
        RECT 700.185 266.825 700.355 266.995 ;
        RECT 702.965 266.835 703.135 267.005 ;
        RECT 703.445 266.835 703.615 267.005 ;
        RECT 703.925 266.835 704.095 267.005 ;
        RECT 704.405 266.835 704.575 267.005 ;
        RECT 704.885 266.835 705.055 267.005 ;
        RECT 705.365 266.835 705.535 267.005 ;
        RECT 705.845 266.835 706.015 267.005 ;
        RECT 708.315 266.855 708.485 267.025 ;
        RECT 708.795 266.855 708.965 267.025 ;
        RECT 709.275 266.855 709.445 267.025 ;
        RECT 709.755 266.855 709.925 267.025 ;
        RECT 710.235 266.855 710.405 267.025 ;
        RECT 710.715 266.855 710.885 267.025 ;
        RECT 711.195 266.855 711.365 267.025 ;
        RECT 714.875 266.925 715.045 267.095 ;
        RECT 715.355 266.925 715.525 267.095 ;
        RECT 715.835 266.925 716.005 267.095 ;
        RECT 716.315 266.925 716.485 267.095 ;
        RECT 716.795 266.925 716.965 267.095 ;
        RECT 717.275 266.925 717.445 267.095 ;
        RECT 717.755 266.925 717.925 267.095 ;
        RECT 720.535 266.935 720.705 267.105 ;
        RECT 721.015 266.935 721.185 267.105 ;
        RECT 721.495 266.935 721.665 267.105 ;
        RECT 721.975 266.935 722.145 267.105 ;
        RECT 722.455 266.935 722.625 267.105 ;
        RECT 722.935 266.935 723.105 267.105 ;
        RECT 723.415 266.935 723.585 267.105 ;
        RECT 725.885 266.955 726.055 267.125 ;
        RECT 726.365 266.955 726.535 267.125 ;
        RECT 726.845 266.955 727.015 267.125 ;
        RECT 727.325 266.955 727.495 267.125 ;
        RECT 727.805 266.955 727.975 267.125 ;
        RECT 728.285 266.955 728.455 267.125 ;
        RECT 728.765 266.955 728.935 267.125 ;
        RECT 732.045 266.955 732.215 267.125 ;
        RECT 732.525 266.955 732.695 267.125 ;
        RECT 733.005 266.955 733.175 267.125 ;
        RECT 733.485 266.955 733.655 267.125 ;
        RECT 733.965 266.955 734.135 267.125 ;
        RECT 734.445 266.955 734.615 267.125 ;
        RECT 734.925 266.955 735.095 267.125 ;
        RECT 737.705 266.965 737.875 267.135 ;
        RECT 738.185 266.965 738.355 267.135 ;
        RECT 738.665 266.965 738.835 267.135 ;
        RECT 739.145 266.965 739.315 267.135 ;
        RECT 739.625 266.965 739.795 267.135 ;
        RECT 740.105 266.965 740.275 267.135 ;
        RECT 740.585 266.965 740.755 267.135 ;
        RECT 743.055 266.985 743.225 267.155 ;
        RECT 743.535 266.985 743.705 267.155 ;
        RECT 744.015 266.985 744.185 267.155 ;
        RECT 744.495 266.985 744.665 267.155 ;
        RECT 744.975 266.985 745.145 267.155 ;
        RECT 745.455 266.985 745.625 267.155 ;
        RECT 745.935 266.985 746.105 267.155 ;
        RECT 749.855 267.015 750.025 267.185 ;
        RECT 750.335 267.015 750.505 267.185 ;
        RECT 750.815 267.015 750.985 267.185 ;
        RECT 751.295 267.015 751.465 267.185 ;
        RECT 751.775 267.015 751.945 267.185 ;
        RECT 752.255 267.015 752.425 267.185 ;
        RECT 752.735 267.015 752.905 267.185 ;
        RECT 755.515 267.025 755.685 267.195 ;
        RECT 755.995 267.025 756.165 267.195 ;
        RECT 756.475 267.025 756.645 267.195 ;
        RECT 756.955 267.025 757.125 267.195 ;
        RECT 757.435 267.025 757.605 267.195 ;
        RECT 757.915 267.025 758.085 267.195 ;
        RECT 758.395 267.025 758.565 267.195 ;
        RECT 760.865 267.045 761.035 267.215 ;
        RECT 761.345 267.045 761.515 267.215 ;
        RECT 761.825 267.045 761.995 267.215 ;
        RECT 762.305 267.045 762.475 267.215 ;
        RECT 762.785 267.045 762.955 267.215 ;
        RECT 763.265 267.045 763.435 267.215 ;
        RECT 763.745 267.045 763.915 267.215 ;
        RECT 840.115 266.245 840.285 266.415 ;
        RECT 840.475 266.245 840.645 266.415 ;
        RECT 840.835 266.245 841.005 266.415 ;
        RECT 838.585 265.765 838.755 265.935 ;
        RECT 839.065 265.765 839.235 265.935 ;
        RECT 839.545 265.765 839.715 265.935 ;
        RECT 840.025 265.765 840.195 265.935 ;
        RECT 840.505 265.765 840.675 265.935 ;
        RECT 840.985 265.765 841.155 265.935 ;
        RECT 841.465 265.765 841.635 265.935 ;
        RECT 118.445 264.780 118.615 264.950 ;
        RECT 118.805 264.780 118.975 264.950 ;
        RECT 121.915 264.780 122.085 264.950 ;
        RECT 122.275 264.780 122.445 264.950 ;
        RECT 125.385 264.780 125.555 264.950 ;
        RECT 125.745 264.780 125.915 264.950 ;
        RECT 128.855 264.780 129.025 264.950 ;
        RECT 129.215 264.780 129.385 264.950 ;
        RECT 132.325 264.780 132.495 264.950 ;
        RECT 132.685 264.780 132.855 264.950 ;
        RECT 135.795 264.780 135.965 264.950 ;
        RECT 136.155 264.780 136.325 264.950 ;
        RECT 139.265 264.780 139.435 264.950 ;
        RECT 139.625 264.780 139.795 264.950 ;
        RECT 142.735 264.780 142.905 264.950 ;
        RECT 143.095 264.780 143.265 264.950 ;
        RECT 146.205 264.780 146.375 264.950 ;
        RECT 146.565 264.780 146.735 264.950 ;
        RECT 149.675 264.780 149.845 264.950 ;
        RECT 150.035 264.780 150.205 264.950 ;
        RECT 152.000 264.945 152.170 265.115 ;
        RECT 781.560 264.245 781.730 264.415 ;
        RECT 781.920 264.245 782.090 264.415 ;
        RECT 782.280 264.245 782.450 264.415 ;
        RECT 783.200 264.245 783.370 264.415 ;
        RECT 783.560 264.245 783.730 264.415 ;
        RECT 788.160 264.245 788.330 264.415 ;
        RECT 788.520 264.245 788.690 264.415 ;
        RECT 788.880 264.245 789.050 264.415 ;
        RECT 792.130 264.245 792.300 264.415 ;
        RECT 792.490 264.245 792.660 264.415 ;
        RECT 792.850 264.245 793.020 264.415 ;
        RECT 794.735 264.245 794.905 264.415 ;
        RECT 795.095 264.245 795.265 264.415 ;
        RECT 795.455 264.245 795.625 264.415 ;
        RECT 800.090 264.305 800.260 264.475 ;
        RECT 800.450 264.305 800.620 264.475 ;
        RECT 800.810 264.305 800.980 264.475 ;
        RECT 801.730 264.305 801.900 264.475 ;
        RECT 802.090 264.305 802.260 264.475 ;
        RECT 806.690 264.305 806.860 264.475 ;
        RECT 807.050 264.305 807.220 264.475 ;
        RECT 807.410 264.305 807.580 264.475 ;
        RECT 810.660 264.305 810.830 264.475 ;
        RECT 811.020 264.305 811.190 264.475 ;
        RECT 811.380 264.305 811.550 264.475 ;
        RECT 857.695 265.085 857.865 265.255 ;
        RECT 858.055 265.085 858.225 265.255 ;
        RECT 858.415 265.085 858.585 265.255 ;
        RECT 856.165 264.605 856.335 264.775 ;
        RECT 856.645 264.605 856.815 264.775 ;
        RECT 857.125 264.605 857.295 264.775 ;
        RECT 857.605 264.605 857.775 264.775 ;
        RECT 858.085 264.605 858.255 264.775 ;
        RECT 858.565 264.605 858.735 264.775 ;
        RECT 859.045 264.605 859.215 264.775 ;
        RECT 813.265 264.305 813.435 264.475 ;
        RECT 813.625 264.305 813.795 264.475 ;
        RECT 813.985 264.305 814.155 264.475 ;
        RECT 781.125 263.765 781.295 263.935 ;
        RECT 781.605 263.765 781.775 263.935 ;
        RECT 782.085 263.765 782.255 263.935 ;
        RECT 782.565 263.765 782.735 263.935 ;
        RECT 783.045 263.765 783.215 263.935 ;
        RECT 783.525 263.765 783.695 263.935 ;
        RECT 784.005 263.765 784.175 263.935 ;
        RECT 784.485 263.765 784.655 263.935 ;
        RECT 784.965 263.765 785.135 263.935 ;
        RECT 785.445 263.765 785.615 263.935 ;
        RECT 785.925 263.765 786.095 263.935 ;
        RECT 786.405 263.765 786.575 263.935 ;
        RECT 786.885 263.765 787.055 263.935 ;
        RECT 787.365 263.765 787.535 263.935 ;
        RECT 787.845 263.765 788.015 263.935 ;
        RECT 788.325 263.765 788.495 263.935 ;
        RECT 788.805 263.765 788.975 263.935 ;
        RECT 789.285 263.765 789.455 263.935 ;
        RECT 789.765 263.765 789.935 263.935 ;
        RECT 790.245 263.765 790.415 263.935 ;
        RECT 790.725 263.765 790.895 263.935 ;
        RECT 791.205 263.765 791.375 263.935 ;
        RECT 791.685 263.765 791.855 263.935 ;
        RECT 792.165 263.765 792.335 263.935 ;
        RECT 792.645 263.765 792.815 263.935 ;
        RECT 793.125 263.765 793.295 263.935 ;
        RECT 793.605 263.765 793.775 263.935 ;
        RECT 794.085 263.765 794.255 263.935 ;
        RECT 794.565 263.765 794.735 263.935 ;
        RECT 795.045 263.765 795.215 263.935 ;
        RECT 795.525 263.765 795.695 263.935 ;
        RECT 796.005 263.765 796.175 263.935 ;
        RECT 799.655 263.825 799.825 263.995 ;
        RECT 800.135 263.825 800.305 263.995 ;
        RECT 800.615 263.825 800.785 263.995 ;
        RECT 801.095 263.825 801.265 263.995 ;
        RECT 801.575 263.825 801.745 263.995 ;
        RECT 802.055 263.825 802.225 263.995 ;
        RECT 802.535 263.825 802.705 263.995 ;
        RECT 803.015 263.825 803.185 263.995 ;
        RECT 803.495 263.825 803.665 263.995 ;
        RECT 803.975 263.825 804.145 263.995 ;
        RECT 804.455 263.825 804.625 263.995 ;
        RECT 804.935 263.825 805.105 263.995 ;
        RECT 805.415 263.825 805.585 263.995 ;
        RECT 805.895 263.825 806.065 263.995 ;
        RECT 806.375 263.825 806.545 263.995 ;
        RECT 806.855 263.825 807.025 263.995 ;
        RECT 807.335 263.825 807.505 263.995 ;
        RECT 807.815 263.825 807.985 263.995 ;
        RECT 808.295 263.825 808.465 263.995 ;
        RECT 808.775 263.825 808.945 263.995 ;
        RECT 809.255 263.825 809.425 263.995 ;
        RECT 809.735 263.825 809.905 263.995 ;
        RECT 810.215 263.825 810.385 263.995 ;
        RECT 810.695 263.825 810.865 263.995 ;
        RECT 811.175 263.825 811.345 263.995 ;
        RECT 811.655 263.825 811.825 263.995 ;
        RECT 812.135 263.825 812.305 263.995 ;
        RECT 812.615 263.825 812.785 263.995 ;
        RECT 813.095 263.825 813.265 263.995 ;
        RECT 813.575 263.825 813.745 263.995 ;
        RECT 814.055 263.825 814.225 263.995 ;
        RECT 814.535 263.825 814.705 263.995 ;
        RECT 118.445 261.490 118.615 261.660 ;
        RECT 118.805 261.490 118.975 261.660 ;
        RECT 121.915 261.490 122.085 261.660 ;
        RECT 122.275 261.490 122.445 261.660 ;
        RECT 125.385 261.490 125.555 261.660 ;
        RECT 125.745 261.490 125.915 261.660 ;
        RECT 128.855 261.490 129.025 261.660 ;
        RECT 129.215 261.490 129.385 261.660 ;
        RECT 132.325 261.490 132.495 261.660 ;
        RECT 132.685 261.490 132.855 261.660 ;
        RECT 135.795 261.490 135.965 261.660 ;
        RECT 136.155 261.490 136.325 261.660 ;
        RECT 139.265 261.490 139.435 261.660 ;
        RECT 139.625 261.490 139.795 261.660 ;
        RECT 142.735 261.490 142.905 261.660 ;
        RECT 143.095 261.490 143.265 261.660 ;
        RECT 146.205 261.490 146.375 261.660 ;
        RECT 146.565 261.490 146.735 261.660 ;
        RECT 149.675 261.490 149.845 261.660 ;
        RECT 150.035 261.490 150.205 261.660 ;
        RECT 144.315 260.375 144.485 260.545 ;
        RECT 144.675 260.375 144.845 260.545 ;
        RECT 145.035 260.375 145.205 260.545 ;
        RECT 145.395 260.375 145.565 260.545 ;
        RECT 145.755 260.375 145.925 260.545 ;
        RECT 146.115 260.375 146.285 260.545 ;
        RECT 146.475 260.375 146.645 260.545 ;
        RECT 146.835 260.375 147.005 260.545 ;
        RECT 147.195 260.375 147.365 260.545 ;
        RECT 122.235 259.835 122.405 260.005 ;
        RECT 122.595 259.835 122.765 260.005 ;
        RECT 122.955 259.835 123.125 260.005 ;
        RECT 123.315 259.835 123.485 260.005 ;
        RECT 123.675 259.835 123.845 260.005 ;
        RECT 124.035 259.835 124.205 260.005 ;
        RECT 124.395 259.835 124.565 260.005 ;
        RECT 124.755 259.835 124.925 260.005 ;
        RECT 125.115 259.835 125.285 260.005 ;
        RECT -97.850 234.195 -97.680 234.365 ;
        RECT -97.850 233.835 -97.680 234.005 ;
        RECT -97.850 233.475 -97.680 233.645 ;
        RECT -97.850 233.115 -97.680 233.285 ;
        RECT -95.270 234.195 -95.100 234.365 ;
        RECT -95.270 233.835 -95.100 234.005 ;
        RECT -95.270 233.475 -95.100 233.645 ;
        RECT -95.270 233.115 -95.100 233.285 ;
        RECT -92.690 234.195 -92.520 234.365 ;
        RECT -92.690 233.835 -92.520 234.005 ;
        RECT -92.690 233.475 -92.520 233.645 ;
        RECT -92.690 233.115 -92.520 233.285 ;
        RECT -90.110 234.195 -89.940 234.365 ;
        RECT -90.110 233.835 -89.940 234.005 ;
        RECT -90.110 233.475 -89.940 233.645 ;
        RECT -90.110 233.115 -89.940 233.285 ;
        RECT -87.530 234.195 -87.360 234.365 ;
        RECT -87.530 233.835 -87.360 234.005 ;
        RECT -87.530 233.475 -87.360 233.645 ;
        RECT -87.530 233.115 -87.360 233.285 ;
        RECT -84.950 234.195 -84.780 234.365 ;
        RECT -84.950 233.835 -84.780 234.005 ;
        RECT -84.950 233.475 -84.780 233.645 ;
        RECT -84.950 233.115 -84.780 233.285 ;
        RECT -82.370 234.195 -82.200 234.365 ;
        RECT -82.370 233.835 -82.200 234.005 ;
        RECT -82.370 233.475 -82.200 233.645 ;
        RECT -82.370 233.115 -82.200 233.285 ;
        RECT -79.790 234.195 -79.620 234.365 ;
        RECT -79.790 233.835 -79.620 234.005 ;
        RECT -79.790 233.475 -79.620 233.645 ;
        RECT -79.790 233.115 -79.620 233.285 ;
        RECT -77.210 234.195 -77.040 234.365 ;
        RECT -77.210 233.835 -77.040 234.005 ;
        RECT -77.210 233.475 -77.040 233.645 ;
        RECT -77.210 233.115 -77.040 233.285 ;
        RECT -74.630 234.195 -74.460 234.365 ;
        RECT -74.630 233.835 -74.460 234.005 ;
        RECT -74.630 233.475 -74.460 233.645 ;
        RECT -74.630 233.115 -74.460 233.285 ;
        RECT -72.050 234.195 -71.880 234.365 ;
        RECT -72.050 233.835 -71.880 234.005 ;
        RECT -72.050 233.475 -71.880 233.645 ;
        RECT -72.050 233.115 -71.880 233.285 ;
        RECT -97.205 230.880 -97.035 231.050 ;
        RECT -95.915 230.880 -95.745 231.050 ;
        RECT -94.625 230.880 -94.455 231.050 ;
        RECT -93.335 230.880 -93.165 231.050 ;
        RECT -92.045 230.880 -91.875 231.050 ;
        RECT -90.755 230.880 -90.585 231.050 ;
        RECT -89.465 230.880 -89.295 231.050 ;
        RECT -88.175 230.880 -88.005 231.050 ;
        RECT -86.885 230.880 -86.715 231.050 ;
        RECT -85.595 230.880 -85.425 231.050 ;
        RECT -84.305 230.880 -84.135 231.050 ;
        RECT -83.015 230.880 -82.845 231.050 ;
        RECT -81.725 230.880 -81.555 231.050 ;
        RECT -80.435 230.880 -80.265 231.050 ;
        RECT -79.145 230.880 -78.975 231.050 ;
        RECT -77.855 230.880 -77.685 231.050 ;
        RECT -76.565 230.880 -76.395 231.050 ;
        RECT -75.275 230.880 -75.105 231.050 ;
        RECT -73.985 230.880 -73.815 231.050 ;
        RECT -72.695 230.880 -72.525 231.050 ;
        RECT -91.610 227.995 -78.120 230.325 ;
        RECT 682.310 258.595 682.480 258.765 ;
        RECT 699.610 258.645 699.780 258.815 ;
        RECT 717.400 258.685 717.570 258.855 ;
        RECT 734.660 258.715 734.830 258.885 ;
        RECT 752.130 258.705 752.300 258.875 ;
        RECT 679.490 257.095 679.660 257.265 ;
        RECT 679.850 257.095 680.020 257.265 ;
        RECT 680.710 257.095 680.880 257.265 ;
        RECT 681.070 257.095 681.240 257.265 ;
        RECT 681.430 257.095 681.600 257.265 ;
        RECT 681.790 257.095 681.960 257.265 ;
        RECT 682.150 257.095 682.320 257.265 ;
        RECT 682.510 257.095 682.680 257.265 ;
        RECT 682.870 257.095 683.040 257.265 ;
        RECT 683.950 257.095 684.120 257.265 ;
        RECT 684.310 257.095 684.480 257.265 ;
        RECT 696.770 257.105 696.940 257.275 ;
        RECT 697.130 257.105 697.300 257.275 ;
        RECT 697.990 257.105 698.160 257.275 ;
        RECT 698.350 257.105 698.520 257.275 ;
        RECT 698.710 257.105 698.880 257.275 ;
        RECT 699.070 257.105 699.240 257.275 ;
        RECT 699.430 257.105 699.600 257.275 ;
        RECT 699.790 257.105 699.960 257.275 ;
        RECT 700.150 257.105 700.320 257.275 ;
        RECT 701.230 257.105 701.400 257.275 ;
        RECT 701.590 257.105 701.760 257.275 ;
        RECT 714.540 257.105 714.710 257.275 ;
        RECT 714.900 257.105 715.070 257.275 ;
        RECT 715.760 257.105 715.930 257.275 ;
        RECT 716.120 257.105 716.290 257.275 ;
        RECT 716.480 257.105 716.650 257.275 ;
        RECT 716.840 257.105 717.010 257.275 ;
        RECT 717.200 257.105 717.370 257.275 ;
        RECT 717.560 257.105 717.730 257.275 ;
        RECT 717.920 257.105 718.090 257.275 ;
        RECT 719.000 257.105 719.170 257.275 ;
        RECT 719.360 257.105 719.530 257.275 ;
        RECT 731.780 257.105 731.950 257.275 ;
        RECT 732.140 257.105 732.310 257.275 ;
        RECT 733.000 257.105 733.170 257.275 ;
        RECT 733.360 257.105 733.530 257.275 ;
        RECT 733.720 257.105 733.890 257.275 ;
        RECT 734.080 257.105 734.250 257.275 ;
        RECT 734.440 257.105 734.610 257.275 ;
        RECT 734.800 257.105 734.970 257.275 ;
        RECT 735.160 257.105 735.330 257.275 ;
        RECT 736.240 257.105 736.410 257.275 ;
        RECT 736.600 257.105 736.770 257.275 ;
        RECT 749.260 257.115 749.430 257.285 ;
        RECT 749.620 257.115 749.790 257.285 ;
        RECT 750.480 257.115 750.650 257.285 ;
        RECT 750.840 257.115 751.010 257.285 ;
        RECT 751.200 257.115 751.370 257.285 ;
        RECT 751.560 257.115 751.730 257.285 ;
        RECT 751.920 257.115 752.090 257.285 ;
        RECT 752.280 257.115 752.450 257.285 ;
        RECT 752.640 257.115 752.810 257.285 ;
        RECT 753.720 257.115 753.890 257.285 ;
        RECT 754.080 257.115 754.250 257.285 ;
        RECT 679.525 256.615 679.695 256.785 ;
        RECT 680.005 256.615 680.175 256.785 ;
        RECT 680.485 256.615 680.655 256.785 ;
        RECT 680.965 256.615 681.135 256.785 ;
        RECT 681.445 256.615 681.615 256.785 ;
        RECT 681.925 256.615 682.095 256.785 ;
        RECT 682.405 256.615 682.575 256.785 ;
        RECT 682.885 256.615 683.055 256.785 ;
        RECT 683.365 256.615 683.535 256.785 ;
        RECT 683.845 256.615 684.015 256.785 ;
        RECT 684.325 256.615 684.495 256.785 ;
        RECT 696.805 256.625 696.975 256.795 ;
        RECT 697.285 256.625 697.455 256.795 ;
        RECT 697.765 256.625 697.935 256.795 ;
        RECT 698.245 256.625 698.415 256.795 ;
        RECT 698.725 256.625 698.895 256.795 ;
        RECT 699.205 256.625 699.375 256.795 ;
        RECT 699.685 256.625 699.855 256.795 ;
        RECT 700.165 256.625 700.335 256.795 ;
        RECT 700.645 256.625 700.815 256.795 ;
        RECT 701.125 256.625 701.295 256.795 ;
        RECT 701.605 256.625 701.775 256.795 ;
        RECT 714.575 256.625 714.745 256.795 ;
        RECT 715.055 256.625 715.225 256.795 ;
        RECT 715.535 256.625 715.705 256.795 ;
        RECT 716.015 256.625 716.185 256.795 ;
        RECT 716.495 256.625 716.665 256.795 ;
        RECT 716.975 256.625 717.145 256.795 ;
        RECT 717.455 256.625 717.625 256.795 ;
        RECT 717.935 256.625 718.105 256.795 ;
        RECT 718.415 256.625 718.585 256.795 ;
        RECT 718.895 256.625 719.065 256.795 ;
        RECT 719.375 256.625 719.545 256.795 ;
        RECT 731.815 256.625 731.985 256.795 ;
        RECT 732.295 256.625 732.465 256.795 ;
        RECT 732.775 256.625 732.945 256.795 ;
        RECT 733.255 256.625 733.425 256.795 ;
        RECT 733.735 256.625 733.905 256.795 ;
        RECT 734.215 256.625 734.385 256.795 ;
        RECT 734.695 256.625 734.865 256.795 ;
        RECT 735.175 256.625 735.345 256.795 ;
        RECT 735.655 256.625 735.825 256.795 ;
        RECT 736.135 256.625 736.305 256.795 ;
        RECT 736.615 256.625 736.785 256.795 ;
        RECT 749.295 256.635 749.465 256.805 ;
        RECT 749.775 256.635 749.945 256.805 ;
        RECT 750.255 256.635 750.425 256.805 ;
        RECT 750.735 256.635 750.905 256.805 ;
        RECT 751.215 256.635 751.385 256.805 ;
        RECT 751.695 256.635 751.865 256.805 ;
        RECT 752.175 256.635 752.345 256.805 ;
        RECT 752.655 256.635 752.825 256.805 ;
        RECT 753.135 256.635 753.305 256.805 ;
        RECT 753.615 256.635 753.785 256.805 ;
        RECT 754.095 256.635 754.265 256.805 ;
        RECT 857.565 255.775 857.735 255.945 ;
        RECT 857.925 255.775 858.095 255.945 ;
        RECT 858.285 255.775 858.455 255.945 ;
        RECT 856.035 255.295 856.205 255.465 ;
        RECT 856.515 255.295 856.685 255.465 ;
        RECT 856.995 255.295 857.165 255.465 ;
        RECT 857.475 255.295 857.645 255.465 ;
        RECT 857.955 255.295 858.125 255.465 ;
        RECT 858.435 255.295 858.605 255.465 ;
        RECT 858.915 255.295 859.085 255.465 ;
        RECT 634.950 254.005 635.120 254.175 ;
        RECT 635.310 254.005 635.480 254.175 ;
        RECT 639.140 254.095 639.310 254.265 ;
        RECT 639.500 254.095 639.670 254.265 ;
        RECT 643.240 254.075 643.410 254.245 ;
        RECT 643.600 254.075 643.770 254.245 ;
        RECT 595.730 253.555 595.900 253.725 ;
        RECT 596.090 253.555 596.260 253.725 ;
        RECT 595.095 253.075 595.265 253.245 ;
        RECT 595.575 253.075 595.745 253.245 ;
        RECT 596.055 253.075 596.225 253.245 ;
        RECT 596.200 252.355 596.370 252.525 ;
        RECT 596.560 252.355 596.730 252.525 ;
        RECT 605.065 249.345 605.595 252.755 ;
        RECT 634.985 253.525 635.155 253.695 ;
        RECT 635.465 253.525 635.635 253.695 ;
        RECT 635.945 253.525 636.115 253.695 ;
        RECT 639.175 253.615 639.345 253.785 ;
        RECT 639.655 253.615 639.825 253.785 ;
        RECT 640.135 253.615 640.305 253.785 ;
        RECT 643.275 253.595 643.445 253.765 ;
        RECT 643.755 253.595 643.925 253.765 ;
        RECT 644.235 253.595 644.405 253.765 ;
        RECT 751.645 253.190 751.815 253.360 ;
        RECT 861.290 253.285 861.460 253.455 ;
        RECT 861.650 253.285 861.820 253.455 ;
        RECT 862.010 253.285 862.180 253.455 ;
        RECT 625.470 252.685 625.640 252.855 ;
        RECT 681.865 252.980 682.035 253.150 ;
        RECT 863.260 253.285 863.430 253.455 ;
        RECT 863.620 253.285 863.790 253.455 ;
        RECT 760.295 252.800 760.465 252.970 ;
        RECT 861.345 252.805 861.515 252.975 ;
        RECT 861.825 252.805 861.995 252.975 ;
        RECT 862.305 252.805 862.475 252.975 ;
        RECT 862.785 252.805 862.955 252.975 ;
        RECT 863.265 252.805 863.435 252.975 ;
        RECT 863.745 252.805 863.915 252.975 ;
        RECT 864.225 252.805 864.395 252.975 ;
        RECT 625.470 252.325 625.640 252.495 ;
        RECT 625.470 251.965 625.640 252.135 ;
        RECT 625.470 251.605 625.640 251.775 ;
        RECT 625.470 251.245 625.640 251.415 ;
        RECT 679.900 251.435 680.070 251.605 ;
        RECT 680.260 251.435 680.430 251.605 ;
        RECT 681.120 251.435 681.290 251.605 ;
        RECT 681.480 251.435 681.650 251.605 ;
        RECT 681.840 251.435 682.010 251.605 ;
        RECT 682.200 251.435 682.370 251.605 ;
        RECT 682.560 251.435 682.730 251.605 ;
        RECT 682.920 251.435 683.090 251.605 ;
        RECT 683.280 251.435 683.450 251.605 ;
        RECT 684.360 251.435 684.530 251.605 ;
        RECT 684.720 251.435 684.890 251.605 ;
        RECT 687.140 251.395 687.310 251.565 ;
        RECT 687.500 251.395 687.670 251.565 ;
        RECT 688.360 251.395 688.530 251.565 ;
        RECT 688.720 251.395 688.890 251.565 ;
        RECT 689.080 251.395 689.250 251.565 ;
        RECT 689.440 251.395 689.610 251.565 ;
        RECT 689.800 251.395 689.970 251.565 ;
        RECT 690.160 251.395 690.330 251.565 ;
        RECT 690.520 251.395 690.690 251.565 ;
        RECT 691.600 251.395 691.770 251.565 ;
        RECT 691.960 251.395 692.130 251.565 ;
        RECT 697.130 251.455 697.300 251.625 ;
        RECT 697.490 251.455 697.660 251.625 ;
        RECT 698.350 251.455 698.520 251.625 ;
        RECT 698.710 251.455 698.880 251.625 ;
        RECT 699.070 251.455 699.240 251.625 ;
        RECT 699.430 251.455 699.600 251.625 ;
        RECT 699.790 251.455 699.960 251.625 ;
        RECT 700.150 251.455 700.320 251.625 ;
        RECT 700.510 251.455 700.680 251.625 ;
        RECT 701.590 251.455 701.760 251.625 ;
        RECT 701.950 251.455 702.120 251.625 ;
        RECT 704.370 251.415 704.540 251.585 ;
        RECT 704.730 251.415 704.900 251.585 ;
        RECT 705.590 251.415 705.760 251.585 ;
        RECT 705.950 251.415 706.120 251.585 ;
        RECT 706.310 251.415 706.480 251.585 ;
        RECT 706.670 251.415 706.840 251.585 ;
        RECT 707.030 251.415 707.200 251.585 ;
        RECT 707.390 251.415 707.560 251.585 ;
        RECT 707.750 251.415 707.920 251.585 ;
        RECT 708.830 251.415 709.000 251.585 ;
        RECT 709.190 251.415 709.360 251.585 ;
        RECT 714.700 251.555 714.870 251.725 ;
        RECT 715.060 251.555 715.230 251.725 ;
        RECT 715.920 251.555 716.090 251.725 ;
        RECT 716.280 251.555 716.450 251.725 ;
        RECT 716.640 251.555 716.810 251.725 ;
        RECT 717.000 251.555 717.170 251.725 ;
        RECT 717.360 251.555 717.530 251.725 ;
        RECT 717.720 251.555 717.890 251.725 ;
        RECT 718.080 251.555 718.250 251.725 ;
        RECT 719.160 251.555 719.330 251.725 ;
        RECT 719.520 251.555 719.690 251.725 ;
        RECT 721.940 251.515 722.110 251.685 ;
        RECT 722.300 251.515 722.470 251.685 ;
        RECT 723.160 251.515 723.330 251.685 ;
        RECT 723.520 251.515 723.690 251.685 ;
        RECT 723.880 251.515 724.050 251.685 ;
        RECT 724.240 251.515 724.410 251.685 ;
        RECT 724.600 251.515 724.770 251.685 ;
        RECT 724.960 251.515 725.130 251.685 ;
        RECT 725.320 251.515 725.490 251.685 ;
        RECT 726.400 251.515 726.570 251.685 ;
        RECT 726.760 251.515 726.930 251.685 ;
        RECT 731.870 251.585 732.040 251.755 ;
        RECT 732.230 251.585 732.400 251.755 ;
        RECT 733.090 251.585 733.260 251.755 ;
        RECT 733.450 251.585 733.620 251.755 ;
        RECT 733.810 251.585 733.980 251.755 ;
        RECT 734.170 251.585 734.340 251.755 ;
        RECT 734.530 251.585 734.700 251.755 ;
        RECT 734.890 251.585 735.060 251.755 ;
        RECT 735.250 251.585 735.420 251.755 ;
        RECT 736.330 251.585 736.500 251.755 ;
        RECT 736.690 251.585 736.860 251.755 ;
        RECT 739.110 251.545 739.280 251.715 ;
        RECT 739.470 251.545 739.640 251.715 ;
        RECT 740.330 251.545 740.500 251.715 ;
        RECT 740.690 251.545 740.860 251.715 ;
        RECT 741.050 251.545 741.220 251.715 ;
        RECT 741.410 251.545 741.580 251.715 ;
        RECT 741.770 251.545 741.940 251.715 ;
        RECT 742.130 251.545 742.300 251.715 ;
        RECT 742.490 251.545 742.660 251.715 ;
        RECT 743.570 251.545 743.740 251.715 ;
        RECT 743.930 251.545 744.100 251.715 ;
        RECT 749.680 251.645 749.850 251.815 ;
        RECT 750.040 251.645 750.210 251.815 ;
        RECT 750.900 251.645 751.070 251.815 ;
        RECT 751.260 251.645 751.430 251.815 ;
        RECT 751.620 251.645 751.790 251.815 ;
        RECT 751.980 251.645 752.150 251.815 ;
        RECT 752.340 251.645 752.510 251.815 ;
        RECT 752.700 251.645 752.870 251.815 ;
        RECT 753.060 251.645 753.230 251.815 ;
        RECT 754.140 251.645 754.310 251.815 ;
        RECT 754.500 251.645 754.670 251.815 ;
        RECT 756.920 251.605 757.090 251.775 ;
        RECT 757.280 251.605 757.450 251.775 ;
        RECT 758.140 251.605 758.310 251.775 ;
        RECT 758.500 251.605 758.670 251.775 ;
        RECT 758.860 251.605 759.030 251.775 ;
        RECT 759.220 251.605 759.390 251.775 ;
        RECT 759.580 251.605 759.750 251.775 ;
        RECT 759.940 251.605 760.110 251.775 ;
        RECT 760.300 251.605 760.470 251.775 ;
        RECT 761.380 251.605 761.550 251.775 ;
        RECT 761.740 251.605 761.910 251.775 ;
        RECT 614.590 250.875 614.760 251.045 ;
        RECT 616.170 250.875 616.340 251.045 ;
        RECT 625.470 250.885 625.640 251.055 ;
        RECT 679.935 250.955 680.105 251.125 ;
        RECT 680.415 250.955 680.585 251.125 ;
        RECT 680.895 250.955 681.065 251.125 ;
        RECT 681.375 250.955 681.545 251.125 ;
        RECT 681.855 250.955 682.025 251.125 ;
        RECT 682.335 250.955 682.505 251.125 ;
        RECT 682.815 250.955 682.985 251.125 ;
        RECT 683.295 250.955 683.465 251.125 ;
        RECT 683.775 250.955 683.945 251.125 ;
        RECT 684.255 250.955 684.425 251.125 ;
        RECT 684.735 250.955 684.905 251.125 ;
        RECT 687.175 250.915 687.345 251.085 ;
        RECT 687.655 250.915 687.825 251.085 ;
        RECT 688.135 250.915 688.305 251.085 ;
        RECT 688.615 250.915 688.785 251.085 ;
        RECT 689.095 250.915 689.265 251.085 ;
        RECT 689.575 250.915 689.745 251.085 ;
        RECT 690.055 250.915 690.225 251.085 ;
        RECT 690.535 250.915 690.705 251.085 ;
        RECT 691.015 250.915 691.185 251.085 ;
        RECT 691.495 250.915 691.665 251.085 ;
        RECT 691.975 250.915 692.145 251.085 ;
        RECT 697.165 250.975 697.335 251.145 ;
        RECT 697.645 250.975 697.815 251.145 ;
        RECT 698.125 250.975 698.295 251.145 ;
        RECT 698.605 250.975 698.775 251.145 ;
        RECT 699.085 250.975 699.255 251.145 ;
        RECT 699.565 250.975 699.735 251.145 ;
        RECT 700.045 250.975 700.215 251.145 ;
        RECT 700.525 250.975 700.695 251.145 ;
        RECT 701.005 250.975 701.175 251.145 ;
        RECT 701.485 250.975 701.655 251.145 ;
        RECT 701.965 250.975 702.135 251.145 ;
        RECT 704.405 250.935 704.575 251.105 ;
        RECT 704.885 250.935 705.055 251.105 ;
        RECT 705.365 250.935 705.535 251.105 ;
        RECT 705.845 250.935 706.015 251.105 ;
        RECT 706.325 250.935 706.495 251.105 ;
        RECT 706.805 250.935 706.975 251.105 ;
        RECT 707.285 250.935 707.455 251.105 ;
        RECT 707.765 250.935 707.935 251.105 ;
        RECT 708.245 250.935 708.415 251.105 ;
        RECT 708.725 250.935 708.895 251.105 ;
        RECT 709.205 250.935 709.375 251.105 ;
        RECT 714.735 251.075 714.905 251.245 ;
        RECT 715.215 251.075 715.385 251.245 ;
        RECT 715.695 251.075 715.865 251.245 ;
        RECT 716.175 251.075 716.345 251.245 ;
        RECT 716.655 251.075 716.825 251.245 ;
        RECT 717.135 251.075 717.305 251.245 ;
        RECT 717.615 251.075 717.785 251.245 ;
        RECT 718.095 251.075 718.265 251.245 ;
        RECT 718.575 251.075 718.745 251.245 ;
        RECT 719.055 251.075 719.225 251.245 ;
        RECT 719.535 251.075 719.705 251.245 ;
        RECT 721.975 251.035 722.145 251.205 ;
        RECT 722.455 251.035 722.625 251.205 ;
        RECT 722.935 251.035 723.105 251.205 ;
        RECT 723.415 251.035 723.585 251.205 ;
        RECT 723.895 251.035 724.065 251.205 ;
        RECT 724.375 251.035 724.545 251.205 ;
        RECT 724.855 251.035 725.025 251.205 ;
        RECT 725.335 251.035 725.505 251.205 ;
        RECT 725.815 251.035 725.985 251.205 ;
        RECT 726.295 251.035 726.465 251.205 ;
        RECT 726.775 251.035 726.945 251.205 ;
        RECT 731.905 251.105 732.075 251.275 ;
        RECT 732.385 251.105 732.555 251.275 ;
        RECT 732.865 251.105 733.035 251.275 ;
        RECT 733.345 251.105 733.515 251.275 ;
        RECT 733.825 251.105 733.995 251.275 ;
        RECT 734.305 251.105 734.475 251.275 ;
        RECT 734.785 251.105 734.955 251.275 ;
        RECT 735.265 251.105 735.435 251.275 ;
        RECT 735.745 251.105 735.915 251.275 ;
        RECT 736.225 251.105 736.395 251.275 ;
        RECT 736.705 251.105 736.875 251.275 ;
        RECT 739.145 251.065 739.315 251.235 ;
        RECT 739.625 251.065 739.795 251.235 ;
        RECT 740.105 251.065 740.275 251.235 ;
        RECT 740.585 251.065 740.755 251.235 ;
        RECT 741.065 251.065 741.235 251.235 ;
        RECT 741.545 251.065 741.715 251.235 ;
        RECT 742.025 251.065 742.195 251.235 ;
        RECT 742.505 251.065 742.675 251.235 ;
        RECT 742.985 251.065 743.155 251.235 ;
        RECT 743.465 251.065 743.635 251.235 ;
        RECT 743.945 251.065 744.115 251.235 ;
        RECT 749.715 251.165 749.885 251.335 ;
        RECT 750.195 251.165 750.365 251.335 ;
        RECT 750.675 251.165 750.845 251.335 ;
        RECT 751.155 251.165 751.325 251.335 ;
        RECT 751.635 251.165 751.805 251.335 ;
        RECT 752.115 251.165 752.285 251.335 ;
        RECT 752.595 251.165 752.765 251.335 ;
        RECT 753.075 251.165 753.245 251.335 ;
        RECT 753.555 251.165 753.725 251.335 ;
        RECT 754.035 251.165 754.205 251.335 ;
        RECT 754.515 251.165 754.685 251.335 ;
        RECT 756.955 251.125 757.125 251.295 ;
        RECT 757.435 251.125 757.605 251.295 ;
        RECT 757.915 251.125 758.085 251.295 ;
        RECT 758.395 251.125 758.565 251.295 ;
        RECT 758.875 251.125 759.045 251.295 ;
        RECT 759.355 251.125 759.525 251.295 ;
        RECT 759.835 251.125 760.005 251.295 ;
        RECT 760.315 251.125 760.485 251.295 ;
        RECT 760.795 251.125 760.965 251.295 ;
        RECT 761.275 251.125 761.445 251.295 ;
        RECT 761.755 251.125 761.925 251.295 ;
        RECT 625.470 250.525 625.640 250.695 ;
        RECT 625.470 250.165 625.640 250.335 ;
        RECT 625.470 249.805 625.640 249.975 ;
        RECT 639.940 249.985 640.110 250.155 ;
        RECT 643.990 250.035 644.160 250.205 ;
        RECT 857.625 250.005 857.795 250.175 ;
        RECT 857.985 250.005 858.155 250.175 ;
        RECT 858.345 250.005 858.515 250.175 ;
        RECT 614.590 249.405 614.760 249.575 ;
        RECT 616.170 249.405 616.340 249.575 ;
        RECT 856.095 249.525 856.265 249.695 ;
        RECT 856.575 249.525 856.745 249.695 ;
        RECT 857.055 249.525 857.225 249.695 ;
        RECT 857.535 249.525 857.705 249.695 ;
        RECT 858.015 249.525 858.185 249.695 ;
        RECT 858.495 249.525 858.665 249.695 ;
        RECT 858.975 249.525 859.145 249.695 ;
        RECT 601.830 248.515 602.000 248.685 ;
        RECT 602.190 248.515 602.360 248.685 ;
        RECT 591.520 247.115 591.690 247.285 ;
        RECT 591.520 246.755 591.690 246.925 ;
        RECT 591.520 246.395 591.690 246.565 ;
        RECT 680.125 246.810 680.295 246.980 ;
        RECT 749.905 247.020 750.075 247.190 ;
        RECT 591.520 246.035 591.690 246.205 ;
        RECT 591.520 245.675 591.690 245.845 ;
        RECT 681.585 245.755 681.755 245.925 ;
        RECT 681.945 245.755 682.115 245.925 ;
        RECT 682.305 245.755 682.475 245.925 ;
        RECT 687.245 245.765 687.415 245.935 ;
        RECT 687.605 245.765 687.775 245.935 ;
        RECT 687.965 245.765 688.135 245.935 ;
        RECT 691.010 245.785 691.180 245.955 ;
        RECT 691.370 245.785 691.540 245.955 ;
        RECT 691.730 245.785 691.900 245.955 ;
        RECT 692.980 245.785 693.150 245.955 ;
        RECT 693.340 245.785 693.510 245.955 ;
        RECT 698.815 245.775 698.985 245.945 ;
        RECT 699.175 245.775 699.345 245.945 ;
        RECT 699.535 245.775 699.705 245.945 ;
        RECT 704.475 245.785 704.645 245.955 ;
        RECT 704.835 245.785 705.005 245.955 ;
        RECT 705.195 245.785 705.365 245.955 ;
        RECT 708.240 245.805 708.410 245.975 ;
        RECT 708.600 245.805 708.770 245.975 ;
        RECT 708.960 245.805 709.130 245.975 ;
        RECT 710.210 245.805 710.380 245.975 ;
        RECT 710.570 245.805 710.740 245.975 ;
        RECT 716.385 245.875 716.555 246.045 ;
        RECT 716.745 245.875 716.915 246.045 ;
        RECT 717.105 245.875 717.275 246.045 ;
        RECT 722.045 245.885 722.215 246.055 ;
        RECT 722.405 245.885 722.575 246.055 ;
        RECT 722.765 245.885 722.935 246.055 ;
        RECT 725.810 245.905 725.980 246.075 ;
        RECT 726.170 245.905 726.340 246.075 ;
        RECT 726.530 245.905 726.700 246.075 ;
        RECT 727.780 245.905 727.950 246.075 ;
        RECT 728.140 245.905 728.310 246.075 ;
        RECT 733.555 245.905 733.725 246.075 ;
        RECT 733.915 245.905 734.085 246.075 ;
        RECT 734.275 245.905 734.445 246.075 ;
        RECT 739.215 245.915 739.385 246.085 ;
        RECT 739.575 245.915 739.745 246.085 ;
        RECT 739.935 245.915 740.105 246.085 ;
        RECT 742.980 245.935 743.150 246.105 ;
        RECT 743.340 245.935 743.510 246.105 ;
        RECT 743.700 245.935 743.870 246.105 ;
        RECT 756.535 246.915 756.705 247.085 ;
        RECT 744.950 245.935 745.120 246.105 ;
        RECT 745.310 245.935 745.480 246.105 ;
        RECT 756.535 246.555 756.705 246.725 ;
        RECT 751.365 245.965 751.535 246.135 ;
        RECT 751.725 245.965 751.895 246.135 ;
        RECT 752.085 245.965 752.255 246.135 ;
        RECT 757.025 245.975 757.195 246.145 ;
        RECT 757.385 245.975 757.555 246.145 ;
        RECT 757.745 245.975 757.915 246.145 ;
        RECT 760.790 245.995 760.960 246.165 ;
        RECT 761.150 245.995 761.320 246.165 ;
        RECT 761.510 245.995 761.680 246.165 ;
        RECT 762.760 245.995 762.930 246.165 ;
        RECT 763.120 245.995 763.290 246.165 ;
        RECT 591.520 245.315 591.690 245.485 ;
        RECT 680.055 245.275 680.225 245.445 ;
        RECT 680.535 245.275 680.705 245.445 ;
        RECT 681.015 245.275 681.185 245.445 ;
        RECT 681.495 245.275 681.665 245.445 ;
        RECT 681.975 245.275 682.145 245.445 ;
        RECT 682.455 245.275 682.625 245.445 ;
        RECT 682.935 245.275 683.105 245.445 ;
        RECT 685.715 245.285 685.885 245.455 ;
        RECT 686.195 245.285 686.365 245.455 ;
        RECT 686.675 245.285 686.845 245.455 ;
        RECT 687.155 245.285 687.325 245.455 ;
        RECT 687.635 245.285 687.805 245.455 ;
        RECT 688.115 245.285 688.285 245.455 ;
        RECT 688.595 245.285 688.765 245.455 ;
        RECT 691.065 245.305 691.235 245.475 ;
        RECT 691.545 245.305 691.715 245.475 ;
        RECT 692.025 245.305 692.195 245.475 ;
        RECT 692.505 245.305 692.675 245.475 ;
        RECT 692.985 245.305 693.155 245.475 ;
        RECT 693.465 245.305 693.635 245.475 ;
        RECT 693.945 245.305 694.115 245.475 ;
        RECT 697.285 245.295 697.455 245.465 ;
        RECT 697.765 245.295 697.935 245.465 ;
        RECT 698.245 245.295 698.415 245.465 ;
        RECT 698.725 245.295 698.895 245.465 ;
        RECT 699.205 245.295 699.375 245.465 ;
        RECT 699.685 245.295 699.855 245.465 ;
        RECT 700.165 245.295 700.335 245.465 ;
        RECT 702.945 245.305 703.115 245.475 ;
        RECT 703.425 245.305 703.595 245.475 ;
        RECT 703.905 245.305 704.075 245.475 ;
        RECT 704.385 245.305 704.555 245.475 ;
        RECT 704.865 245.305 705.035 245.475 ;
        RECT 705.345 245.305 705.515 245.475 ;
        RECT 705.825 245.305 705.995 245.475 ;
        RECT 708.295 245.325 708.465 245.495 ;
        RECT 708.775 245.325 708.945 245.495 ;
        RECT 709.255 245.325 709.425 245.495 ;
        RECT 709.735 245.325 709.905 245.495 ;
        RECT 710.215 245.325 710.385 245.495 ;
        RECT 710.695 245.325 710.865 245.495 ;
        RECT 711.175 245.325 711.345 245.495 ;
        RECT 714.855 245.395 715.025 245.565 ;
        RECT 715.335 245.395 715.505 245.565 ;
        RECT 715.815 245.395 715.985 245.565 ;
        RECT 716.295 245.395 716.465 245.565 ;
        RECT 716.775 245.395 716.945 245.565 ;
        RECT 717.255 245.395 717.425 245.565 ;
        RECT 717.735 245.395 717.905 245.565 ;
        RECT 720.515 245.405 720.685 245.575 ;
        RECT 720.995 245.405 721.165 245.575 ;
        RECT 721.475 245.405 721.645 245.575 ;
        RECT 721.955 245.405 722.125 245.575 ;
        RECT 722.435 245.405 722.605 245.575 ;
        RECT 722.915 245.405 723.085 245.575 ;
        RECT 723.395 245.405 723.565 245.575 ;
        RECT 725.865 245.425 726.035 245.595 ;
        RECT 726.345 245.425 726.515 245.595 ;
        RECT 726.825 245.425 726.995 245.595 ;
        RECT 727.305 245.425 727.475 245.595 ;
        RECT 727.785 245.425 727.955 245.595 ;
        RECT 728.265 245.425 728.435 245.595 ;
        RECT 728.745 245.425 728.915 245.595 ;
        RECT 732.025 245.425 732.195 245.595 ;
        RECT 732.505 245.425 732.675 245.595 ;
        RECT 732.985 245.425 733.155 245.595 ;
        RECT 733.465 245.425 733.635 245.595 ;
        RECT 733.945 245.425 734.115 245.595 ;
        RECT 734.425 245.425 734.595 245.595 ;
        RECT 734.905 245.425 735.075 245.595 ;
        RECT 737.685 245.435 737.855 245.605 ;
        RECT 738.165 245.435 738.335 245.605 ;
        RECT 738.645 245.435 738.815 245.605 ;
        RECT 739.125 245.435 739.295 245.605 ;
        RECT 739.605 245.435 739.775 245.605 ;
        RECT 740.085 245.435 740.255 245.605 ;
        RECT 740.565 245.435 740.735 245.605 ;
        RECT 743.035 245.455 743.205 245.625 ;
        RECT 743.515 245.455 743.685 245.625 ;
        RECT 743.995 245.455 744.165 245.625 ;
        RECT 744.475 245.455 744.645 245.625 ;
        RECT 744.955 245.455 745.125 245.625 ;
        RECT 745.435 245.455 745.605 245.625 ;
        RECT 745.915 245.455 746.085 245.625 ;
        RECT 749.835 245.485 750.005 245.655 ;
        RECT 750.315 245.485 750.485 245.655 ;
        RECT 750.795 245.485 750.965 245.655 ;
        RECT 751.275 245.485 751.445 245.655 ;
        RECT 751.755 245.485 751.925 245.655 ;
        RECT 752.235 245.485 752.405 245.655 ;
        RECT 752.715 245.485 752.885 245.655 ;
        RECT 755.495 245.495 755.665 245.665 ;
        RECT 755.975 245.495 756.145 245.665 ;
        RECT 756.455 245.495 756.625 245.665 ;
        RECT 756.935 245.495 757.105 245.665 ;
        RECT 757.415 245.495 757.585 245.665 ;
        RECT 757.895 245.495 758.065 245.665 ;
        RECT 758.375 245.495 758.545 245.665 ;
        RECT 760.845 245.515 761.015 245.685 ;
        RECT 761.325 245.515 761.495 245.685 ;
        RECT 761.805 245.515 761.975 245.685 ;
        RECT 762.285 245.515 762.455 245.685 ;
        RECT 762.765 245.515 762.935 245.685 ;
        RECT 763.245 245.515 763.415 245.685 ;
        RECT 763.725 245.515 763.895 245.685 ;
        RECT 122.030 223.575 125.800 224.825 ;
        RECT -97.160 222.095 -96.990 222.265 ;
        RECT -97.160 221.735 -96.990 221.905 ;
        RECT -97.160 221.375 -96.990 221.545 ;
        RECT -97.160 221.015 -96.990 221.185 ;
        RECT -94.580 222.095 -94.410 222.265 ;
        RECT -94.580 221.735 -94.410 221.905 ;
        RECT -94.580 221.375 -94.410 221.545 ;
        RECT -94.580 221.015 -94.410 221.185 ;
        RECT -92.000 222.095 -91.830 222.265 ;
        RECT -92.000 221.735 -91.830 221.905 ;
        RECT -92.000 221.375 -91.830 221.545 ;
        RECT -92.000 221.015 -91.830 221.185 ;
        RECT -89.420 222.095 -89.250 222.265 ;
        RECT -89.420 221.735 -89.250 221.905 ;
        RECT -89.420 221.375 -89.250 221.545 ;
        RECT -89.420 221.015 -89.250 221.185 ;
        RECT -86.840 222.095 -86.670 222.265 ;
        RECT -86.840 221.735 -86.670 221.905 ;
        RECT -86.840 221.375 -86.670 221.545 ;
        RECT -86.840 221.015 -86.670 221.185 ;
        RECT -84.260 222.095 -84.090 222.265 ;
        RECT -84.260 221.735 -84.090 221.905 ;
        RECT -84.260 221.375 -84.090 221.545 ;
        RECT -84.260 221.015 -84.090 221.185 ;
        RECT -81.680 222.095 -81.510 222.265 ;
        RECT -81.680 221.735 -81.510 221.905 ;
        RECT -81.680 221.375 -81.510 221.545 ;
        RECT -81.680 221.015 -81.510 221.185 ;
        RECT -79.100 222.095 -78.930 222.265 ;
        RECT -79.100 221.735 -78.930 221.905 ;
        RECT -79.100 221.375 -78.930 221.545 ;
        RECT -79.100 221.015 -78.930 221.185 ;
        RECT -76.520 222.095 -76.350 222.265 ;
        RECT -76.520 221.735 -76.350 221.905 ;
        RECT -76.520 221.375 -76.350 221.545 ;
        RECT -76.520 221.015 -76.350 221.185 ;
        RECT -73.940 222.095 -73.770 222.265 ;
        RECT -73.940 221.735 -73.770 221.905 ;
        RECT -73.940 221.375 -73.770 221.545 ;
        RECT -73.940 221.015 -73.770 221.185 ;
        RECT -71.360 222.095 -71.190 222.265 ;
        RECT -71.360 221.735 -71.190 221.905 ;
        RECT -71.360 221.375 -71.190 221.545 ;
        RECT -71.360 221.015 -71.190 221.185 ;
        RECT 197.090 222.225 208.420 224.915 ;
        RECT -96.515 218.780 -96.345 218.950 ;
        RECT -95.225 218.780 -95.055 218.950 ;
        RECT -93.935 218.780 -93.765 218.950 ;
        RECT -92.645 218.780 -92.475 218.950 ;
        RECT -91.355 218.780 -91.185 218.950 ;
        RECT -90.065 218.780 -89.895 218.950 ;
        RECT -88.775 218.780 -88.605 218.950 ;
        RECT -87.485 218.780 -87.315 218.950 ;
        RECT -86.195 218.780 -86.025 218.950 ;
        RECT -84.905 218.780 -84.735 218.950 ;
        RECT -83.615 218.780 -83.445 218.950 ;
        RECT -82.325 218.780 -82.155 218.950 ;
        RECT -81.035 218.780 -80.865 218.950 ;
        RECT -79.745 218.780 -79.575 218.950 ;
        RECT -78.455 218.780 -78.285 218.950 ;
        RECT -77.165 218.780 -76.995 218.950 ;
        RECT -75.875 218.780 -75.705 218.950 ;
        RECT -74.585 218.780 -74.415 218.950 ;
        RECT -73.295 218.780 -73.125 218.950 ;
        RECT -72.005 218.780 -71.835 218.950 ;
        RECT -90.980 215.875 -77.490 218.205 ;
        RECT 55.460 218.300 55.630 218.470 ;
        RECT 55.820 218.300 55.990 218.470 ;
        RECT 248.275 218.755 249.165 219.285 ;
        RECT 342.200 219.330 342.370 219.500 ;
        RECT 342.560 219.330 342.730 219.500 ;
        RECT 342.920 219.330 343.090 219.500 ;
        RECT 343.280 219.330 343.450 219.500 ;
        RECT 343.640 219.330 343.810 219.500 ;
        RECT 344.000 219.330 344.170 219.500 ;
        RECT 319.320 217.500 320.570 218.030 ;
        RECT 9.790 214.985 9.960 215.155 ;
        RECT 9.790 214.625 9.960 214.795 ;
        RECT 15.080 214.985 15.250 215.155 ;
        RECT 20.370 214.985 20.540 215.155 ;
        RECT 25.660 214.985 25.830 215.155 ;
        RECT 30.950 214.985 31.120 215.155 ;
        RECT 9.790 214.265 9.960 214.435 ;
        RECT 9.790 213.905 9.960 214.075 ;
        RECT 9.790 209.515 9.960 209.685 ;
        RECT 9.790 209.155 9.960 209.325 ;
        RECT 9.790 208.795 9.960 208.965 ;
        RECT 9.790 208.435 9.960 208.605 ;
        RECT 6.780 207.395 6.950 207.565 ;
        RECT 6.780 207.035 6.950 207.205 ;
        RECT 6.780 206.675 6.950 206.845 ;
        RECT 6.780 206.315 6.950 206.485 ;
        RECT 6.780 205.955 6.950 206.125 ;
        RECT 6.780 205.595 6.950 205.765 ;
        RECT 6.780 205.235 6.950 205.405 ;
        RECT 6.780 204.875 6.950 205.045 ;
        RECT 6.780 204.515 6.950 204.685 ;
        RECT 6.780 204.155 6.950 204.325 ;
        RECT 6.780 203.795 6.950 203.965 ;
        RECT 6.780 203.435 6.950 203.605 ;
        RECT 6.780 203.075 6.950 203.245 ;
        RECT 6.780 202.715 6.950 202.885 ;
        RECT 6.780 202.355 6.950 202.525 ;
        RECT 6.780 201.995 6.950 202.165 ;
        RECT 6.780 201.635 6.950 201.805 ;
        RECT 9.790 204.045 9.960 204.215 ;
        RECT 9.790 203.685 9.960 203.855 ;
        RECT 9.790 203.325 9.960 203.495 ;
        RECT 9.790 202.965 9.960 203.135 ;
        RECT 9.790 198.575 9.960 198.745 ;
        RECT 9.790 198.215 9.960 198.385 ;
        RECT 9.790 197.855 9.960 198.025 ;
        RECT 9.790 197.495 9.960 197.665 ;
        RECT 9.790 193.105 9.960 193.275 ;
        RECT 15.080 214.625 15.250 214.795 ;
        RECT 15.080 214.265 15.250 214.435 ;
        RECT 15.080 213.905 15.250 214.075 ;
        RECT 15.080 209.515 15.250 209.685 ;
        RECT 15.080 209.155 15.250 209.325 ;
        RECT 15.080 208.795 15.250 208.965 ;
        RECT 15.080 208.435 15.250 208.605 ;
        RECT 15.080 204.045 15.250 204.215 ;
        RECT 15.080 203.685 15.250 203.855 ;
        RECT 15.080 203.325 15.250 203.495 ;
        RECT 15.080 202.965 15.250 203.135 ;
        RECT 15.080 198.575 15.250 198.745 ;
        RECT 15.080 198.215 15.250 198.385 ;
        RECT 15.080 197.855 15.250 198.025 ;
        RECT 15.080 197.495 15.250 197.665 ;
        RECT 15.080 193.105 15.250 193.275 ;
        RECT 20.370 214.625 20.540 214.795 ;
        RECT 20.370 214.265 20.540 214.435 ;
        RECT 20.370 213.905 20.540 214.075 ;
        RECT 20.370 209.515 20.540 209.685 ;
        RECT 20.370 209.155 20.540 209.325 ;
        RECT 20.370 208.795 20.540 208.965 ;
        RECT 20.370 208.435 20.540 208.605 ;
        RECT 20.370 204.045 20.540 204.215 ;
        RECT 20.370 203.685 20.540 203.855 ;
        RECT 20.370 203.325 20.540 203.495 ;
        RECT 20.370 202.965 20.540 203.135 ;
        RECT 20.370 198.575 20.540 198.745 ;
        RECT 20.370 198.215 20.540 198.385 ;
        RECT 20.370 197.855 20.540 198.025 ;
        RECT 20.370 197.495 20.540 197.665 ;
        RECT 20.370 193.105 20.540 193.275 ;
        RECT 36.240 214.985 36.410 215.155 ;
        RECT 25.660 214.625 25.830 214.795 ;
        RECT 25.660 214.265 25.830 214.435 ;
        RECT 25.660 213.905 25.830 214.075 ;
        RECT 25.660 209.515 25.830 209.685 ;
        RECT 25.660 209.155 25.830 209.325 ;
        RECT 25.660 208.795 25.830 208.965 ;
        RECT 25.660 208.435 25.830 208.605 ;
        RECT 25.660 204.045 25.830 204.215 ;
        RECT 25.660 203.685 25.830 203.855 ;
        RECT 25.660 203.325 25.830 203.495 ;
        RECT 25.660 202.965 25.830 203.135 ;
        RECT 25.660 198.575 25.830 198.745 ;
        RECT 25.660 198.215 25.830 198.385 ;
        RECT 25.660 197.855 25.830 198.025 ;
        RECT 25.660 197.495 25.830 197.665 ;
        RECT 25.660 193.105 25.830 193.275 ;
        RECT 30.950 214.625 31.120 214.795 ;
        RECT 30.950 214.265 31.120 214.435 ;
        RECT 30.950 213.905 31.120 214.075 ;
        RECT 30.950 209.515 31.120 209.685 ;
        RECT 30.950 209.155 31.120 209.325 ;
        RECT 30.950 208.795 31.120 208.965 ;
        RECT 30.950 208.435 31.120 208.605 ;
        RECT 30.950 204.045 31.120 204.215 ;
        RECT 30.950 203.685 31.120 203.855 ;
        RECT 30.950 203.325 31.120 203.495 ;
        RECT 30.950 202.965 31.120 203.135 ;
        RECT 30.950 198.575 31.120 198.745 ;
        RECT 30.950 198.215 31.120 198.385 ;
        RECT 30.950 197.855 31.120 198.025 ;
        RECT 30.950 197.495 31.120 197.665 ;
        RECT 9.790 192.745 9.960 192.915 ;
        RECT 9.790 192.385 9.960 192.555 ;
        RECT 15.080 192.745 15.250 192.915 ;
        RECT 9.790 192.025 9.960 192.195 ;
        RECT 15.080 192.385 15.250 192.555 ;
        RECT 20.370 192.745 20.540 192.915 ;
        RECT 15.080 192.025 15.250 192.195 ;
        RECT 20.370 192.385 20.540 192.555 ;
        RECT 30.950 193.105 31.120 193.275 ;
        RECT 36.240 214.625 36.410 214.795 ;
        RECT 36.240 214.265 36.410 214.435 ;
        RECT 36.240 213.905 36.410 214.075 ;
        RECT 42.360 215.025 42.530 215.195 ;
        RECT 42.360 214.665 42.530 214.835 ;
        RECT 47.650 215.025 47.820 215.195 ;
        RECT 52.940 215.025 53.110 215.195 ;
        RECT 58.230 215.025 58.400 215.195 ;
        RECT 63.520 215.025 63.690 215.195 ;
        RECT 42.360 214.305 42.530 214.475 ;
        RECT 42.360 213.945 42.530 214.115 ;
        RECT 36.240 209.515 36.410 209.685 ;
        RECT 36.240 209.155 36.410 209.325 ;
        RECT 36.240 208.795 36.410 208.965 ;
        RECT 36.240 208.435 36.410 208.605 ;
        RECT 36.240 204.045 36.410 204.215 ;
        RECT 36.240 203.685 36.410 203.855 ;
        RECT 36.240 203.325 36.410 203.495 ;
        RECT 36.240 202.965 36.410 203.135 ;
        RECT 36.240 198.575 36.410 198.745 ;
        RECT 36.240 198.215 36.410 198.385 ;
        RECT 36.240 197.855 36.410 198.025 ;
        RECT 36.240 197.495 36.410 197.665 ;
        RECT 25.660 192.745 25.830 192.915 ;
        RECT 25.660 192.385 25.830 192.555 ;
        RECT 30.950 192.745 31.120 192.915 ;
        RECT 30.950 192.385 31.120 192.555 ;
        RECT 36.240 193.105 36.410 193.275 ;
        RECT 36.240 192.745 36.410 192.915 ;
        RECT 20.370 192.025 20.540 192.195 ;
        RECT 25.660 192.025 25.830 192.195 ;
        RECT 30.950 192.025 31.120 192.195 ;
        RECT 36.240 192.385 36.410 192.555 ;
        RECT 36.240 192.025 36.410 192.195 ;
        RECT 39.350 207.435 39.520 207.605 ;
        RECT 39.350 207.075 39.520 207.245 ;
        RECT 39.350 206.715 39.520 206.885 ;
        RECT 39.350 206.355 39.520 206.525 ;
        RECT 39.350 205.995 39.520 206.165 ;
        RECT 39.350 205.635 39.520 205.805 ;
        RECT 39.350 205.275 39.520 205.445 ;
        RECT 39.350 204.915 39.520 205.085 ;
        RECT 39.350 204.555 39.520 204.725 ;
        RECT 39.350 204.195 39.520 204.365 ;
        RECT 39.350 203.835 39.520 204.005 ;
        RECT 39.350 203.475 39.520 203.645 ;
        RECT 39.350 203.115 39.520 203.285 ;
        RECT 39.350 202.755 39.520 202.925 ;
        RECT 39.350 202.395 39.520 202.565 ;
        RECT 39.350 202.035 39.520 202.205 ;
        RECT 39.350 201.675 39.520 201.845 ;
        RECT 9.790 185.905 9.960 186.075 ;
        RECT 9.790 185.545 9.960 185.715 ;
        RECT 15.080 185.905 15.250 186.075 ;
        RECT 20.370 185.905 20.540 186.075 ;
        RECT 25.660 185.905 25.830 186.075 ;
        RECT 30.950 185.905 31.120 186.075 ;
        RECT 9.790 185.185 9.960 185.355 ;
        RECT 9.790 184.825 9.960 184.995 ;
        RECT 9.790 180.435 9.960 180.605 ;
        RECT 9.790 180.075 9.960 180.245 ;
        RECT 9.790 179.715 9.960 179.885 ;
        RECT 9.790 179.355 9.960 179.525 ;
        RECT 6.780 178.315 6.950 178.485 ;
        RECT 6.780 177.955 6.950 178.125 ;
        RECT 6.780 177.595 6.950 177.765 ;
        RECT 6.780 177.235 6.950 177.405 ;
        RECT 6.780 176.875 6.950 177.045 ;
        RECT 6.780 176.515 6.950 176.685 ;
        RECT 6.780 176.155 6.950 176.325 ;
        RECT 6.780 175.795 6.950 175.965 ;
        RECT 6.780 175.435 6.950 175.605 ;
        RECT 6.780 175.075 6.950 175.245 ;
        RECT 6.780 174.715 6.950 174.885 ;
        RECT 6.780 174.355 6.950 174.525 ;
        RECT 6.780 173.995 6.950 174.165 ;
        RECT 6.780 173.635 6.950 173.805 ;
        RECT 6.780 173.275 6.950 173.445 ;
        RECT 6.780 172.915 6.950 173.085 ;
        RECT 6.780 172.555 6.950 172.725 ;
        RECT 9.790 174.965 9.960 175.135 ;
        RECT 9.790 174.605 9.960 174.775 ;
        RECT 9.790 174.245 9.960 174.415 ;
        RECT 9.790 173.885 9.960 174.055 ;
        RECT 9.790 169.495 9.960 169.665 ;
        RECT 9.790 169.135 9.960 169.305 ;
        RECT 9.790 168.775 9.960 168.945 ;
        RECT 9.790 168.415 9.960 168.585 ;
        RECT 9.790 164.025 9.960 164.195 ;
        RECT 15.080 185.545 15.250 185.715 ;
        RECT 15.080 185.185 15.250 185.355 ;
        RECT 15.080 184.825 15.250 184.995 ;
        RECT 15.080 180.435 15.250 180.605 ;
        RECT 15.080 180.075 15.250 180.245 ;
        RECT 15.080 179.715 15.250 179.885 ;
        RECT 15.080 179.355 15.250 179.525 ;
        RECT 15.080 174.965 15.250 175.135 ;
        RECT 15.080 174.605 15.250 174.775 ;
        RECT 15.080 174.245 15.250 174.415 ;
        RECT 15.080 173.885 15.250 174.055 ;
        RECT 15.080 169.495 15.250 169.665 ;
        RECT 15.080 169.135 15.250 169.305 ;
        RECT 15.080 168.775 15.250 168.945 ;
        RECT 15.080 168.415 15.250 168.585 ;
        RECT 15.080 164.025 15.250 164.195 ;
        RECT 20.370 185.545 20.540 185.715 ;
        RECT 20.370 185.185 20.540 185.355 ;
        RECT 20.370 184.825 20.540 184.995 ;
        RECT 20.370 180.435 20.540 180.605 ;
        RECT 20.370 180.075 20.540 180.245 ;
        RECT 20.370 179.715 20.540 179.885 ;
        RECT 20.370 179.355 20.540 179.525 ;
        RECT 20.370 174.965 20.540 175.135 ;
        RECT 20.370 174.605 20.540 174.775 ;
        RECT 20.370 174.245 20.540 174.415 ;
        RECT 20.370 173.885 20.540 174.055 ;
        RECT 20.370 169.495 20.540 169.665 ;
        RECT 20.370 169.135 20.540 169.305 ;
        RECT 20.370 168.775 20.540 168.945 ;
        RECT 20.370 168.415 20.540 168.585 ;
        RECT 20.370 164.025 20.540 164.195 ;
        RECT 36.240 185.905 36.410 186.075 ;
        RECT 25.660 185.545 25.830 185.715 ;
        RECT 25.660 185.185 25.830 185.355 ;
        RECT 25.660 184.825 25.830 184.995 ;
        RECT 25.660 180.435 25.830 180.605 ;
        RECT 25.660 180.075 25.830 180.245 ;
        RECT 25.660 179.715 25.830 179.885 ;
        RECT 25.660 179.355 25.830 179.525 ;
        RECT 25.660 174.965 25.830 175.135 ;
        RECT 25.660 174.605 25.830 174.775 ;
        RECT 25.660 174.245 25.830 174.415 ;
        RECT 25.660 173.885 25.830 174.055 ;
        RECT 25.660 169.495 25.830 169.665 ;
        RECT 25.660 169.135 25.830 169.305 ;
        RECT 25.660 168.775 25.830 168.945 ;
        RECT 25.660 168.415 25.830 168.585 ;
        RECT 25.660 164.025 25.830 164.195 ;
        RECT 30.950 185.545 31.120 185.715 ;
        RECT 30.950 185.185 31.120 185.355 ;
        RECT 30.950 184.825 31.120 184.995 ;
        RECT 30.950 180.435 31.120 180.605 ;
        RECT 30.950 180.075 31.120 180.245 ;
        RECT 30.950 179.715 31.120 179.885 ;
        RECT 30.950 179.355 31.120 179.525 ;
        RECT 30.950 174.965 31.120 175.135 ;
        RECT 30.950 174.605 31.120 174.775 ;
        RECT 30.950 174.245 31.120 174.415 ;
        RECT 30.950 173.885 31.120 174.055 ;
        RECT 30.950 169.495 31.120 169.665 ;
        RECT 30.950 169.135 31.120 169.305 ;
        RECT 30.950 168.775 31.120 168.945 ;
        RECT 30.950 168.415 31.120 168.585 ;
        RECT 9.790 163.665 9.960 163.835 ;
        RECT 9.790 163.305 9.960 163.475 ;
        RECT 15.080 163.665 15.250 163.835 ;
        RECT 9.790 162.945 9.960 163.115 ;
        RECT 15.080 163.305 15.250 163.475 ;
        RECT 20.370 163.665 20.540 163.835 ;
        RECT 15.080 162.945 15.250 163.115 ;
        RECT 20.370 163.305 20.540 163.475 ;
        RECT 30.950 164.025 31.120 164.195 ;
        RECT 36.240 185.545 36.410 185.715 ;
        RECT 36.240 185.185 36.410 185.355 ;
        RECT 36.240 184.825 36.410 184.995 ;
        RECT 36.240 180.435 36.410 180.605 ;
        RECT 36.240 180.075 36.410 180.245 ;
        RECT 36.240 179.715 36.410 179.885 ;
        RECT 36.240 179.355 36.410 179.525 ;
        RECT 36.240 174.965 36.410 175.135 ;
        RECT 36.240 174.605 36.410 174.775 ;
        RECT 36.240 174.245 36.410 174.415 ;
        RECT 36.240 173.885 36.410 174.055 ;
        RECT 36.240 169.495 36.410 169.665 ;
        RECT 36.240 169.135 36.410 169.305 ;
        RECT 36.240 168.775 36.410 168.945 ;
        RECT 36.240 168.415 36.410 168.585 ;
        RECT 25.660 163.665 25.830 163.835 ;
        RECT 25.660 163.305 25.830 163.475 ;
        RECT 30.950 163.665 31.120 163.835 ;
        RECT 30.950 163.305 31.120 163.475 ;
        RECT 36.240 164.025 36.410 164.195 ;
        RECT 36.240 163.665 36.410 163.835 ;
        RECT 20.370 162.945 20.540 163.115 ;
        RECT 25.660 162.945 25.830 163.115 ;
        RECT 30.950 162.945 31.120 163.115 ;
        RECT 36.240 163.305 36.410 163.475 ;
        RECT 36.240 162.945 36.410 163.115 ;
        RECT 42.360 209.555 42.530 209.725 ;
        RECT 42.360 209.195 42.530 209.365 ;
        RECT 42.360 208.835 42.530 209.005 ;
        RECT 42.360 208.475 42.530 208.645 ;
        RECT 42.360 204.085 42.530 204.255 ;
        RECT 42.360 203.725 42.530 203.895 ;
        RECT 42.360 203.365 42.530 203.535 ;
        RECT 42.360 203.005 42.530 203.175 ;
        RECT 42.360 198.615 42.530 198.785 ;
        RECT 42.360 198.255 42.530 198.425 ;
        RECT 42.360 197.895 42.530 198.065 ;
        RECT 42.360 197.535 42.530 197.705 ;
        RECT 42.360 193.145 42.530 193.315 ;
        RECT 47.650 214.665 47.820 214.835 ;
        RECT 47.650 214.305 47.820 214.475 ;
        RECT 47.650 213.945 47.820 214.115 ;
        RECT 47.650 209.555 47.820 209.725 ;
        RECT 47.650 209.195 47.820 209.365 ;
        RECT 47.650 208.835 47.820 209.005 ;
        RECT 47.650 208.475 47.820 208.645 ;
        RECT 47.650 204.085 47.820 204.255 ;
        RECT 47.650 203.725 47.820 203.895 ;
        RECT 47.650 203.365 47.820 203.535 ;
        RECT 47.650 203.005 47.820 203.175 ;
        RECT 47.650 198.615 47.820 198.785 ;
        RECT 47.650 198.255 47.820 198.425 ;
        RECT 47.650 197.895 47.820 198.065 ;
        RECT 47.650 197.535 47.820 197.705 ;
        RECT 47.650 193.145 47.820 193.315 ;
        RECT 52.940 214.665 53.110 214.835 ;
        RECT 52.940 214.305 53.110 214.475 ;
        RECT 52.940 213.945 53.110 214.115 ;
        RECT 52.940 209.555 53.110 209.725 ;
        RECT 52.940 209.195 53.110 209.365 ;
        RECT 52.940 208.835 53.110 209.005 ;
        RECT 52.940 208.475 53.110 208.645 ;
        RECT 52.940 204.085 53.110 204.255 ;
        RECT 52.940 203.725 53.110 203.895 ;
        RECT 52.940 203.365 53.110 203.535 ;
        RECT 52.940 203.005 53.110 203.175 ;
        RECT 52.940 198.615 53.110 198.785 ;
        RECT 52.940 198.255 53.110 198.425 ;
        RECT 52.940 197.895 53.110 198.065 ;
        RECT 52.940 197.535 53.110 197.705 ;
        RECT 52.940 193.145 53.110 193.315 ;
        RECT 68.810 215.025 68.980 215.195 ;
        RECT 74.890 215.065 75.060 215.235 ;
        RECT 58.230 214.665 58.400 214.835 ;
        RECT 58.230 214.305 58.400 214.475 ;
        RECT 58.230 213.945 58.400 214.115 ;
        RECT 58.230 209.555 58.400 209.725 ;
        RECT 58.230 209.195 58.400 209.365 ;
        RECT 58.230 208.835 58.400 209.005 ;
        RECT 58.230 208.475 58.400 208.645 ;
        RECT 58.230 204.085 58.400 204.255 ;
        RECT 58.230 203.725 58.400 203.895 ;
        RECT 58.230 203.365 58.400 203.535 ;
        RECT 58.230 203.005 58.400 203.175 ;
        RECT 58.230 198.615 58.400 198.785 ;
        RECT 58.230 198.255 58.400 198.425 ;
        RECT 58.230 197.895 58.400 198.065 ;
        RECT 58.230 197.535 58.400 197.705 ;
        RECT 58.230 193.145 58.400 193.315 ;
        RECT 63.520 214.665 63.690 214.835 ;
        RECT 63.520 214.305 63.690 214.475 ;
        RECT 63.520 213.945 63.690 214.115 ;
        RECT 63.520 209.555 63.690 209.725 ;
        RECT 63.520 209.195 63.690 209.365 ;
        RECT 63.520 208.835 63.690 209.005 ;
        RECT 63.520 208.475 63.690 208.645 ;
        RECT 63.520 204.085 63.690 204.255 ;
        RECT 63.520 203.725 63.690 203.895 ;
        RECT 63.520 203.365 63.690 203.535 ;
        RECT 63.520 203.005 63.690 203.175 ;
        RECT 63.520 198.615 63.690 198.785 ;
        RECT 63.520 198.255 63.690 198.425 ;
        RECT 63.520 197.895 63.690 198.065 ;
        RECT 63.520 197.535 63.690 197.705 ;
        RECT 42.360 192.785 42.530 192.955 ;
        RECT 42.360 192.425 42.530 192.595 ;
        RECT 47.650 192.785 47.820 192.955 ;
        RECT 42.360 192.065 42.530 192.235 ;
        RECT 47.650 192.425 47.820 192.595 ;
        RECT 52.940 192.785 53.110 192.955 ;
        RECT 47.650 192.065 47.820 192.235 ;
        RECT 52.940 192.425 53.110 192.595 ;
        RECT 63.520 193.145 63.690 193.315 ;
        RECT 68.810 214.665 68.980 214.835 ;
        RECT 68.810 214.305 68.980 214.475 ;
        RECT 68.810 213.945 68.980 214.115 ;
        RECT 68.810 209.555 68.980 209.725 ;
        RECT 68.810 209.195 68.980 209.365 ;
        RECT 68.810 208.835 68.980 209.005 ;
        RECT 68.810 208.475 68.980 208.645 ;
        RECT 74.890 214.705 75.060 214.875 ;
        RECT 80.180 215.065 80.350 215.235 ;
        RECT 85.470 215.065 85.640 215.235 ;
        RECT 90.760 215.065 90.930 215.235 ;
        RECT 96.050 215.065 96.220 215.235 ;
        RECT 74.890 214.345 75.060 214.515 ;
        RECT 74.890 213.985 75.060 214.155 ;
        RECT 74.890 209.595 75.060 209.765 ;
        RECT 74.890 209.235 75.060 209.405 ;
        RECT 74.890 208.875 75.060 209.045 ;
        RECT 74.890 208.515 75.060 208.685 ;
        RECT 68.810 204.085 68.980 204.255 ;
        RECT 68.810 203.725 68.980 203.895 ;
        RECT 68.810 203.365 68.980 203.535 ;
        RECT 68.810 203.005 68.980 203.175 ;
        RECT 68.810 198.615 68.980 198.785 ;
        RECT 68.810 198.255 68.980 198.425 ;
        RECT 68.810 197.895 68.980 198.065 ;
        RECT 68.810 197.535 68.980 197.705 ;
        RECT 58.230 192.785 58.400 192.955 ;
        RECT 58.230 192.425 58.400 192.595 ;
        RECT 68.810 193.145 68.980 193.315 ;
        RECT 63.520 192.785 63.690 192.955 ;
        RECT 63.520 192.425 63.690 192.595 ;
        RECT 68.810 192.785 68.980 192.955 ;
        RECT 52.940 192.065 53.110 192.235 ;
        RECT 58.230 192.065 58.400 192.235 ;
        RECT 63.520 192.065 63.690 192.235 ;
        RECT 68.810 192.425 68.980 192.595 ;
        RECT 68.810 192.065 68.980 192.235 ;
        RECT 71.880 207.475 72.050 207.645 ;
        RECT 71.880 207.115 72.050 207.285 ;
        RECT 71.880 206.755 72.050 206.925 ;
        RECT 71.880 206.395 72.050 206.565 ;
        RECT 71.880 206.035 72.050 206.205 ;
        RECT 71.880 205.675 72.050 205.845 ;
        RECT 71.880 205.315 72.050 205.485 ;
        RECT 71.880 204.955 72.050 205.125 ;
        RECT 71.880 204.595 72.050 204.765 ;
        RECT 71.880 204.235 72.050 204.405 ;
        RECT 71.880 203.875 72.050 204.045 ;
        RECT 71.880 203.515 72.050 203.685 ;
        RECT 71.880 203.155 72.050 203.325 ;
        RECT 71.880 202.795 72.050 202.965 ;
        RECT 71.880 202.435 72.050 202.605 ;
        RECT 71.880 202.075 72.050 202.245 ;
        RECT 71.880 201.715 72.050 201.885 ;
        RECT 39.350 178.355 39.520 178.525 ;
        RECT 39.350 177.995 39.520 178.165 ;
        RECT 39.350 177.635 39.520 177.805 ;
        RECT 39.350 177.275 39.520 177.445 ;
        RECT 39.350 176.915 39.520 177.085 ;
        RECT 39.350 176.555 39.520 176.725 ;
        RECT 39.350 176.195 39.520 176.365 ;
        RECT 39.350 175.835 39.520 176.005 ;
        RECT 39.350 175.475 39.520 175.645 ;
        RECT 39.350 175.115 39.520 175.285 ;
        RECT 39.350 174.755 39.520 174.925 ;
        RECT 39.350 174.395 39.520 174.565 ;
        RECT 39.350 174.035 39.520 174.205 ;
        RECT 39.350 173.675 39.520 173.845 ;
        RECT 39.350 173.315 39.520 173.485 ;
        RECT 39.350 172.955 39.520 173.125 ;
        RECT 39.350 172.595 39.520 172.765 ;
        RECT 9.790 156.735 9.960 156.905 ;
        RECT 9.790 156.375 9.960 156.545 ;
        RECT 15.080 156.735 15.250 156.905 ;
        RECT 20.370 156.735 20.540 156.905 ;
        RECT 25.660 156.735 25.830 156.905 ;
        RECT 30.950 156.735 31.120 156.905 ;
        RECT 9.790 156.015 9.960 156.185 ;
        RECT 9.790 155.655 9.960 155.825 ;
        RECT 9.790 151.265 9.960 151.435 ;
        RECT 9.790 150.905 9.960 151.075 ;
        RECT 9.790 150.545 9.960 150.715 ;
        RECT 9.790 150.185 9.960 150.355 ;
        RECT 6.780 149.145 6.950 149.315 ;
        RECT 6.780 148.785 6.950 148.955 ;
        RECT 6.780 148.425 6.950 148.595 ;
        RECT 6.780 148.065 6.950 148.235 ;
        RECT 6.780 147.705 6.950 147.875 ;
        RECT 6.780 147.345 6.950 147.515 ;
        RECT 6.780 146.985 6.950 147.155 ;
        RECT 6.780 146.625 6.950 146.795 ;
        RECT 6.780 146.265 6.950 146.435 ;
        RECT 6.780 145.905 6.950 146.075 ;
        RECT 6.780 145.545 6.950 145.715 ;
        RECT 6.780 145.185 6.950 145.355 ;
        RECT 6.780 144.825 6.950 144.995 ;
        RECT 6.780 144.465 6.950 144.635 ;
        RECT 6.780 144.105 6.950 144.275 ;
        RECT 6.780 143.745 6.950 143.915 ;
        RECT 6.780 143.385 6.950 143.555 ;
        RECT 9.790 145.795 9.960 145.965 ;
        RECT 9.790 145.435 9.960 145.605 ;
        RECT 9.790 145.075 9.960 145.245 ;
        RECT 9.790 144.715 9.960 144.885 ;
        RECT 9.790 140.325 9.960 140.495 ;
        RECT 9.790 139.965 9.960 140.135 ;
        RECT 9.790 139.605 9.960 139.775 ;
        RECT 9.790 139.245 9.960 139.415 ;
        RECT -97.560 134.345 -97.390 134.515 ;
        RECT -97.560 133.985 -97.390 134.155 ;
        RECT -97.560 133.625 -97.390 133.795 ;
        RECT -97.560 133.265 -97.390 133.435 ;
        RECT -94.980 134.345 -94.810 134.515 ;
        RECT -94.980 133.985 -94.810 134.155 ;
        RECT -94.980 133.625 -94.810 133.795 ;
        RECT -94.980 133.265 -94.810 133.435 ;
        RECT -92.400 134.345 -92.230 134.515 ;
        RECT -92.400 133.985 -92.230 134.155 ;
        RECT -92.400 133.625 -92.230 133.795 ;
        RECT -92.400 133.265 -92.230 133.435 ;
        RECT -89.820 134.345 -89.650 134.515 ;
        RECT -89.820 133.985 -89.650 134.155 ;
        RECT -89.820 133.625 -89.650 133.795 ;
        RECT -89.820 133.265 -89.650 133.435 ;
        RECT -87.240 134.345 -87.070 134.515 ;
        RECT -87.240 133.985 -87.070 134.155 ;
        RECT -87.240 133.625 -87.070 133.795 ;
        RECT -87.240 133.265 -87.070 133.435 ;
        RECT -84.660 134.345 -84.490 134.515 ;
        RECT -84.660 133.985 -84.490 134.155 ;
        RECT -84.660 133.625 -84.490 133.795 ;
        RECT -84.660 133.265 -84.490 133.435 ;
        RECT -82.080 134.345 -81.910 134.515 ;
        RECT -82.080 133.985 -81.910 134.155 ;
        RECT -82.080 133.625 -81.910 133.795 ;
        RECT -82.080 133.265 -81.910 133.435 ;
        RECT -79.500 134.345 -79.330 134.515 ;
        RECT -79.500 133.985 -79.330 134.155 ;
        RECT -79.500 133.625 -79.330 133.795 ;
        RECT -79.500 133.265 -79.330 133.435 ;
        RECT -76.920 134.345 -76.750 134.515 ;
        RECT -76.920 133.985 -76.750 134.155 ;
        RECT -76.920 133.625 -76.750 133.795 ;
        RECT -76.920 133.265 -76.750 133.435 ;
        RECT -74.340 134.345 -74.170 134.515 ;
        RECT -74.340 133.985 -74.170 134.155 ;
        RECT -74.340 133.625 -74.170 133.795 ;
        RECT -74.340 133.265 -74.170 133.435 ;
        RECT -71.760 134.345 -71.590 134.515 ;
        RECT -71.760 133.985 -71.590 134.155 ;
        RECT -71.760 133.625 -71.590 133.795 ;
        RECT -71.760 133.265 -71.590 133.435 ;
        RECT 9.790 134.855 9.960 135.025 ;
        RECT 15.080 156.375 15.250 156.545 ;
        RECT 15.080 156.015 15.250 156.185 ;
        RECT 15.080 155.655 15.250 155.825 ;
        RECT 15.080 151.265 15.250 151.435 ;
        RECT 15.080 150.905 15.250 151.075 ;
        RECT 15.080 150.545 15.250 150.715 ;
        RECT 15.080 150.185 15.250 150.355 ;
        RECT 15.080 145.795 15.250 145.965 ;
        RECT 15.080 145.435 15.250 145.605 ;
        RECT 15.080 145.075 15.250 145.245 ;
        RECT 15.080 144.715 15.250 144.885 ;
        RECT 15.080 140.325 15.250 140.495 ;
        RECT 15.080 139.965 15.250 140.135 ;
        RECT 15.080 139.605 15.250 139.775 ;
        RECT 15.080 139.245 15.250 139.415 ;
        RECT 15.080 134.855 15.250 135.025 ;
        RECT 20.370 156.375 20.540 156.545 ;
        RECT 20.370 156.015 20.540 156.185 ;
        RECT 20.370 155.655 20.540 155.825 ;
        RECT 20.370 151.265 20.540 151.435 ;
        RECT 20.370 150.905 20.540 151.075 ;
        RECT 20.370 150.545 20.540 150.715 ;
        RECT 20.370 150.185 20.540 150.355 ;
        RECT 20.370 145.795 20.540 145.965 ;
        RECT 20.370 145.435 20.540 145.605 ;
        RECT 20.370 145.075 20.540 145.245 ;
        RECT 20.370 144.715 20.540 144.885 ;
        RECT 20.370 140.325 20.540 140.495 ;
        RECT 20.370 139.965 20.540 140.135 ;
        RECT 20.370 139.605 20.540 139.775 ;
        RECT 20.370 139.245 20.540 139.415 ;
        RECT 20.370 134.855 20.540 135.025 ;
        RECT 36.240 156.735 36.410 156.905 ;
        RECT 25.660 156.375 25.830 156.545 ;
        RECT 25.660 156.015 25.830 156.185 ;
        RECT 25.660 155.655 25.830 155.825 ;
        RECT 25.660 151.265 25.830 151.435 ;
        RECT 25.660 150.905 25.830 151.075 ;
        RECT 25.660 150.545 25.830 150.715 ;
        RECT 25.660 150.185 25.830 150.355 ;
        RECT 25.660 145.795 25.830 145.965 ;
        RECT 25.660 145.435 25.830 145.605 ;
        RECT 25.660 145.075 25.830 145.245 ;
        RECT 25.660 144.715 25.830 144.885 ;
        RECT 25.660 140.325 25.830 140.495 ;
        RECT 25.660 139.965 25.830 140.135 ;
        RECT 25.660 139.605 25.830 139.775 ;
        RECT 25.660 139.245 25.830 139.415 ;
        RECT 25.660 134.855 25.830 135.025 ;
        RECT 30.950 156.375 31.120 156.545 ;
        RECT 30.950 156.015 31.120 156.185 ;
        RECT 30.950 155.655 31.120 155.825 ;
        RECT 30.950 151.265 31.120 151.435 ;
        RECT 30.950 150.905 31.120 151.075 ;
        RECT 30.950 150.545 31.120 150.715 ;
        RECT 30.950 150.185 31.120 150.355 ;
        RECT 30.950 145.795 31.120 145.965 ;
        RECT 30.950 145.435 31.120 145.605 ;
        RECT 30.950 145.075 31.120 145.245 ;
        RECT 30.950 144.715 31.120 144.885 ;
        RECT 30.950 140.325 31.120 140.495 ;
        RECT 30.950 139.965 31.120 140.135 ;
        RECT 30.950 139.605 31.120 139.775 ;
        RECT 30.950 139.245 31.120 139.415 ;
        RECT 9.790 134.495 9.960 134.665 ;
        RECT 9.790 134.135 9.960 134.305 ;
        RECT 15.080 134.495 15.250 134.665 ;
        RECT 9.790 133.775 9.960 133.945 ;
        RECT -96.915 131.030 -96.745 131.200 ;
        RECT -95.625 131.030 -95.455 131.200 ;
        RECT -94.335 131.030 -94.165 131.200 ;
        RECT -93.045 131.030 -92.875 131.200 ;
        RECT -91.755 131.030 -91.585 131.200 ;
        RECT -90.465 131.030 -90.295 131.200 ;
        RECT -89.175 131.030 -89.005 131.200 ;
        RECT -87.885 131.030 -87.715 131.200 ;
        RECT -86.595 131.030 -86.425 131.200 ;
        RECT -85.305 131.030 -85.135 131.200 ;
        RECT -84.015 131.030 -83.845 131.200 ;
        RECT -82.725 131.030 -82.555 131.200 ;
        RECT -81.435 131.030 -81.265 131.200 ;
        RECT -80.145 131.030 -79.975 131.200 ;
        RECT -78.855 131.030 -78.685 131.200 ;
        RECT -77.565 131.030 -77.395 131.200 ;
        RECT -76.275 131.030 -76.105 131.200 ;
        RECT -74.985 131.030 -74.815 131.200 ;
        RECT -73.695 131.030 -73.525 131.200 ;
        RECT -72.405 131.030 -72.235 131.200 ;
        RECT -91.440 128.035 -77.950 130.365 ;
        RECT 15.080 134.135 15.250 134.305 ;
        RECT 20.370 134.495 20.540 134.665 ;
        RECT 15.080 133.775 15.250 133.945 ;
        RECT 20.370 134.135 20.540 134.305 ;
        RECT 30.950 134.855 31.120 135.025 ;
        RECT 36.240 156.375 36.410 156.545 ;
        RECT 36.240 156.015 36.410 156.185 ;
        RECT 36.240 155.655 36.410 155.825 ;
        RECT 36.240 151.265 36.410 151.435 ;
        RECT 36.240 150.905 36.410 151.075 ;
        RECT 36.240 150.545 36.410 150.715 ;
        RECT 36.240 150.185 36.410 150.355 ;
        RECT 36.240 145.795 36.410 145.965 ;
        RECT 36.240 145.435 36.410 145.605 ;
        RECT 36.240 145.075 36.410 145.245 ;
        RECT 36.240 144.715 36.410 144.885 ;
        RECT 36.240 140.325 36.410 140.495 ;
        RECT 36.240 139.965 36.410 140.135 ;
        RECT 36.240 139.605 36.410 139.775 ;
        RECT 36.240 139.245 36.410 139.415 ;
        RECT 25.660 134.495 25.830 134.665 ;
        RECT 25.660 134.135 25.830 134.305 ;
        RECT 30.950 134.495 31.120 134.665 ;
        RECT 30.950 134.135 31.120 134.305 ;
        RECT 36.240 134.855 36.410 135.025 ;
        RECT 36.240 134.495 36.410 134.665 ;
        RECT 20.370 133.775 20.540 133.945 ;
        RECT 25.660 133.775 25.830 133.945 ;
        RECT 30.950 133.775 31.120 133.945 ;
        RECT 36.240 134.135 36.410 134.305 ;
        RECT 36.240 133.775 36.410 133.945 ;
        RECT 42.360 185.945 42.530 186.115 ;
        RECT 42.360 185.585 42.530 185.755 ;
        RECT 47.650 185.945 47.820 186.115 ;
        RECT 52.940 185.945 53.110 186.115 ;
        RECT 58.230 185.945 58.400 186.115 ;
        RECT 63.520 185.945 63.690 186.115 ;
        RECT 42.360 185.225 42.530 185.395 ;
        RECT 42.360 184.865 42.530 185.035 ;
        RECT 42.360 180.475 42.530 180.645 ;
        RECT 42.360 180.115 42.530 180.285 ;
        RECT 42.360 179.755 42.530 179.925 ;
        RECT 42.360 179.395 42.530 179.565 ;
        RECT 42.360 175.005 42.530 175.175 ;
        RECT 42.360 174.645 42.530 174.815 ;
        RECT 42.360 174.285 42.530 174.455 ;
        RECT 42.360 173.925 42.530 174.095 ;
        RECT 42.360 169.535 42.530 169.705 ;
        RECT 42.360 169.175 42.530 169.345 ;
        RECT 42.360 168.815 42.530 168.985 ;
        RECT 42.360 168.455 42.530 168.625 ;
        RECT 42.360 164.065 42.530 164.235 ;
        RECT 47.650 185.585 47.820 185.755 ;
        RECT 47.650 185.225 47.820 185.395 ;
        RECT 47.650 184.865 47.820 185.035 ;
        RECT 47.650 180.475 47.820 180.645 ;
        RECT 47.650 180.115 47.820 180.285 ;
        RECT 47.650 179.755 47.820 179.925 ;
        RECT 47.650 179.395 47.820 179.565 ;
        RECT 47.650 175.005 47.820 175.175 ;
        RECT 47.650 174.645 47.820 174.815 ;
        RECT 47.650 174.285 47.820 174.455 ;
        RECT 47.650 173.925 47.820 174.095 ;
        RECT 47.650 169.535 47.820 169.705 ;
        RECT 47.650 169.175 47.820 169.345 ;
        RECT 47.650 168.815 47.820 168.985 ;
        RECT 47.650 168.455 47.820 168.625 ;
        RECT 47.650 164.065 47.820 164.235 ;
        RECT 52.940 185.585 53.110 185.755 ;
        RECT 52.940 185.225 53.110 185.395 ;
        RECT 52.940 184.865 53.110 185.035 ;
        RECT 52.940 180.475 53.110 180.645 ;
        RECT 52.940 180.115 53.110 180.285 ;
        RECT 52.940 179.755 53.110 179.925 ;
        RECT 52.940 179.395 53.110 179.565 ;
        RECT 52.940 175.005 53.110 175.175 ;
        RECT 52.940 174.645 53.110 174.815 ;
        RECT 52.940 174.285 53.110 174.455 ;
        RECT 52.940 173.925 53.110 174.095 ;
        RECT 52.940 169.535 53.110 169.705 ;
        RECT 52.940 169.175 53.110 169.345 ;
        RECT 52.940 168.815 53.110 168.985 ;
        RECT 52.940 168.455 53.110 168.625 ;
        RECT 52.940 164.065 53.110 164.235 ;
        RECT 68.810 185.945 68.980 186.115 ;
        RECT 58.230 185.585 58.400 185.755 ;
        RECT 58.230 185.225 58.400 185.395 ;
        RECT 58.230 184.865 58.400 185.035 ;
        RECT 58.230 180.475 58.400 180.645 ;
        RECT 58.230 180.115 58.400 180.285 ;
        RECT 58.230 179.755 58.400 179.925 ;
        RECT 58.230 179.395 58.400 179.565 ;
        RECT 58.230 175.005 58.400 175.175 ;
        RECT 58.230 174.645 58.400 174.815 ;
        RECT 58.230 174.285 58.400 174.455 ;
        RECT 58.230 173.925 58.400 174.095 ;
        RECT 58.230 169.535 58.400 169.705 ;
        RECT 58.230 169.175 58.400 169.345 ;
        RECT 58.230 168.815 58.400 168.985 ;
        RECT 58.230 168.455 58.400 168.625 ;
        RECT 58.230 164.065 58.400 164.235 ;
        RECT 63.520 185.585 63.690 185.755 ;
        RECT 63.520 185.225 63.690 185.395 ;
        RECT 63.520 184.865 63.690 185.035 ;
        RECT 63.520 180.475 63.690 180.645 ;
        RECT 63.520 180.115 63.690 180.285 ;
        RECT 63.520 179.755 63.690 179.925 ;
        RECT 63.520 179.395 63.690 179.565 ;
        RECT 63.520 175.005 63.690 175.175 ;
        RECT 63.520 174.645 63.690 174.815 ;
        RECT 63.520 174.285 63.690 174.455 ;
        RECT 63.520 173.925 63.690 174.095 ;
        RECT 63.520 169.535 63.690 169.705 ;
        RECT 63.520 169.175 63.690 169.345 ;
        RECT 63.520 168.815 63.690 168.985 ;
        RECT 63.520 168.455 63.690 168.625 ;
        RECT 42.360 163.705 42.530 163.875 ;
        RECT 42.360 163.345 42.530 163.515 ;
        RECT 47.650 163.705 47.820 163.875 ;
        RECT 42.360 162.985 42.530 163.155 ;
        RECT 47.650 163.345 47.820 163.515 ;
        RECT 52.940 163.705 53.110 163.875 ;
        RECT 47.650 162.985 47.820 163.155 ;
        RECT 52.940 163.345 53.110 163.515 ;
        RECT 63.520 164.065 63.690 164.235 ;
        RECT 68.810 185.585 68.980 185.755 ;
        RECT 68.810 185.225 68.980 185.395 ;
        RECT 68.810 184.865 68.980 185.035 ;
        RECT 68.810 180.475 68.980 180.645 ;
        RECT 68.810 180.115 68.980 180.285 ;
        RECT 68.810 179.755 68.980 179.925 ;
        RECT 68.810 179.395 68.980 179.565 ;
        RECT 68.810 175.005 68.980 175.175 ;
        RECT 68.810 174.645 68.980 174.815 ;
        RECT 68.810 174.285 68.980 174.455 ;
        RECT 68.810 173.925 68.980 174.095 ;
        RECT 68.810 169.535 68.980 169.705 ;
        RECT 68.810 169.175 68.980 169.345 ;
        RECT 68.810 168.815 68.980 168.985 ;
        RECT 68.810 168.455 68.980 168.625 ;
        RECT 58.230 163.705 58.400 163.875 ;
        RECT 58.230 163.345 58.400 163.515 ;
        RECT 68.810 164.065 68.980 164.235 ;
        RECT 63.520 163.705 63.690 163.875 ;
        RECT 63.520 163.345 63.690 163.515 ;
        RECT 68.810 163.705 68.980 163.875 ;
        RECT 52.940 162.985 53.110 163.155 ;
        RECT 58.230 162.985 58.400 163.155 ;
        RECT 63.520 162.985 63.690 163.155 ;
        RECT 68.810 163.345 68.980 163.515 ;
        RECT 68.810 162.985 68.980 163.155 ;
        RECT 74.890 204.125 75.060 204.295 ;
        RECT 74.890 203.765 75.060 203.935 ;
        RECT 74.890 203.405 75.060 203.575 ;
        RECT 74.890 203.045 75.060 203.215 ;
        RECT 74.890 198.655 75.060 198.825 ;
        RECT 74.890 198.295 75.060 198.465 ;
        RECT 74.890 197.935 75.060 198.105 ;
        RECT 74.890 197.575 75.060 197.745 ;
        RECT 74.890 193.185 75.060 193.355 ;
        RECT 80.180 214.705 80.350 214.875 ;
        RECT 80.180 214.345 80.350 214.515 ;
        RECT 80.180 213.985 80.350 214.155 ;
        RECT 80.180 209.595 80.350 209.765 ;
        RECT 80.180 209.235 80.350 209.405 ;
        RECT 80.180 208.875 80.350 209.045 ;
        RECT 80.180 208.515 80.350 208.685 ;
        RECT 80.180 204.125 80.350 204.295 ;
        RECT 80.180 203.765 80.350 203.935 ;
        RECT 80.180 203.405 80.350 203.575 ;
        RECT 80.180 203.045 80.350 203.215 ;
        RECT 80.180 198.655 80.350 198.825 ;
        RECT 80.180 198.295 80.350 198.465 ;
        RECT 80.180 197.935 80.350 198.105 ;
        RECT 80.180 197.575 80.350 197.745 ;
        RECT 80.180 193.185 80.350 193.355 ;
        RECT 85.470 214.705 85.640 214.875 ;
        RECT 85.470 214.345 85.640 214.515 ;
        RECT 85.470 213.985 85.640 214.155 ;
        RECT 85.470 209.595 85.640 209.765 ;
        RECT 85.470 209.235 85.640 209.405 ;
        RECT 85.470 208.875 85.640 209.045 ;
        RECT 85.470 208.515 85.640 208.685 ;
        RECT 85.470 204.125 85.640 204.295 ;
        RECT 85.470 203.765 85.640 203.935 ;
        RECT 85.470 203.405 85.640 203.575 ;
        RECT 85.470 203.045 85.640 203.215 ;
        RECT 85.470 198.655 85.640 198.825 ;
        RECT 85.470 198.295 85.640 198.465 ;
        RECT 85.470 197.935 85.640 198.105 ;
        RECT 85.470 197.575 85.640 197.745 ;
        RECT 85.470 193.185 85.640 193.355 ;
        RECT 101.340 215.065 101.510 215.235 ;
        RECT 204.950 215.095 205.120 215.265 ;
        RECT 90.760 214.705 90.930 214.875 ;
        RECT 90.760 214.345 90.930 214.515 ;
        RECT 90.760 213.985 90.930 214.155 ;
        RECT 90.760 209.595 90.930 209.765 ;
        RECT 90.760 209.235 90.930 209.405 ;
        RECT 90.760 208.875 90.930 209.045 ;
        RECT 90.760 208.515 90.930 208.685 ;
        RECT 90.760 204.125 90.930 204.295 ;
        RECT 90.760 203.765 90.930 203.935 ;
        RECT 90.760 203.405 90.930 203.575 ;
        RECT 90.760 203.045 90.930 203.215 ;
        RECT 90.760 198.655 90.930 198.825 ;
        RECT 90.760 198.295 90.930 198.465 ;
        RECT 90.760 197.935 90.930 198.105 ;
        RECT 90.760 197.575 90.930 197.745 ;
        RECT 90.760 193.185 90.930 193.355 ;
        RECT 96.050 214.705 96.220 214.875 ;
        RECT 96.050 214.345 96.220 214.515 ;
        RECT 96.050 213.985 96.220 214.155 ;
        RECT 96.050 209.595 96.220 209.765 ;
        RECT 96.050 209.235 96.220 209.405 ;
        RECT 96.050 208.875 96.220 209.045 ;
        RECT 96.050 208.515 96.220 208.685 ;
        RECT 96.050 204.125 96.220 204.295 ;
        RECT 96.050 203.765 96.220 203.935 ;
        RECT 96.050 203.405 96.220 203.575 ;
        RECT 96.050 203.045 96.220 203.215 ;
        RECT 96.050 198.655 96.220 198.825 ;
        RECT 96.050 198.295 96.220 198.465 ;
        RECT 96.050 197.935 96.220 198.105 ;
        RECT 96.050 197.575 96.220 197.745 ;
        RECT 74.890 192.825 75.060 192.995 ;
        RECT 74.890 192.465 75.060 192.635 ;
        RECT 80.180 192.825 80.350 192.995 ;
        RECT 74.890 192.105 75.060 192.275 ;
        RECT 80.180 192.465 80.350 192.635 ;
        RECT 85.470 192.825 85.640 192.995 ;
        RECT 80.180 192.105 80.350 192.275 ;
        RECT 85.470 192.465 85.640 192.635 ;
        RECT 96.050 193.185 96.220 193.355 ;
        RECT 101.340 214.705 101.510 214.875 ;
        RECT 101.340 214.345 101.510 214.515 ;
        RECT 101.340 213.985 101.510 214.155 ;
        RECT 204.950 214.735 205.120 214.905 ;
        RECT 210.240 215.095 210.410 215.265 ;
        RECT 215.530 215.095 215.700 215.265 ;
        RECT 220.820 215.095 220.990 215.265 ;
        RECT 226.110 215.095 226.280 215.265 ;
        RECT 204.950 214.375 205.120 214.545 ;
        RECT 101.340 209.595 101.510 209.765 ;
        RECT 101.340 209.235 101.510 209.405 ;
        RECT 101.340 208.875 101.510 209.045 ;
        RECT 101.340 208.515 101.510 208.685 ;
        RECT 101.340 204.125 101.510 204.295 ;
        RECT 101.340 203.765 101.510 203.935 ;
        RECT 101.340 203.405 101.510 203.575 ;
        RECT 101.340 203.045 101.510 203.215 ;
        RECT 101.340 198.655 101.510 198.825 ;
        RECT 101.340 198.295 101.510 198.465 ;
        RECT 101.340 197.935 101.510 198.105 ;
        RECT 101.340 197.575 101.510 197.745 ;
        RECT 90.760 192.825 90.930 192.995 ;
        RECT 90.760 192.465 90.930 192.635 ;
        RECT 96.050 192.825 96.220 192.995 ;
        RECT 96.050 192.465 96.220 192.635 ;
        RECT 85.470 192.105 85.640 192.275 ;
        RECT 90.760 192.105 90.930 192.275 ;
        RECT 96.050 192.105 96.220 192.275 ;
        RECT 101.340 193.185 101.510 193.355 ;
        RECT 101.340 192.825 101.510 192.995 ;
        RECT 101.340 192.465 101.510 192.635 ;
        RECT 101.340 192.105 101.510 192.275 ;
        RECT 104.330 207.395 104.500 207.565 ;
        RECT 104.330 207.035 104.500 207.205 ;
        RECT 104.330 206.675 104.500 206.845 ;
        RECT 104.330 206.315 104.500 206.485 ;
        RECT 104.330 205.955 104.500 206.125 ;
        RECT 104.330 205.595 104.500 205.765 ;
        RECT 104.330 205.235 104.500 205.405 ;
        RECT 104.330 204.875 104.500 205.045 ;
        RECT 104.330 204.515 104.500 204.685 ;
        RECT 104.330 204.155 104.500 204.325 ;
        RECT 104.330 203.795 104.500 203.965 ;
        RECT 104.330 203.435 104.500 203.605 ;
        RECT 104.330 203.075 104.500 203.245 ;
        RECT 104.330 202.715 104.500 202.885 ;
        RECT 104.330 202.355 104.500 202.525 ;
        RECT 104.330 201.995 104.500 202.165 ;
        RECT 104.330 201.635 104.500 201.805 ;
        RECT 71.880 178.395 72.050 178.565 ;
        RECT 71.880 178.035 72.050 178.205 ;
        RECT 71.880 177.675 72.050 177.845 ;
        RECT 71.880 177.315 72.050 177.485 ;
        RECT 71.880 176.955 72.050 177.125 ;
        RECT 71.880 176.595 72.050 176.765 ;
        RECT 71.880 176.235 72.050 176.405 ;
        RECT 71.880 175.875 72.050 176.045 ;
        RECT 71.880 175.515 72.050 175.685 ;
        RECT 71.880 175.155 72.050 175.325 ;
        RECT 71.880 174.795 72.050 174.965 ;
        RECT 71.880 174.435 72.050 174.605 ;
        RECT 71.880 174.075 72.050 174.245 ;
        RECT 71.880 173.715 72.050 173.885 ;
        RECT 71.880 173.355 72.050 173.525 ;
        RECT 71.880 172.995 72.050 173.165 ;
        RECT 71.880 172.635 72.050 172.805 ;
        RECT 39.350 149.185 39.520 149.355 ;
        RECT 39.350 148.825 39.520 148.995 ;
        RECT 39.350 148.465 39.520 148.635 ;
        RECT 39.350 148.105 39.520 148.275 ;
        RECT 39.350 147.745 39.520 147.915 ;
        RECT 39.350 147.385 39.520 147.555 ;
        RECT 39.350 147.025 39.520 147.195 ;
        RECT 39.350 146.665 39.520 146.835 ;
        RECT 39.350 146.305 39.520 146.475 ;
        RECT 39.350 145.945 39.520 146.115 ;
        RECT 39.350 145.585 39.520 145.755 ;
        RECT 39.350 145.225 39.520 145.395 ;
        RECT 39.350 144.865 39.520 145.035 ;
        RECT 39.350 144.505 39.520 144.675 ;
        RECT 39.350 144.145 39.520 144.315 ;
        RECT 39.350 143.785 39.520 143.955 ;
        RECT 39.350 143.425 39.520 143.595 ;
        RECT 9.790 127.555 9.960 127.725 ;
        RECT 9.790 127.195 9.960 127.365 ;
        RECT 15.080 127.555 15.250 127.725 ;
        RECT 20.370 127.555 20.540 127.725 ;
        RECT 25.660 127.555 25.830 127.725 ;
        RECT 30.950 127.555 31.120 127.725 ;
        RECT 9.790 126.835 9.960 127.005 ;
        RECT 9.790 126.475 9.960 126.645 ;
        RECT 9.790 122.085 9.960 122.255 ;
        RECT 9.790 121.725 9.960 121.895 ;
        RECT 9.790 121.365 9.960 121.535 ;
        RECT 9.790 121.005 9.960 121.175 ;
        RECT 6.780 119.965 6.950 120.135 ;
        RECT 6.780 119.605 6.950 119.775 ;
        RECT 6.780 119.245 6.950 119.415 ;
        RECT 6.780 118.885 6.950 119.055 ;
        RECT 6.780 118.525 6.950 118.695 ;
        RECT 6.780 118.165 6.950 118.335 ;
        RECT 6.780 117.805 6.950 117.975 ;
        RECT 6.780 117.445 6.950 117.615 ;
        RECT 6.780 117.085 6.950 117.255 ;
        RECT 6.780 116.725 6.950 116.895 ;
        RECT 6.780 116.365 6.950 116.535 ;
        RECT 6.780 116.005 6.950 116.175 ;
        RECT 6.780 115.645 6.950 115.815 ;
        RECT 6.780 115.285 6.950 115.455 ;
        RECT 6.780 114.925 6.950 115.095 ;
        RECT 6.780 114.565 6.950 114.735 ;
        RECT 6.780 114.205 6.950 114.375 ;
        RECT 9.790 116.615 9.960 116.785 ;
        RECT 9.790 116.255 9.960 116.425 ;
        RECT 9.790 115.895 9.960 116.065 ;
        RECT 9.790 115.535 9.960 115.705 ;
        RECT 9.790 111.145 9.960 111.315 ;
        RECT 9.790 110.785 9.960 110.955 ;
        RECT 9.790 110.425 9.960 110.595 ;
        RECT 9.790 110.065 9.960 110.235 ;
        RECT 9.790 105.675 9.960 105.845 ;
        RECT 15.080 127.195 15.250 127.365 ;
        RECT 15.080 126.835 15.250 127.005 ;
        RECT 15.080 126.475 15.250 126.645 ;
        RECT 15.080 122.085 15.250 122.255 ;
        RECT 15.080 121.725 15.250 121.895 ;
        RECT 15.080 121.365 15.250 121.535 ;
        RECT 15.080 121.005 15.250 121.175 ;
        RECT 15.080 116.615 15.250 116.785 ;
        RECT 15.080 116.255 15.250 116.425 ;
        RECT 15.080 115.895 15.250 116.065 ;
        RECT 15.080 115.535 15.250 115.705 ;
        RECT 15.080 111.145 15.250 111.315 ;
        RECT 15.080 110.785 15.250 110.955 ;
        RECT 15.080 110.425 15.250 110.595 ;
        RECT 15.080 110.065 15.250 110.235 ;
        RECT 15.080 105.675 15.250 105.845 ;
        RECT 20.370 127.195 20.540 127.365 ;
        RECT 20.370 126.835 20.540 127.005 ;
        RECT 20.370 126.475 20.540 126.645 ;
        RECT 20.370 122.085 20.540 122.255 ;
        RECT 20.370 121.725 20.540 121.895 ;
        RECT 20.370 121.365 20.540 121.535 ;
        RECT 20.370 121.005 20.540 121.175 ;
        RECT 20.370 116.615 20.540 116.785 ;
        RECT 20.370 116.255 20.540 116.425 ;
        RECT 20.370 115.895 20.540 116.065 ;
        RECT 20.370 115.535 20.540 115.705 ;
        RECT 20.370 111.145 20.540 111.315 ;
        RECT 20.370 110.785 20.540 110.955 ;
        RECT 20.370 110.425 20.540 110.595 ;
        RECT 20.370 110.065 20.540 110.235 ;
        RECT 20.370 105.675 20.540 105.845 ;
        RECT 36.240 127.555 36.410 127.725 ;
        RECT 25.660 127.195 25.830 127.365 ;
        RECT 25.660 126.835 25.830 127.005 ;
        RECT 25.660 126.475 25.830 126.645 ;
        RECT 25.660 122.085 25.830 122.255 ;
        RECT 25.660 121.725 25.830 121.895 ;
        RECT 25.660 121.365 25.830 121.535 ;
        RECT 25.660 121.005 25.830 121.175 ;
        RECT 25.660 116.615 25.830 116.785 ;
        RECT 25.660 116.255 25.830 116.425 ;
        RECT 25.660 115.895 25.830 116.065 ;
        RECT 25.660 115.535 25.830 115.705 ;
        RECT 25.660 111.145 25.830 111.315 ;
        RECT 25.660 110.785 25.830 110.955 ;
        RECT 25.660 110.425 25.830 110.595 ;
        RECT 25.660 110.065 25.830 110.235 ;
        RECT 25.660 105.675 25.830 105.845 ;
        RECT 30.950 127.195 31.120 127.365 ;
        RECT 30.950 126.835 31.120 127.005 ;
        RECT 30.950 126.475 31.120 126.645 ;
        RECT 30.950 122.085 31.120 122.255 ;
        RECT 30.950 121.725 31.120 121.895 ;
        RECT 30.950 121.365 31.120 121.535 ;
        RECT 30.950 121.005 31.120 121.175 ;
        RECT 30.950 116.615 31.120 116.785 ;
        RECT 30.950 116.255 31.120 116.425 ;
        RECT 30.950 115.895 31.120 116.065 ;
        RECT 30.950 115.535 31.120 115.705 ;
        RECT 30.950 111.145 31.120 111.315 ;
        RECT 30.950 110.785 31.120 110.955 ;
        RECT 30.950 110.425 31.120 110.595 ;
        RECT 30.950 110.065 31.120 110.235 ;
        RECT 9.790 105.315 9.960 105.485 ;
        RECT 9.790 104.955 9.960 105.125 ;
        RECT 15.080 105.315 15.250 105.485 ;
        RECT 9.790 104.595 9.960 104.765 ;
        RECT 15.080 104.955 15.250 105.125 ;
        RECT 20.370 105.315 20.540 105.485 ;
        RECT 15.080 104.595 15.250 104.765 ;
        RECT 20.370 104.955 20.540 105.125 ;
        RECT 30.950 105.675 31.120 105.845 ;
        RECT 36.240 127.195 36.410 127.365 ;
        RECT 36.240 126.835 36.410 127.005 ;
        RECT 36.240 126.475 36.410 126.645 ;
        RECT 36.240 122.085 36.410 122.255 ;
        RECT 36.240 121.725 36.410 121.895 ;
        RECT 36.240 121.365 36.410 121.535 ;
        RECT 36.240 121.005 36.410 121.175 ;
        RECT 36.240 116.615 36.410 116.785 ;
        RECT 36.240 116.255 36.410 116.425 ;
        RECT 36.240 115.895 36.410 116.065 ;
        RECT 36.240 115.535 36.410 115.705 ;
        RECT 36.240 111.145 36.410 111.315 ;
        RECT 36.240 110.785 36.410 110.955 ;
        RECT 36.240 110.425 36.410 110.595 ;
        RECT 36.240 110.065 36.410 110.235 ;
        RECT 25.660 105.315 25.830 105.485 ;
        RECT 25.660 104.955 25.830 105.125 ;
        RECT 30.950 105.315 31.120 105.485 ;
        RECT 30.950 104.955 31.120 105.125 ;
        RECT 36.240 105.675 36.410 105.845 ;
        RECT 36.240 105.315 36.410 105.485 ;
        RECT 20.370 104.595 20.540 104.765 ;
        RECT 25.660 104.595 25.830 104.765 ;
        RECT 30.950 104.595 31.120 104.765 ;
        RECT 36.240 104.955 36.410 105.125 ;
        RECT 36.240 104.595 36.410 104.765 ;
        RECT 42.360 156.775 42.530 156.945 ;
        RECT 42.360 156.415 42.530 156.585 ;
        RECT 47.650 156.775 47.820 156.945 ;
        RECT 52.940 156.775 53.110 156.945 ;
        RECT 58.230 156.775 58.400 156.945 ;
        RECT 63.520 156.775 63.690 156.945 ;
        RECT 42.360 156.055 42.530 156.225 ;
        RECT 42.360 155.695 42.530 155.865 ;
        RECT 42.360 151.305 42.530 151.475 ;
        RECT 42.360 150.945 42.530 151.115 ;
        RECT 42.360 150.585 42.530 150.755 ;
        RECT 42.360 150.225 42.530 150.395 ;
        RECT 42.360 145.835 42.530 146.005 ;
        RECT 42.360 145.475 42.530 145.645 ;
        RECT 42.360 145.115 42.530 145.285 ;
        RECT 42.360 144.755 42.530 144.925 ;
        RECT 42.360 140.365 42.530 140.535 ;
        RECT 42.360 140.005 42.530 140.175 ;
        RECT 42.360 139.645 42.530 139.815 ;
        RECT 42.360 139.285 42.530 139.455 ;
        RECT 42.360 134.895 42.530 135.065 ;
        RECT 47.650 156.415 47.820 156.585 ;
        RECT 47.650 156.055 47.820 156.225 ;
        RECT 47.650 155.695 47.820 155.865 ;
        RECT 47.650 151.305 47.820 151.475 ;
        RECT 47.650 150.945 47.820 151.115 ;
        RECT 47.650 150.585 47.820 150.755 ;
        RECT 47.650 150.225 47.820 150.395 ;
        RECT 47.650 145.835 47.820 146.005 ;
        RECT 47.650 145.475 47.820 145.645 ;
        RECT 47.650 145.115 47.820 145.285 ;
        RECT 47.650 144.755 47.820 144.925 ;
        RECT 47.650 140.365 47.820 140.535 ;
        RECT 47.650 140.005 47.820 140.175 ;
        RECT 47.650 139.645 47.820 139.815 ;
        RECT 47.650 139.285 47.820 139.455 ;
        RECT 47.650 134.895 47.820 135.065 ;
        RECT 52.940 156.415 53.110 156.585 ;
        RECT 52.940 156.055 53.110 156.225 ;
        RECT 52.940 155.695 53.110 155.865 ;
        RECT 52.940 151.305 53.110 151.475 ;
        RECT 52.940 150.945 53.110 151.115 ;
        RECT 52.940 150.585 53.110 150.755 ;
        RECT 52.940 150.225 53.110 150.395 ;
        RECT 52.940 145.835 53.110 146.005 ;
        RECT 52.940 145.475 53.110 145.645 ;
        RECT 52.940 145.115 53.110 145.285 ;
        RECT 52.940 144.755 53.110 144.925 ;
        RECT 52.940 140.365 53.110 140.535 ;
        RECT 52.940 140.005 53.110 140.175 ;
        RECT 52.940 139.645 53.110 139.815 ;
        RECT 52.940 139.285 53.110 139.455 ;
        RECT 52.940 134.895 53.110 135.065 ;
        RECT 68.810 156.775 68.980 156.945 ;
        RECT 58.230 156.415 58.400 156.585 ;
        RECT 58.230 156.055 58.400 156.225 ;
        RECT 58.230 155.695 58.400 155.865 ;
        RECT 58.230 151.305 58.400 151.475 ;
        RECT 58.230 150.945 58.400 151.115 ;
        RECT 58.230 150.585 58.400 150.755 ;
        RECT 58.230 150.225 58.400 150.395 ;
        RECT 58.230 145.835 58.400 146.005 ;
        RECT 58.230 145.475 58.400 145.645 ;
        RECT 58.230 145.115 58.400 145.285 ;
        RECT 58.230 144.755 58.400 144.925 ;
        RECT 58.230 140.365 58.400 140.535 ;
        RECT 58.230 140.005 58.400 140.175 ;
        RECT 58.230 139.645 58.400 139.815 ;
        RECT 58.230 139.285 58.400 139.455 ;
        RECT 58.230 134.895 58.400 135.065 ;
        RECT 63.520 156.415 63.690 156.585 ;
        RECT 63.520 156.055 63.690 156.225 ;
        RECT 63.520 155.695 63.690 155.865 ;
        RECT 63.520 151.305 63.690 151.475 ;
        RECT 63.520 150.945 63.690 151.115 ;
        RECT 63.520 150.585 63.690 150.755 ;
        RECT 63.520 150.225 63.690 150.395 ;
        RECT 63.520 145.835 63.690 146.005 ;
        RECT 63.520 145.475 63.690 145.645 ;
        RECT 63.520 145.115 63.690 145.285 ;
        RECT 63.520 144.755 63.690 144.925 ;
        RECT 63.520 140.365 63.690 140.535 ;
        RECT 63.520 140.005 63.690 140.175 ;
        RECT 63.520 139.645 63.690 139.815 ;
        RECT 63.520 139.285 63.690 139.455 ;
        RECT 42.360 134.535 42.530 134.705 ;
        RECT 42.360 134.175 42.530 134.345 ;
        RECT 47.650 134.535 47.820 134.705 ;
        RECT 42.360 133.815 42.530 133.985 ;
        RECT 47.650 134.175 47.820 134.345 ;
        RECT 52.940 134.535 53.110 134.705 ;
        RECT 47.650 133.815 47.820 133.985 ;
        RECT 52.940 134.175 53.110 134.345 ;
        RECT 63.520 134.895 63.690 135.065 ;
        RECT 68.810 156.415 68.980 156.585 ;
        RECT 68.810 156.055 68.980 156.225 ;
        RECT 68.810 155.695 68.980 155.865 ;
        RECT 68.810 151.305 68.980 151.475 ;
        RECT 68.810 150.945 68.980 151.115 ;
        RECT 68.810 150.585 68.980 150.755 ;
        RECT 68.810 150.225 68.980 150.395 ;
        RECT 68.810 145.835 68.980 146.005 ;
        RECT 68.810 145.475 68.980 145.645 ;
        RECT 68.810 145.115 68.980 145.285 ;
        RECT 68.810 144.755 68.980 144.925 ;
        RECT 68.810 140.365 68.980 140.535 ;
        RECT 68.810 140.005 68.980 140.175 ;
        RECT 68.810 139.645 68.980 139.815 ;
        RECT 68.810 139.285 68.980 139.455 ;
        RECT 58.230 134.535 58.400 134.705 ;
        RECT 58.230 134.175 58.400 134.345 ;
        RECT 68.810 134.895 68.980 135.065 ;
        RECT 63.520 134.535 63.690 134.705 ;
        RECT 63.520 134.175 63.690 134.345 ;
        RECT 68.810 134.535 68.980 134.705 ;
        RECT 52.940 133.815 53.110 133.985 ;
        RECT 58.230 133.815 58.400 133.985 ;
        RECT 63.520 133.815 63.690 133.985 ;
        RECT 68.810 134.175 68.980 134.345 ;
        RECT 68.810 133.815 68.980 133.985 ;
        RECT 74.890 185.985 75.060 186.155 ;
        RECT 74.890 185.625 75.060 185.795 ;
        RECT 80.180 185.985 80.350 186.155 ;
        RECT 85.470 185.985 85.640 186.155 ;
        RECT 90.760 185.985 90.930 186.155 ;
        RECT 96.050 185.985 96.220 186.155 ;
        RECT 74.890 185.265 75.060 185.435 ;
        RECT 74.890 184.905 75.060 185.075 ;
        RECT 74.890 180.515 75.060 180.685 ;
        RECT 74.890 180.155 75.060 180.325 ;
        RECT 74.890 179.795 75.060 179.965 ;
        RECT 74.890 179.435 75.060 179.605 ;
        RECT 74.890 175.045 75.060 175.215 ;
        RECT 74.890 174.685 75.060 174.855 ;
        RECT 74.890 174.325 75.060 174.495 ;
        RECT 74.890 173.965 75.060 174.135 ;
        RECT 74.890 169.575 75.060 169.745 ;
        RECT 74.890 169.215 75.060 169.385 ;
        RECT 74.890 168.855 75.060 169.025 ;
        RECT 74.890 168.495 75.060 168.665 ;
        RECT 74.890 164.105 75.060 164.275 ;
        RECT 80.180 185.625 80.350 185.795 ;
        RECT 80.180 185.265 80.350 185.435 ;
        RECT 80.180 184.905 80.350 185.075 ;
        RECT 80.180 180.515 80.350 180.685 ;
        RECT 80.180 180.155 80.350 180.325 ;
        RECT 80.180 179.795 80.350 179.965 ;
        RECT 80.180 179.435 80.350 179.605 ;
        RECT 80.180 175.045 80.350 175.215 ;
        RECT 80.180 174.685 80.350 174.855 ;
        RECT 80.180 174.325 80.350 174.495 ;
        RECT 80.180 173.965 80.350 174.135 ;
        RECT 80.180 169.575 80.350 169.745 ;
        RECT 80.180 169.215 80.350 169.385 ;
        RECT 80.180 168.855 80.350 169.025 ;
        RECT 80.180 168.495 80.350 168.665 ;
        RECT 80.180 164.105 80.350 164.275 ;
        RECT 85.470 185.625 85.640 185.795 ;
        RECT 85.470 185.265 85.640 185.435 ;
        RECT 85.470 184.905 85.640 185.075 ;
        RECT 85.470 180.515 85.640 180.685 ;
        RECT 85.470 180.155 85.640 180.325 ;
        RECT 85.470 179.795 85.640 179.965 ;
        RECT 85.470 179.435 85.640 179.605 ;
        RECT 85.470 175.045 85.640 175.215 ;
        RECT 85.470 174.685 85.640 174.855 ;
        RECT 85.470 174.325 85.640 174.495 ;
        RECT 85.470 173.965 85.640 174.135 ;
        RECT 85.470 169.575 85.640 169.745 ;
        RECT 85.470 169.215 85.640 169.385 ;
        RECT 85.470 168.855 85.640 169.025 ;
        RECT 85.470 168.495 85.640 168.665 ;
        RECT 85.470 164.105 85.640 164.275 ;
        RECT 101.340 185.985 101.510 186.155 ;
        RECT 90.760 185.625 90.930 185.795 ;
        RECT 90.760 185.265 90.930 185.435 ;
        RECT 90.760 184.905 90.930 185.075 ;
        RECT 90.760 180.515 90.930 180.685 ;
        RECT 90.760 180.155 90.930 180.325 ;
        RECT 90.760 179.795 90.930 179.965 ;
        RECT 90.760 179.435 90.930 179.605 ;
        RECT 90.760 175.045 90.930 175.215 ;
        RECT 90.760 174.685 90.930 174.855 ;
        RECT 90.760 174.325 90.930 174.495 ;
        RECT 90.760 173.965 90.930 174.135 ;
        RECT 90.760 169.575 90.930 169.745 ;
        RECT 90.760 169.215 90.930 169.385 ;
        RECT 90.760 168.855 90.930 169.025 ;
        RECT 90.760 168.495 90.930 168.665 ;
        RECT 90.760 164.105 90.930 164.275 ;
        RECT 96.050 185.625 96.220 185.795 ;
        RECT 96.050 185.265 96.220 185.435 ;
        RECT 96.050 184.905 96.220 185.075 ;
        RECT 96.050 180.515 96.220 180.685 ;
        RECT 96.050 180.155 96.220 180.325 ;
        RECT 96.050 179.795 96.220 179.965 ;
        RECT 96.050 179.435 96.220 179.605 ;
        RECT 96.050 175.045 96.220 175.215 ;
        RECT 96.050 174.685 96.220 174.855 ;
        RECT 96.050 174.325 96.220 174.495 ;
        RECT 96.050 173.965 96.220 174.135 ;
        RECT 96.050 169.575 96.220 169.745 ;
        RECT 96.050 169.215 96.220 169.385 ;
        RECT 96.050 168.855 96.220 169.025 ;
        RECT 96.050 168.495 96.220 168.665 ;
        RECT 74.890 163.745 75.060 163.915 ;
        RECT 74.890 163.385 75.060 163.555 ;
        RECT 80.180 163.745 80.350 163.915 ;
        RECT 74.890 163.025 75.060 163.195 ;
        RECT 80.180 163.385 80.350 163.555 ;
        RECT 85.470 163.745 85.640 163.915 ;
        RECT 80.180 163.025 80.350 163.195 ;
        RECT 85.470 163.385 85.640 163.555 ;
        RECT 96.050 164.105 96.220 164.275 ;
        RECT 101.340 185.625 101.510 185.795 ;
        RECT 101.340 185.265 101.510 185.435 ;
        RECT 101.340 184.905 101.510 185.075 ;
        RECT 101.340 180.515 101.510 180.685 ;
        RECT 101.340 180.155 101.510 180.325 ;
        RECT 101.340 179.795 101.510 179.965 ;
        RECT 101.340 179.435 101.510 179.605 ;
        RECT 101.340 175.045 101.510 175.215 ;
        RECT 101.340 174.685 101.510 174.855 ;
        RECT 101.340 174.325 101.510 174.495 ;
        RECT 101.340 173.965 101.510 174.135 ;
        RECT 101.340 169.575 101.510 169.745 ;
        RECT 101.340 169.215 101.510 169.385 ;
        RECT 101.340 168.855 101.510 169.025 ;
        RECT 101.340 168.495 101.510 168.665 ;
        RECT 90.760 163.745 90.930 163.915 ;
        RECT 90.760 163.385 90.930 163.555 ;
        RECT 96.050 163.745 96.220 163.915 ;
        RECT 96.050 163.385 96.220 163.555 ;
        RECT 85.470 163.025 85.640 163.195 ;
        RECT 90.760 163.025 90.930 163.195 ;
        RECT 96.050 163.025 96.220 163.195 ;
        RECT 101.340 164.105 101.510 164.275 ;
        RECT 101.340 163.745 101.510 163.915 ;
        RECT 104.330 178.315 104.500 178.485 ;
        RECT 104.330 177.955 104.500 178.125 ;
        RECT 104.330 177.595 104.500 177.765 ;
        RECT 104.330 177.235 104.500 177.405 ;
        RECT 104.330 176.875 104.500 177.045 ;
        RECT 104.330 176.515 104.500 176.685 ;
        RECT 104.330 176.155 104.500 176.325 ;
        RECT 104.330 175.795 104.500 175.965 ;
        RECT 104.330 175.435 104.500 175.605 ;
        RECT 104.330 175.075 104.500 175.245 ;
        RECT 104.330 174.715 104.500 174.885 ;
        RECT 104.330 174.355 104.500 174.525 ;
        RECT 104.330 173.995 104.500 174.165 ;
        RECT 104.330 173.635 104.500 173.805 ;
        RECT 104.330 173.275 104.500 173.445 ;
        RECT 104.330 172.915 104.500 173.085 ;
        RECT 104.330 172.555 104.500 172.725 ;
        RECT 101.340 163.385 101.510 163.555 ;
        RECT 101.340 163.025 101.510 163.195 ;
        RECT 71.880 149.225 72.050 149.395 ;
        RECT 71.880 148.865 72.050 149.035 ;
        RECT 71.880 148.505 72.050 148.675 ;
        RECT 71.880 148.145 72.050 148.315 ;
        RECT 71.880 147.785 72.050 147.955 ;
        RECT 71.880 147.425 72.050 147.595 ;
        RECT 71.880 147.065 72.050 147.235 ;
        RECT 71.880 146.705 72.050 146.875 ;
        RECT 71.880 146.345 72.050 146.515 ;
        RECT 71.880 145.985 72.050 146.155 ;
        RECT 71.880 145.625 72.050 145.795 ;
        RECT 71.880 145.265 72.050 145.435 ;
        RECT 71.880 144.905 72.050 145.075 ;
        RECT 71.880 144.545 72.050 144.715 ;
        RECT 71.880 144.185 72.050 144.355 ;
        RECT 71.880 143.825 72.050 143.995 ;
        RECT 71.880 143.465 72.050 143.635 ;
        RECT 39.350 120.005 39.520 120.175 ;
        RECT 39.350 119.645 39.520 119.815 ;
        RECT 39.350 119.285 39.520 119.455 ;
        RECT 39.350 118.925 39.520 119.095 ;
        RECT 39.350 118.565 39.520 118.735 ;
        RECT 39.350 118.205 39.520 118.375 ;
        RECT 39.350 117.845 39.520 118.015 ;
        RECT 39.350 117.485 39.520 117.655 ;
        RECT 39.350 117.125 39.520 117.295 ;
        RECT 39.350 116.765 39.520 116.935 ;
        RECT 39.350 116.405 39.520 116.575 ;
        RECT 39.350 116.045 39.520 116.215 ;
        RECT 39.350 115.685 39.520 115.855 ;
        RECT 39.350 115.325 39.520 115.495 ;
        RECT 39.350 114.965 39.520 115.135 ;
        RECT 39.350 114.605 39.520 114.775 ;
        RECT 39.350 114.245 39.520 114.415 ;
        RECT 9.790 98.235 9.960 98.405 ;
        RECT 9.790 97.875 9.960 98.045 ;
        RECT 15.080 98.235 15.250 98.405 ;
        RECT 20.370 98.235 20.540 98.405 ;
        RECT 25.660 98.235 25.830 98.405 ;
        RECT 30.950 98.235 31.120 98.405 ;
        RECT 9.790 97.515 9.960 97.685 ;
        RECT 9.790 97.155 9.960 97.325 ;
        RECT 9.790 92.765 9.960 92.935 ;
        RECT 9.790 92.405 9.960 92.575 ;
        RECT 9.790 92.045 9.960 92.215 ;
        RECT 9.790 91.685 9.960 91.855 ;
        RECT 6.780 90.645 6.950 90.815 ;
        RECT 6.780 90.285 6.950 90.455 ;
        RECT 6.780 89.925 6.950 90.095 ;
        RECT 6.780 89.565 6.950 89.735 ;
        RECT 6.780 89.205 6.950 89.375 ;
        RECT 6.780 88.845 6.950 89.015 ;
        RECT 6.780 88.485 6.950 88.655 ;
        RECT 6.780 88.125 6.950 88.295 ;
        RECT 6.780 87.765 6.950 87.935 ;
        RECT 6.780 87.405 6.950 87.575 ;
        RECT 6.780 87.045 6.950 87.215 ;
        RECT 6.780 86.685 6.950 86.855 ;
        RECT 6.780 86.325 6.950 86.495 ;
        RECT 6.780 85.965 6.950 86.135 ;
        RECT 6.780 85.605 6.950 85.775 ;
        RECT 6.780 85.245 6.950 85.415 ;
        RECT 6.780 84.885 6.950 85.055 ;
        RECT 9.790 87.295 9.960 87.465 ;
        RECT 9.790 86.935 9.960 87.105 ;
        RECT 9.790 86.575 9.960 86.745 ;
        RECT 9.790 86.215 9.960 86.385 ;
        RECT 9.790 81.825 9.960 81.995 ;
        RECT 9.790 81.465 9.960 81.635 ;
        RECT 9.790 81.105 9.960 81.275 ;
        RECT 9.790 80.745 9.960 80.915 ;
        RECT 9.790 76.355 9.960 76.525 ;
        RECT 15.080 97.875 15.250 98.045 ;
        RECT 15.080 97.515 15.250 97.685 ;
        RECT 15.080 97.155 15.250 97.325 ;
        RECT 15.080 92.765 15.250 92.935 ;
        RECT 15.080 92.405 15.250 92.575 ;
        RECT 15.080 92.045 15.250 92.215 ;
        RECT 15.080 91.685 15.250 91.855 ;
        RECT 15.080 87.295 15.250 87.465 ;
        RECT 15.080 86.935 15.250 87.105 ;
        RECT 15.080 86.575 15.250 86.745 ;
        RECT 15.080 86.215 15.250 86.385 ;
        RECT 15.080 81.825 15.250 81.995 ;
        RECT 15.080 81.465 15.250 81.635 ;
        RECT 15.080 81.105 15.250 81.275 ;
        RECT 15.080 80.745 15.250 80.915 ;
        RECT 15.080 76.355 15.250 76.525 ;
        RECT 20.370 97.875 20.540 98.045 ;
        RECT 20.370 97.515 20.540 97.685 ;
        RECT 20.370 97.155 20.540 97.325 ;
        RECT 20.370 92.765 20.540 92.935 ;
        RECT 20.370 92.405 20.540 92.575 ;
        RECT 20.370 92.045 20.540 92.215 ;
        RECT 20.370 91.685 20.540 91.855 ;
        RECT 20.370 87.295 20.540 87.465 ;
        RECT 20.370 86.935 20.540 87.105 ;
        RECT 20.370 86.575 20.540 86.745 ;
        RECT 20.370 86.215 20.540 86.385 ;
        RECT 20.370 81.825 20.540 81.995 ;
        RECT 20.370 81.465 20.540 81.635 ;
        RECT 20.370 81.105 20.540 81.275 ;
        RECT 20.370 80.745 20.540 80.915 ;
        RECT 20.370 76.355 20.540 76.525 ;
        RECT 36.240 98.235 36.410 98.405 ;
        RECT 25.660 97.875 25.830 98.045 ;
        RECT 25.660 97.515 25.830 97.685 ;
        RECT 25.660 97.155 25.830 97.325 ;
        RECT 25.660 92.765 25.830 92.935 ;
        RECT 25.660 92.405 25.830 92.575 ;
        RECT 25.660 92.045 25.830 92.215 ;
        RECT 25.660 91.685 25.830 91.855 ;
        RECT 25.660 87.295 25.830 87.465 ;
        RECT 25.660 86.935 25.830 87.105 ;
        RECT 25.660 86.575 25.830 86.745 ;
        RECT 25.660 86.215 25.830 86.385 ;
        RECT 25.660 81.825 25.830 81.995 ;
        RECT 25.660 81.465 25.830 81.635 ;
        RECT 25.660 81.105 25.830 81.275 ;
        RECT 25.660 80.745 25.830 80.915 ;
        RECT 25.660 76.355 25.830 76.525 ;
        RECT 30.950 97.875 31.120 98.045 ;
        RECT 30.950 97.515 31.120 97.685 ;
        RECT 30.950 97.155 31.120 97.325 ;
        RECT 30.950 92.765 31.120 92.935 ;
        RECT 30.950 92.405 31.120 92.575 ;
        RECT 30.950 92.045 31.120 92.215 ;
        RECT 30.950 91.685 31.120 91.855 ;
        RECT 30.950 87.295 31.120 87.465 ;
        RECT 30.950 86.935 31.120 87.105 ;
        RECT 30.950 86.575 31.120 86.745 ;
        RECT 30.950 86.215 31.120 86.385 ;
        RECT 30.950 81.825 31.120 81.995 ;
        RECT 30.950 81.465 31.120 81.635 ;
        RECT 30.950 81.105 31.120 81.275 ;
        RECT 30.950 80.745 31.120 80.915 ;
        RECT 9.790 75.995 9.960 76.165 ;
        RECT 9.790 75.635 9.960 75.805 ;
        RECT 15.080 75.995 15.250 76.165 ;
        RECT 9.790 75.275 9.960 75.445 ;
        RECT 15.080 75.635 15.250 75.805 ;
        RECT 20.370 75.995 20.540 76.165 ;
        RECT 15.080 75.275 15.250 75.445 ;
        RECT 20.370 75.635 20.540 75.805 ;
        RECT 30.950 76.355 31.120 76.525 ;
        RECT 36.240 97.875 36.410 98.045 ;
        RECT 36.240 97.515 36.410 97.685 ;
        RECT 36.240 97.155 36.410 97.325 ;
        RECT 36.240 92.765 36.410 92.935 ;
        RECT 36.240 92.405 36.410 92.575 ;
        RECT 36.240 92.045 36.410 92.215 ;
        RECT 36.240 91.685 36.410 91.855 ;
        RECT 36.240 87.295 36.410 87.465 ;
        RECT 36.240 86.935 36.410 87.105 ;
        RECT 36.240 86.575 36.410 86.745 ;
        RECT 36.240 86.215 36.410 86.385 ;
        RECT 36.240 81.825 36.410 81.995 ;
        RECT 36.240 81.465 36.410 81.635 ;
        RECT 36.240 81.105 36.410 81.275 ;
        RECT 36.240 80.745 36.410 80.915 ;
        RECT 25.660 75.995 25.830 76.165 ;
        RECT 25.660 75.635 25.830 75.805 ;
        RECT 30.950 75.995 31.120 76.165 ;
        RECT 30.950 75.635 31.120 75.805 ;
        RECT 36.240 76.355 36.410 76.525 ;
        RECT 36.240 75.995 36.410 76.165 ;
        RECT 20.370 75.275 20.540 75.445 ;
        RECT 25.660 75.275 25.830 75.445 ;
        RECT 30.950 75.275 31.120 75.445 ;
        RECT 36.240 75.635 36.410 75.805 ;
        RECT 36.240 75.275 36.410 75.445 ;
        RECT 42.360 127.595 42.530 127.765 ;
        RECT 42.360 127.235 42.530 127.405 ;
        RECT 47.650 127.595 47.820 127.765 ;
        RECT 52.940 127.595 53.110 127.765 ;
        RECT 58.230 127.595 58.400 127.765 ;
        RECT 63.520 127.595 63.690 127.765 ;
        RECT 42.360 126.875 42.530 127.045 ;
        RECT 42.360 126.515 42.530 126.685 ;
        RECT 42.360 122.125 42.530 122.295 ;
        RECT 42.360 121.765 42.530 121.935 ;
        RECT 42.360 121.405 42.530 121.575 ;
        RECT 42.360 121.045 42.530 121.215 ;
        RECT 42.360 116.655 42.530 116.825 ;
        RECT 42.360 116.295 42.530 116.465 ;
        RECT 42.360 115.935 42.530 116.105 ;
        RECT 42.360 115.575 42.530 115.745 ;
        RECT 42.360 111.185 42.530 111.355 ;
        RECT 42.360 110.825 42.530 110.995 ;
        RECT 42.360 110.465 42.530 110.635 ;
        RECT 42.360 110.105 42.530 110.275 ;
        RECT 42.360 105.715 42.530 105.885 ;
        RECT 47.650 127.235 47.820 127.405 ;
        RECT 47.650 126.875 47.820 127.045 ;
        RECT 47.650 126.515 47.820 126.685 ;
        RECT 47.650 122.125 47.820 122.295 ;
        RECT 47.650 121.765 47.820 121.935 ;
        RECT 47.650 121.405 47.820 121.575 ;
        RECT 47.650 121.045 47.820 121.215 ;
        RECT 47.650 116.655 47.820 116.825 ;
        RECT 47.650 116.295 47.820 116.465 ;
        RECT 47.650 115.935 47.820 116.105 ;
        RECT 47.650 115.575 47.820 115.745 ;
        RECT 47.650 111.185 47.820 111.355 ;
        RECT 47.650 110.825 47.820 110.995 ;
        RECT 47.650 110.465 47.820 110.635 ;
        RECT 47.650 110.105 47.820 110.275 ;
        RECT 47.650 105.715 47.820 105.885 ;
        RECT 52.940 127.235 53.110 127.405 ;
        RECT 52.940 126.875 53.110 127.045 ;
        RECT 52.940 126.515 53.110 126.685 ;
        RECT 52.940 122.125 53.110 122.295 ;
        RECT 52.940 121.765 53.110 121.935 ;
        RECT 52.940 121.405 53.110 121.575 ;
        RECT 52.940 121.045 53.110 121.215 ;
        RECT 52.940 116.655 53.110 116.825 ;
        RECT 52.940 116.295 53.110 116.465 ;
        RECT 52.940 115.935 53.110 116.105 ;
        RECT 52.940 115.575 53.110 115.745 ;
        RECT 52.940 111.185 53.110 111.355 ;
        RECT 52.940 110.825 53.110 110.995 ;
        RECT 52.940 110.465 53.110 110.635 ;
        RECT 52.940 110.105 53.110 110.275 ;
        RECT 52.940 105.715 53.110 105.885 ;
        RECT 68.810 127.595 68.980 127.765 ;
        RECT 58.230 127.235 58.400 127.405 ;
        RECT 58.230 126.875 58.400 127.045 ;
        RECT 58.230 126.515 58.400 126.685 ;
        RECT 58.230 122.125 58.400 122.295 ;
        RECT 58.230 121.765 58.400 121.935 ;
        RECT 58.230 121.405 58.400 121.575 ;
        RECT 58.230 121.045 58.400 121.215 ;
        RECT 58.230 116.655 58.400 116.825 ;
        RECT 58.230 116.295 58.400 116.465 ;
        RECT 58.230 115.935 58.400 116.105 ;
        RECT 58.230 115.575 58.400 115.745 ;
        RECT 58.230 111.185 58.400 111.355 ;
        RECT 58.230 110.825 58.400 110.995 ;
        RECT 58.230 110.465 58.400 110.635 ;
        RECT 58.230 110.105 58.400 110.275 ;
        RECT 58.230 105.715 58.400 105.885 ;
        RECT 63.520 127.235 63.690 127.405 ;
        RECT 63.520 126.875 63.690 127.045 ;
        RECT 63.520 126.515 63.690 126.685 ;
        RECT 63.520 122.125 63.690 122.295 ;
        RECT 63.520 121.765 63.690 121.935 ;
        RECT 63.520 121.405 63.690 121.575 ;
        RECT 63.520 121.045 63.690 121.215 ;
        RECT 63.520 116.655 63.690 116.825 ;
        RECT 63.520 116.295 63.690 116.465 ;
        RECT 63.520 115.935 63.690 116.105 ;
        RECT 63.520 115.575 63.690 115.745 ;
        RECT 63.520 111.185 63.690 111.355 ;
        RECT 63.520 110.825 63.690 110.995 ;
        RECT 63.520 110.465 63.690 110.635 ;
        RECT 63.520 110.105 63.690 110.275 ;
        RECT 42.360 105.355 42.530 105.525 ;
        RECT 42.360 104.995 42.530 105.165 ;
        RECT 47.650 105.355 47.820 105.525 ;
        RECT 42.360 104.635 42.530 104.805 ;
        RECT 47.650 104.995 47.820 105.165 ;
        RECT 52.940 105.355 53.110 105.525 ;
        RECT 47.650 104.635 47.820 104.805 ;
        RECT 52.940 104.995 53.110 105.165 ;
        RECT 63.520 105.715 63.690 105.885 ;
        RECT 68.810 127.235 68.980 127.405 ;
        RECT 68.810 126.875 68.980 127.045 ;
        RECT 68.810 126.515 68.980 126.685 ;
        RECT 68.810 122.125 68.980 122.295 ;
        RECT 68.810 121.765 68.980 121.935 ;
        RECT 68.810 121.405 68.980 121.575 ;
        RECT 68.810 121.045 68.980 121.215 ;
        RECT 68.810 116.655 68.980 116.825 ;
        RECT 68.810 116.295 68.980 116.465 ;
        RECT 68.810 115.935 68.980 116.105 ;
        RECT 68.810 115.575 68.980 115.745 ;
        RECT 68.810 111.185 68.980 111.355 ;
        RECT 68.810 110.825 68.980 110.995 ;
        RECT 68.810 110.465 68.980 110.635 ;
        RECT 68.810 110.105 68.980 110.275 ;
        RECT 58.230 105.355 58.400 105.525 ;
        RECT 58.230 104.995 58.400 105.165 ;
        RECT 68.810 105.715 68.980 105.885 ;
        RECT 63.520 105.355 63.690 105.525 ;
        RECT 63.520 104.995 63.690 105.165 ;
        RECT 68.810 105.355 68.980 105.525 ;
        RECT 52.940 104.635 53.110 104.805 ;
        RECT 58.230 104.635 58.400 104.805 ;
        RECT 63.520 104.635 63.690 104.805 ;
        RECT 68.810 104.995 68.980 105.165 ;
        RECT 68.810 104.635 68.980 104.805 ;
        RECT 74.890 156.815 75.060 156.985 ;
        RECT 74.890 156.455 75.060 156.625 ;
        RECT 80.180 156.815 80.350 156.985 ;
        RECT 85.470 156.815 85.640 156.985 ;
        RECT 90.760 156.815 90.930 156.985 ;
        RECT 96.050 156.815 96.220 156.985 ;
        RECT 74.890 156.095 75.060 156.265 ;
        RECT 74.890 155.735 75.060 155.905 ;
        RECT 74.890 151.345 75.060 151.515 ;
        RECT 74.890 150.985 75.060 151.155 ;
        RECT 74.890 150.625 75.060 150.795 ;
        RECT 74.890 150.265 75.060 150.435 ;
        RECT 74.890 145.875 75.060 146.045 ;
        RECT 74.890 145.515 75.060 145.685 ;
        RECT 74.890 145.155 75.060 145.325 ;
        RECT 74.890 144.795 75.060 144.965 ;
        RECT 74.890 140.405 75.060 140.575 ;
        RECT 74.890 140.045 75.060 140.215 ;
        RECT 74.890 139.685 75.060 139.855 ;
        RECT 74.890 139.325 75.060 139.495 ;
        RECT 74.890 134.935 75.060 135.105 ;
        RECT 80.180 156.455 80.350 156.625 ;
        RECT 80.180 156.095 80.350 156.265 ;
        RECT 80.180 155.735 80.350 155.905 ;
        RECT 80.180 151.345 80.350 151.515 ;
        RECT 80.180 150.985 80.350 151.155 ;
        RECT 80.180 150.625 80.350 150.795 ;
        RECT 80.180 150.265 80.350 150.435 ;
        RECT 80.180 145.875 80.350 146.045 ;
        RECT 80.180 145.515 80.350 145.685 ;
        RECT 80.180 145.155 80.350 145.325 ;
        RECT 80.180 144.795 80.350 144.965 ;
        RECT 80.180 140.405 80.350 140.575 ;
        RECT 80.180 140.045 80.350 140.215 ;
        RECT 80.180 139.685 80.350 139.855 ;
        RECT 80.180 139.325 80.350 139.495 ;
        RECT 80.180 134.935 80.350 135.105 ;
        RECT 85.470 156.455 85.640 156.625 ;
        RECT 85.470 156.095 85.640 156.265 ;
        RECT 85.470 155.735 85.640 155.905 ;
        RECT 85.470 151.345 85.640 151.515 ;
        RECT 85.470 150.985 85.640 151.155 ;
        RECT 85.470 150.625 85.640 150.795 ;
        RECT 85.470 150.265 85.640 150.435 ;
        RECT 85.470 145.875 85.640 146.045 ;
        RECT 85.470 145.515 85.640 145.685 ;
        RECT 85.470 145.155 85.640 145.325 ;
        RECT 85.470 144.795 85.640 144.965 ;
        RECT 85.470 140.405 85.640 140.575 ;
        RECT 85.470 140.045 85.640 140.215 ;
        RECT 85.470 139.685 85.640 139.855 ;
        RECT 85.470 139.325 85.640 139.495 ;
        RECT 85.470 134.935 85.640 135.105 ;
        RECT 101.340 156.815 101.510 156.985 ;
        RECT 90.760 156.455 90.930 156.625 ;
        RECT 90.760 156.095 90.930 156.265 ;
        RECT 90.760 155.735 90.930 155.905 ;
        RECT 90.760 151.345 90.930 151.515 ;
        RECT 90.760 150.985 90.930 151.155 ;
        RECT 90.760 150.625 90.930 150.795 ;
        RECT 90.760 150.265 90.930 150.435 ;
        RECT 90.760 145.875 90.930 146.045 ;
        RECT 90.760 145.515 90.930 145.685 ;
        RECT 90.760 145.155 90.930 145.325 ;
        RECT 90.760 144.795 90.930 144.965 ;
        RECT 90.760 140.405 90.930 140.575 ;
        RECT 90.760 140.045 90.930 140.215 ;
        RECT 90.760 139.685 90.930 139.855 ;
        RECT 90.760 139.325 90.930 139.495 ;
        RECT 90.760 134.935 90.930 135.105 ;
        RECT 96.050 156.455 96.220 156.625 ;
        RECT 96.050 156.095 96.220 156.265 ;
        RECT 96.050 155.735 96.220 155.905 ;
        RECT 96.050 151.345 96.220 151.515 ;
        RECT 96.050 150.985 96.220 151.155 ;
        RECT 96.050 150.625 96.220 150.795 ;
        RECT 96.050 150.265 96.220 150.435 ;
        RECT 96.050 145.875 96.220 146.045 ;
        RECT 96.050 145.515 96.220 145.685 ;
        RECT 96.050 145.155 96.220 145.325 ;
        RECT 96.050 144.795 96.220 144.965 ;
        RECT 96.050 140.405 96.220 140.575 ;
        RECT 96.050 140.045 96.220 140.215 ;
        RECT 96.050 139.685 96.220 139.855 ;
        RECT 96.050 139.325 96.220 139.495 ;
        RECT 74.890 134.575 75.060 134.745 ;
        RECT 74.890 134.215 75.060 134.385 ;
        RECT 80.180 134.575 80.350 134.745 ;
        RECT 74.890 133.855 75.060 134.025 ;
        RECT 80.180 134.215 80.350 134.385 ;
        RECT 85.470 134.575 85.640 134.745 ;
        RECT 80.180 133.855 80.350 134.025 ;
        RECT 85.470 134.215 85.640 134.385 ;
        RECT 96.050 134.935 96.220 135.105 ;
        RECT 101.340 156.455 101.510 156.625 ;
        RECT 101.340 156.095 101.510 156.265 ;
        RECT 101.340 155.735 101.510 155.905 ;
        RECT 101.340 151.345 101.510 151.515 ;
        RECT 101.340 150.985 101.510 151.155 ;
        RECT 101.340 150.625 101.510 150.795 ;
        RECT 101.340 150.265 101.510 150.435 ;
        RECT 101.340 145.875 101.510 146.045 ;
        RECT 101.340 145.515 101.510 145.685 ;
        RECT 101.340 145.155 101.510 145.325 ;
        RECT 101.340 144.795 101.510 144.965 ;
        RECT 101.340 140.405 101.510 140.575 ;
        RECT 101.340 140.045 101.510 140.215 ;
        RECT 101.340 139.685 101.510 139.855 ;
        RECT 101.340 139.325 101.510 139.495 ;
        RECT 90.760 134.575 90.930 134.745 ;
        RECT 90.760 134.215 90.930 134.385 ;
        RECT 96.050 134.575 96.220 134.745 ;
        RECT 96.050 134.215 96.220 134.385 ;
        RECT 101.340 134.935 101.510 135.105 ;
        RECT 101.340 134.575 101.510 134.745 ;
        RECT 85.470 133.855 85.640 134.025 ;
        RECT 90.760 133.855 90.930 134.025 ;
        RECT 96.050 133.855 96.220 134.025 ;
        RECT 101.340 134.215 101.510 134.385 ;
        RECT 104.330 149.145 104.500 149.315 ;
        RECT 104.330 148.785 104.500 148.955 ;
        RECT 104.330 148.425 104.500 148.595 ;
        RECT 104.330 148.065 104.500 148.235 ;
        RECT 104.330 147.705 104.500 147.875 ;
        RECT 104.330 147.345 104.500 147.515 ;
        RECT 104.330 146.985 104.500 147.155 ;
        RECT 104.330 146.625 104.500 146.795 ;
        RECT 104.330 146.265 104.500 146.435 ;
        RECT 104.330 145.905 104.500 146.075 ;
        RECT 104.330 145.545 104.500 145.715 ;
        RECT 104.330 145.185 104.500 145.355 ;
        RECT 104.330 144.825 104.500 144.995 ;
        RECT 104.330 144.465 104.500 144.635 ;
        RECT 104.330 144.105 104.500 144.275 ;
        RECT 104.330 143.745 104.500 143.915 ;
        RECT 104.330 143.385 104.500 143.555 ;
        RECT 101.340 133.855 101.510 134.025 ;
        RECT 71.880 120.045 72.050 120.215 ;
        RECT 71.880 119.685 72.050 119.855 ;
        RECT 71.880 119.325 72.050 119.495 ;
        RECT 71.880 118.965 72.050 119.135 ;
        RECT 71.880 118.605 72.050 118.775 ;
        RECT 71.880 118.245 72.050 118.415 ;
        RECT 71.880 117.885 72.050 118.055 ;
        RECT 71.880 117.525 72.050 117.695 ;
        RECT 71.880 117.165 72.050 117.335 ;
        RECT 71.880 116.805 72.050 116.975 ;
        RECT 71.880 116.445 72.050 116.615 ;
        RECT 71.880 116.085 72.050 116.255 ;
        RECT 71.880 115.725 72.050 115.895 ;
        RECT 71.880 115.365 72.050 115.535 ;
        RECT 71.880 115.005 72.050 115.175 ;
        RECT 71.880 114.645 72.050 114.815 ;
        RECT 71.880 114.285 72.050 114.455 ;
        RECT 39.350 90.685 39.520 90.855 ;
        RECT 39.350 90.325 39.520 90.495 ;
        RECT 39.350 89.965 39.520 90.135 ;
        RECT 39.350 89.605 39.520 89.775 ;
        RECT 39.350 89.245 39.520 89.415 ;
        RECT 39.350 88.885 39.520 89.055 ;
        RECT 39.350 88.525 39.520 88.695 ;
        RECT 39.350 88.165 39.520 88.335 ;
        RECT 39.350 87.805 39.520 87.975 ;
        RECT 39.350 87.445 39.520 87.615 ;
        RECT 39.350 87.085 39.520 87.255 ;
        RECT 39.350 86.725 39.520 86.895 ;
        RECT 39.350 86.365 39.520 86.535 ;
        RECT 39.350 86.005 39.520 86.175 ;
        RECT 39.350 85.645 39.520 85.815 ;
        RECT 39.350 85.285 39.520 85.455 ;
        RECT 39.350 84.925 39.520 85.095 ;
        RECT 9.840 68.955 10.010 69.125 ;
        RECT 9.840 68.595 10.010 68.765 ;
        RECT 15.130 68.955 15.300 69.125 ;
        RECT 20.420 68.955 20.590 69.125 ;
        RECT 25.710 68.955 25.880 69.125 ;
        RECT 31.000 68.955 31.170 69.125 ;
        RECT 9.840 68.235 10.010 68.405 ;
        RECT 9.840 67.875 10.010 68.045 ;
        RECT 9.840 63.485 10.010 63.655 ;
        RECT 9.840 63.125 10.010 63.295 ;
        RECT 9.840 62.765 10.010 62.935 ;
        RECT 9.840 62.405 10.010 62.575 ;
        RECT 6.830 61.365 7.000 61.535 ;
        RECT 6.830 61.005 7.000 61.175 ;
        RECT 6.830 60.645 7.000 60.815 ;
        RECT 6.830 60.285 7.000 60.455 ;
        RECT 6.830 59.925 7.000 60.095 ;
        RECT 6.830 59.565 7.000 59.735 ;
        RECT 6.830 59.205 7.000 59.375 ;
        RECT 6.830 58.845 7.000 59.015 ;
        RECT 6.830 58.485 7.000 58.655 ;
        RECT 6.830 58.125 7.000 58.295 ;
        RECT 6.830 57.765 7.000 57.935 ;
        RECT 6.830 57.405 7.000 57.575 ;
        RECT 6.830 57.045 7.000 57.215 ;
        RECT 6.830 56.685 7.000 56.855 ;
        RECT 6.830 56.325 7.000 56.495 ;
        RECT 6.830 55.965 7.000 56.135 ;
        RECT 6.830 55.605 7.000 55.775 ;
        RECT 9.840 58.015 10.010 58.185 ;
        RECT 9.840 57.655 10.010 57.825 ;
        RECT 9.840 57.295 10.010 57.465 ;
        RECT 9.840 56.935 10.010 57.105 ;
        RECT 9.840 52.545 10.010 52.715 ;
        RECT 9.840 52.185 10.010 52.355 ;
        RECT 9.840 51.825 10.010 51.995 ;
        RECT 9.840 51.465 10.010 51.635 ;
        RECT 9.840 47.075 10.010 47.245 ;
        RECT 15.130 68.595 15.300 68.765 ;
        RECT 15.130 68.235 15.300 68.405 ;
        RECT 15.130 67.875 15.300 68.045 ;
        RECT 15.130 63.485 15.300 63.655 ;
        RECT 15.130 63.125 15.300 63.295 ;
        RECT 15.130 62.765 15.300 62.935 ;
        RECT 15.130 62.405 15.300 62.575 ;
        RECT 15.130 58.015 15.300 58.185 ;
        RECT 15.130 57.655 15.300 57.825 ;
        RECT 15.130 57.295 15.300 57.465 ;
        RECT 15.130 56.935 15.300 57.105 ;
        RECT 15.130 52.545 15.300 52.715 ;
        RECT 15.130 52.185 15.300 52.355 ;
        RECT 15.130 51.825 15.300 51.995 ;
        RECT 15.130 51.465 15.300 51.635 ;
        RECT 15.130 47.075 15.300 47.245 ;
        RECT 20.420 68.595 20.590 68.765 ;
        RECT 20.420 68.235 20.590 68.405 ;
        RECT 20.420 67.875 20.590 68.045 ;
        RECT 20.420 63.485 20.590 63.655 ;
        RECT 20.420 63.125 20.590 63.295 ;
        RECT 20.420 62.765 20.590 62.935 ;
        RECT 20.420 62.405 20.590 62.575 ;
        RECT 20.420 58.015 20.590 58.185 ;
        RECT 20.420 57.655 20.590 57.825 ;
        RECT 20.420 57.295 20.590 57.465 ;
        RECT 20.420 56.935 20.590 57.105 ;
        RECT 20.420 52.545 20.590 52.715 ;
        RECT 20.420 52.185 20.590 52.355 ;
        RECT 20.420 51.825 20.590 51.995 ;
        RECT 20.420 51.465 20.590 51.635 ;
        RECT 20.420 47.075 20.590 47.245 ;
        RECT 36.290 68.955 36.460 69.125 ;
        RECT 25.710 68.595 25.880 68.765 ;
        RECT 25.710 68.235 25.880 68.405 ;
        RECT 25.710 67.875 25.880 68.045 ;
        RECT 25.710 63.485 25.880 63.655 ;
        RECT 25.710 63.125 25.880 63.295 ;
        RECT 25.710 62.765 25.880 62.935 ;
        RECT 25.710 62.405 25.880 62.575 ;
        RECT 25.710 58.015 25.880 58.185 ;
        RECT 25.710 57.655 25.880 57.825 ;
        RECT 25.710 57.295 25.880 57.465 ;
        RECT 25.710 56.935 25.880 57.105 ;
        RECT 25.710 52.545 25.880 52.715 ;
        RECT 25.710 52.185 25.880 52.355 ;
        RECT 25.710 51.825 25.880 51.995 ;
        RECT 25.710 51.465 25.880 51.635 ;
        RECT 25.710 47.075 25.880 47.245 ;
        RECT 31.000 68.595 31.170 68.765 ;
        RECT 31.000 68.235 31.170 68.405 ;
        RECT 31.000 67.875 31.170 68.045 ;
        RECT 31.000 63.485 31.170 63.655 ;
        RECT 31.000 63.125 31.170 63.295 ;
        RECT 31.000 62.765 31.170 62.935 ;
        RECT 31.000 62.405 31.170 62.575 ;
        RECT 31.000 58.015 31.170 58.185 ;
        RECT 31.000 57.655 31.170 57.825 ;
        RECT 31.000 57.295 31.170 57.465 ;
        RECT 31.000 56.935 31.170 57.105 ;
        RECT 31.000 52.545 31.170 52.715 ;
        RECT 31.000 52.185 31.170 52.355 ;
        RECT 31.000 51.825 31.170 51.995 ;
        RECT 31.000 51.465 31.170 51.635 ;
        RECT 9.840 46.715 10.010 46.885 ;
        RECT 9.840 46.355 10.010 46.525 ;
        RECT 15.130 46.715 15.300 46.885 ;
        RECT 9.840 45.995 10.010 46.165 ;
        RECT 15.130 46.355 15.300 46.525 ;
        RECT 20.420 46.715 20.590 46.885 ;
        RECT 15.130 45.995 15.300 46.165 ;
        RECT 20.420 46.355 20.590 46.525 ;
        RECT 31.000 47.075 31.170 47.245 ;
        RECT 36.290 68.595 36.460 68.765 ;
        RECT 36.290 68.235 36.460 68.405 ;
        RECT 36.290 67.875 36.460 68.045 ;
        RECT 36.290 63.485 36.460 63.655 ;
        RECT 36.290 63.125 36.460 63.295 ;
        RECT 36.290 62.765 36.460 62.935 ;
        RECT 36.290 62.405 36.460 62.575 ;
        RECT 36.290 58.015 36.460 58.185 ;
        RECT 36.290 57.655 36.460 57.825 ;
        RECT 36.290 57.295 36.460 57.465 ;
        RECT 36.290 56.935 36.460 57.105 ;
        RECT 36.290 52.545 36.460 52.715 ;
        RECT 36.290 52.185 36.460 52.355 ;
        RECT 36.290 51.825 36.460 51.995 ;
        RECT 36.290 51.465 36.460 51.635 ;
        RECT 25.710 46.715 25.880 46.885 ;
        RECT 25.710 46.355 25.880 46.525 ;
        RECT 31.000 46.715 31.170 46.885 ;
        RECT 31.000 46.355 31.170 46.525 ;
        RECT 36.290 47.075 36.460 47.245 ;
        RECT 36.290 46.715 36.460 46.885 ;
        RECT 20.420 45.995 20.590 46.165 ;
        RECT 25.710 45.995 25.880 46.165 ;
        RECT 31.000 45.995 31.170 46.165 ;
        RECT 36.290 46.355 36.460 46.525 ;
        RECT 36.290 45.995 36.460 46.165 ;
        RECT 42.360 98.275 42.530 98.445 ;
        RECT 42.360 97.915 42.530 98.085 ;
        RECT 47.650 98.275 47.820 98.445 ;
        RECT 52.940 98.275 53.110 98.445 ;
        RECT 58.230 98.275 58.400 98.445 ;
        RECT 63.520 98.275 63.690 98.445 ;
        RECT 42.360 97.555 42.530 97.725 ;
        RECT 42.360 97.195 42.530 97.365 ;
        RECT 42.360 92.805 42.530 92.975 ;
        RECT 42.360 92.445 42.530 92.615 ;
        RECT 42.360 92.085 42.530 92.255 ;
        RECT 42.360 91.725 42.530 91.895 ;
        RECT 42.360 87.335 42.530 87.505 ;
        RECT 42.360 86.975 42.530 87.145 ;
        RECT 42.360 86.615 42.530 86.785 ;
        RECT 42.360 86.255 42.530 86.425 ;
        RECT 42.360 81.865 42.530 82.035 ;
        RECT 42.360 81.505 42.530 81.675 ;
        RECT 42.360 81.145 42.530 81.315 ;
        RECT 42.360 80.785 42.530 80.955 ;
        RECT 42.360 76.395 42.530 76.565 ;
        RECT 47.650 97.915 47.820 98.085 ;
        RECT 47.650 97.555 47.820 97.725 ;
        RECT 47.650 97.195 47.820 97.365 ;
        RECT 47.650 92.805 47.820 92.975 ;
        RECT 47.650 92.445 47.820 92.615 ;
        RECT 47.650 92.085 47.820 92.255 ;
        RECT 47.650 91.725 47.820 91.895 ;
        RECT 47.650 87.335 47.820 87.505 ;
        RECT 47.650 86.975 47.820 87.145 ;
        RECT 47.650 86.615 47.820 86.785 ;
        RECT 47.650 86.255 47.820 86.425 ;
        RECT 47.650 81.865 47.820 82.035 ;
        RECT 47.650 81.505 47.820 81.675 ;
        RECT 47.650 81.145 47.820 81.315 ;
        RECT 47.650 80.785 47.820 80.955 ;
        RECT 47.650 76.395 47.820 76.565 ;
        RECT 52.940 97.915 53.110 98.085 ;
        RECT 52.940 97.555 53.110 97.725 ;
        RECT 52.940 97.195 53.110 97.365 ;
        RECT 52.940 92.805 53.110 92.975 ;
        RECT 52.940 92.445 53.110 92.615 ;
        RECT 52.940 92.085 53.110 92.255 ;
        RECT 52.940 91.725 53.110 91.895 ;
        RECT 52.940 87.335 53.110 87.505 ;
        RECT 52.940 86.975 53.110 87.145 ;
        RECT 52.940 86.615 53.110 86.785 ;
        RECT 52.940 86.255 53.110 86.425 ;
        RECT 52.940 81.865 53.110 82.035 ;
        RECT 52.940 81.505 53.110 81.675 ;
        RECT 52.940 81.145 53.110 81.315 ;
        RECT 52.940 80.785 53.110 80.955 ;
        RECT 52.940 76.395 53.110 76.565 ;
        RECT 68.810 98.275 68.980 98.445 ;
        RECT 58.230 97.915 58.400 98.085 ;
        RECT 58.230 97.555 58.400 97.725 ;
        RECT 58.230 97.195 58.400 97.365 ;
        RECT 58.230 92.805 58.400 92.975 ;
        RECT 58.230 92.445 58.400 92.615 ;
        RECT 58.230 92.085 58.400 92.255 ;
        RECT 58.230 91.725 58.400 91.895 ;
        RECT 58.230 87.335 58.400 87.505 ;
        RECT 58.230 86.975 58.400 87.145 ;
        RECT 58.230 86.615 58.400 86.785 ;
        RECT 58.230 86.255 58.400 86.425 ;
        RECT 58.230 81.865 58.400 82.035 ;
        RECT 58.230 81.505 58.400 81.675 ;
        RECT 58.230 81.145 58.400 81.315 ;
        RECT 58.230 80.785 58.400 80.955 ;
        RECT 58.230 76.395 58.400 76.565 ;
        RECT 63.520 97.915 63.690 98.085 ;
        RECT 63.520 97.555 63.690 97.725 ;
        RECT 63.520 97.195 63.690 97.365 ;
        RECT 63.520 92.805 63.690 92.975 ;
        RECT 63.520 92.445 63.690 92.615 ;
        RECT 63.520 92.085 63.690 92.255 ;
        RECT 63.520 91.725 63.690 91.895 ;
        RECT 63.520 87.335 63.690 87.505 ;
        RECT 63.520 86.975 63.690 87.145 ;
        RECT 63.520 86.615 63.690 86.785 ;
        RECT 63.520 86.255 63.690 86.425 ;
        RECT 63.520 81.865 63.690 82.035 ;
        RECT 63.520 81.505 63.690 81.675 ;
        RECT 63.520 81.145 63.690 81.315 ;
        RECT 63.520 80.785 63.690 80.955 ;
        RECT 42.360 76.035 42.530 76.205 ;
        RECT 42.360 75.675 42.530 75.845 ;
        RECT 47.650 76.035 47.820 76.205 ;
        RECT 42.360 75.315 42.530 75.485 ;
        RECT 47.650 75.675 47.820 75.845 ;
        RECT 52.940 76.035 53.110 76.205 ;
        RECT 47.650 75.315 47.820 75.485 ;
        RECT 52.940 75.675 53.110 75.845 ;
        RECT 63.520 76.395 63.690 76.565 ;
        RECT 68.810 97.915 68.980 98.085 ;
        RECT 68.810 97.555 68.980 97.725 ;
        RECT 68.810 97.195 68.980 97.365 ;
        RECT 68.810 92.805 68.980 92.975 ;
        RECT 68.810 92.445 68.980 92.615 ;
        RECT 68.810 92.085 68.980 92.255 ;
        RECT 68.810 91.725 68.980 91.895 ;
        RECT 68.810 87.335 68.980 87.505 ;
        RECT 68.810 86.975 68.980 87.145 ;
        RECT 68.810 86.615 68.980 86.785 ;
        RECT 68.810 86.255 68.980 86.425 ;
        RECT 68.810 81.865 68.980 82.035 ;
        RECT 68.810 81.505 68.980 81.675 ;
        RECT 68.810 81.145 68.980 81.315 ;
        RECT 68.810 80.785 68.980 80.955 ;
        RECT 58.230 76.035 58.400 76.205 ;
        RECT 58.230 75.675 58.400 75.845 ;
        RECT 68.810 76.395 68.980 76.565 ;
        RECT 63.520 76.035 63.690 76.205 ;
        RECT 63.520 75.675 63.690 75.845 ;
        RECT 68.810 76.035 68.980 76.205 ;
        RECT 52.940 75.315 53.110 75.485 ;
        RECT 58.230 75.315 58.400 75.485 ;
        RECT 63.520 75.315 63.690 75.485 ;
        RECT 68.810 75.675 68.980 75.845 ;
        RECT 68.810 75.315 68.980 75.485 ;
        RECT 74.890 127.635 75.060 127.805 ;
        RECT 74.890 127.275 75.060 127.445 ;
        RECT 80.180 127.635 80.350 127.805 ;
        RECT 85.470 127.635 85.640 127.805 ;
        RECT 90.760 127.635 90.930 127.805 ;
        RECT 96.050 127.635 96.220 127.805 ;
        RECT 74.890 126.915 75.060 127.085 ;
        RECT 74.890 126.555 75.060 126.725 ;
        RECT 74.890 122.165 75.060 122.335 ;
        RECT 74.890 121.805 75.060 121.975 ;
        RECT 74.890 121.445 75.060 121.615 ;
        RECT 74.890 121.085 75.060 121.255 ;
        RECT 74.890 116.695 75.060 116.865 ;
        RECT 74.890 116.335 75.060 116.505 ;
        RECT 74.890 115.975 75.060 116.145 ;
        RECT 74.890 115.615 75.060 115.785 ;
        RECT 74.890 111.225 75.060 111.395 ;
        RECT 74.890 110.865 75.060 111.035 ;
        RECT 74.890 110.505 75.060 110.675 ;
        RECT 74.890 110.145 75.060 110.315 ;
        RECT 74.890 105.755 75.060 105.925 ;
        RECT 80.180 127.275 80.350 127.445 ;
        RECT 80.180 126.915 80.350 127.085 ;
        RECT 80.180 126.555 80.350 126.725 ;
        RECT 80.180 122.165 80.350 122.335 ;
        RECT 80.180 121.805 80.350 121.975 ;
        RECT 80.180 121.445 80.350 121.615 ;
        RECT 80.180 121.085 80.350 121.255 ;
        RECT 80.180 116.695 80.350 116.865 ;
        RECT 80.180 116.335 80.350 116.505 ;
        RECT 80.180 115.975 80.350 116.145 ;
        RECT 80.180 115.615 80.350 115.785 ;
        RECT 80.180 111.225 80.350 111.395 ;
        RECT 80.180 110.865 80.350 111.035 ;
        RECT 80.180 110.505 80.350 110.675 ;
        RECT 80.180 110.145 80.350 110.315 ;
        RECT 80.180 105.755 80.350 105.925 ;
        RECT 85.470 127.275 85.640 127.445 ;
        RECT 85.470 126.915 85.640 127.085 ;
        RECT 85.470 126.555 85.640 126.725 ;
        RECT 85.470 122.165 85.640 122.335 ;
        RECT 85.470 121.805 85.640 121.975 ;
        RECT 85.470 121.445 85.640 121.615 ;
        RECT 85.470 121.085 85.640 121.255 ;
        RECT 85.470 116.695 85.640 116.865 ;
        RECT 85.470 116.335 85.640 116.505 ;
        RECT 85.470 115.975 85.640 116.145 ;
        RECT 85.470 115.615 85.640 115.785 ;
        RECT 85.470 111.225 85.640 111.395 ;
        RECT 85.470 110.865 85.640 111.035 ;
        RECT 85.470 110.505 85.640 110.675 ;
        RECT 85.470 110.145 85.640 110.315 ;
        RECT 85.470 105.755 85.640 105.925 ;
        RECT 101.340 127.635 101.510 127.805 ;
        RECT 90.760 127.275 90.930 127.445 ;
        RECT 90.760 126.915 90.930 127.085 ;
        RECT 90.760 126.555 90.930 126.725 ;
        RECT 90.760 122.165 90.930 122.335 ;
        RECT 90.760 121.805 90.930 121.975 ;
        RECT 90.760 121.445 90.930 121.615 ;
        RECT 90.760 121.085 90.930 121.255 ;
        RECT 90.760 116.695 90.930 116.865 ;
        RECT 90.760 116.335 90.930 116.505 ;
        RECT 90.760 115.975 90.930 116.145 ;
        RECT 90.760 115.615 90.930 115.785 ;
        RECT 90.760 111.225 90.930 111.395 ;
        RECT 90.760 110.865 90.930 111.035 ;
        RECT 90.760 110.505 90.930 110.675 ;
        RECT 90.760 110.145 90.930 110.315 ;
        RECT 90.760 105.755 90.930 105.925 ;
        RECT 96.050 127.275 96.220 127.445 ;
        RECT 96.050 126.915 96.220 127.085 ;
        RECT 96.050 126.555 96.220 126.725 ;
        RECT 96.050 122.165 96.220 122.335 ;
        RECT 96.050 121.805 96.220 121.975 ;
        RECT 96.050 121.445 96.220 121.615 ;
        RECT 96.050 121.085 96.220 121.255 ;
        RECT 96.050 116.695 96.220 116.865 ;
        RECT 96.050 116.335 96.220 116.505 ;
        RECT 96.050 115.975 96.220 116.145 ;
        RECT 96.050 115.615 96.220 115.785 ;
        RECT 96.050 111.225 96.220 111.395 ;
        RECT 96.050 110.865 96.220 111.035 ;
        RECT 96.050 110.505 96.220 110.675 ;
        RECT 96.050 110.145 96.220 110.315 ;
        RECT 74.890 105.395 75.060 105.565 ;
        RECT 74.890 105.035 75.060 105.205 ;
        RECT 80.180 105.395 80.350 105.565 ;
        RECT 74.890 104.675 75.060 104.845 ;
        RECT 80.180 105.035 80.350 105.205 ;
        RECT 85.470 105.395 85.640 105.565 ;
        RECT 80.180 104.675 80.350 104.845 ;
        RECT 85.470 105.035 85.640 105.205 ;
        RECT 96.050 105.755 96.220 105.925 ;
        RECT 101.340 127.275 101.510 127.445 ;
        RECT 101.340 126.915 101.510 127.085 ;
        RECT 101.340 126.555 101.510 126.725 ;
        RECT 101.340 122.165 101.510 122.335 ;
        RECT 101.340 121.805 101.510 121.975 ;
        RECT 101.340 121.445 101.510 121.615 ;
        RECT 101.340 121.085 101.510 121.255 ;
        RECT 101.340 116.695 101.510 116.865 ;
        RECT 101.340 116.335 101.510 116.505 ;
        RECT 101.340 115.975 101.510 116.145 ;
        RECT 101.340 115.615 101.510 115.785 ;
        RECT 101.340 111.225 101.510 111.395 ;
        RECT 101.340 110.865 101.510 111.035 ;
        RECT 101.340 110.505 101.510 110.675 ;
        RECT 101.340 110.145 101.510 110.315 ;
        RECT 90.760 105.395 90.930 105.565 ;
        RECT 90.760 105.035 90.930 105.205 ;
        RECT 96.050 105.395 96.220 105.565 ;
        RECT 96.050 105.035 96.220 105.205 ;
        RECT 85.470 104.675 85.640 104.845 ;
        RECT 90.760 104.675 90.930 104.845 ;
        RECT 96.050 104.675 96.220 104.845 ;
        RECT 101.340 105.755 101.510 105.925 ;
        RECT 101.340 105.395 101.510 105.565 ;
        RECT 101.340 105.035 101.510 105.205 ;
        RECT 101.340 104.675 101.510 104.845 ;
        RECT 104.330 119.965 104.500 120.135 ;
        RECT 104.330 119.605 104.500 119.775 ;
        RECT 104.330 119.245 104.500 119.415 ;
        RECT 104.330 118.885 104.500 119.055 ;
        RECT 104.330 118.525 104.500 118.695 ;
        RECT 104.330 118.165 104.500 118.335 ;
        RECT 104.330 117.805 104.500 117.975 ;
        RECT 104.330 117.445 104.500 117.615 ;
        RECT 104.330 117.085 104.500 117.255 ;
        RECT 104.330 116.725 104.500 116.895 ;
        RECT 104.330 116.365 104.500 116.535 ;
        RECT 104.330 116.005 104.500 116.175 ;
        RECT 104.330 115.645 104.500 115.815 ;
        RECT 104.330 115.285 104.500 115.455 ;
        RECT 104.330 114.925 104.500 115.095 ;
        RECT 104.330 114.565 104.500 114.735 ;
        RECT 104.330 114.205 104.500 114.375 ;
        RECT 71.880 90.725 72.050 90.895 ;
        RECT 71.880 90.365 72.050 90.535 ;
        RECT 71.880 90.005 72.050 90.175 ;
        RECT 71.880 89.645 72.050 89.815 ;
        RECT 71.880 89.285 72.050 89.455 ;
        RECT 71.880 88.925 72.050 89.095 ;
        RECT 71.880 88.565 72.050 88.735 ;
        RECT 71.880 88.205 72.050 88.375 ;
        RECT 71.880 87.845 72.050 88.015 ;
        RECT 71.880 87.485 72.050 87.655 ;
        RECT 71.880 87.125 72.050 87.295 ;
        RECT 71.880 86.765 72.050 86.935 ;
        RECT 71.880 86.405 72.050 86.575 ;
        RECT 71.880 86.045 72.050 86.215 ;
        RECT 71.880 85.685 72.050 85.855 ;
        RECT 71.880 85.325 72.050 85.495 ;
        RECT 71.880 84.965 72.050 85.135 ;
        RECT 39.400 61.405 39.570 61.575 ;
        RECT 39.400 61.045 39.570 61.215 ;
        RECT 39.400 60.685 39.570 60.855 ;
        RECT 39.400 60.325 39.570 60.495 ;
        RECT 39.400 59.965 39.570 60.135 ;
        RECT 39.400 59.605 39.570 59.775 ;
        RECT 39.400 59.245 39.570 59.415 ;
        RECT 39.400 58.885 39.570 59.055 ;
        RECT 39.400 58.525 39.570 58.695 ;
        RECT 39.400 58.165 39.570 58.335 ;
        RECT 39.400 57.805 39.570 57.975 ;
        RECT 39.400 57.445 39.570 57.615 ;
        RECT 39.400 57.085 39.570 57.255 ;
        RECT 39.400 56.725 39.570 56.895 ;
        RECT 39.400 56.365 39.570 56.535 ;
        RECT 39.400 56.005 39.570 56.175 ;
        RECT 39.400 55.645 39.570 55.815 ;
        RECT 9.930 39.415 10.100 39.585 ;
        RECT 9.930 39.055 10.100 39.225 ;
        RECT 15.220 39.415 15.390 39.585 ;
        RECT 20.510 39.415 20.680 39.585 ;
        RECT 25.800 39.415 25.970 39.585 ;
        RECT 31.090 39.415 31.260 39.585 ;
        RECT 9.930 38.695 10.100 38.865 ;
        RECT 9.930 38.335 10.100 38.505 ;
        RECT 15.220 39.055 15.390 39.225 ;
        RECT 15.220 38.695 15.390 38.865 ;
        RECT 15.220 38.335 15.390 38.505 ;
        RECT 9.930 33.945 10.100 34.115 ;
        RECT 9.930 33.585 10.100 33.755 ;
        RECT 9.930 33.225 10.100 33.395 ;
        RECT 9.930 32.865 10.100 33.035 ;
        RECT 15.220 33.945 15.390 34.115 ;
        RECT 15.220 33.585 15.390 33.755 ;
        RECT 15.220 33.225 15.390 33.395 ;
        RECT 15.220 32.865 15.390 33.035 ;
        RECT 6.920 31.825 7.090 31.995 ;
        RECT 6.920 31.465 7.090 31.635 ;
        RECT 6.920 31.105 7.090 31.275 ;
        RECT 6.920 30.745 7.090 30.915 ;
        RECT 6.920 30.385 7.090 30.555 ;
        RECT 6.920 30.025 7.090 30.195 ;
        RECT 6.920 29.665 7.090 29.835 ;
        RECT 6.920 29.305 7.090 29.475 ;
        RECT 6.920 28.945 7.090 29.115 ;
        RECT 6.920 28.585 7.090 28.755 ;
        RECT 6.920 28.225 7.090 28.395 ;
        RECT 6.920 27.865 7.090 28.035 ;
        RECT 6.920 27.505 7.090 27.675 ;
        RECT 6.920 27.145 7.090 27.315 ;
        RECT 6.920 26.785 7.090 26.955 ;
        RECT 6.920 26.425 7.090 26.595 ;
        RECT 6.920 26.065 7.090 26.235 ;
        RECT 9.930 28.475 10.100 28.645 ;
        RECT 9.930 28.115 10.100 28.285 ;
        RECT 9.930 27.755 10.100 27.925 ;
        RECT 9.930 27.395 10.100 27.565 ;
        RECT 15.220 28.475 15.390 28.645 ;
        RECT 15.220 28.115 15.390 28.285 ;
        RECT 15.220 27.755 15.390 27.925 ;
        RECT 15.220 27.395 15.390 27.565 ;
        RECT 9.930 23.005 10.100 23.175 ;
        RECT 9.930 22.645 10.100 22.815 ;
        RECT 9.930 22.285 10.100 22.455 ;
        RECT 9.930 21.925 10.100 22.095 ;
        RECT 15.220 23.005 15.390 23.175 ;
        RECT 15.220 22.645 15.390 22.815 ;
        RECT 15.220 22.285 15.390 22.455 ;
        RECT 15.220 21.925 15.390 22.095 ;
        RECT 9.930 17.535 10.100 17.705 ;
        RECT 15.220 17.535 15.390 17.705 ;
        RECT 20.510 39.055 20.680 39.225 ;
        RECT 20.510 38.695 20.680 38.865 ;
        RECT 20.510 38.335 20.680 38.505 ;
        RECT 20.510 33.945 20.680 34.115 ;
        RECT 20.510 33.585 20.680 33.755 ;
        RECT 20.510 33.225 20.680 33.395 ;
        RECT 20.510 32.865 20.680 33.035 ;
        RECT 20.510 28.475 20.680 28.645 ;
        RECT 20.510 28.115 20.680 28.285 ;
        RECT 20.510 27.755 20.680 27.925 ;
        RECT 20.510 27.395 20.680 27.565 ;
        RECT 20.510 23.005 20.680 23.175 ;
        RECT 20.510 22.645 20.680 22.815 ;
        RECT 20.510 22.285 20.680 22.455 ;
        RECT 20.510 21.925 20.680 22.095 ;
        RECT 20.510 17.535 20.680 17.705 ;
        RECT 36.380 39.415 36.550 39.585 ;
        RECT 25.800 39.055 25.970 39.225 ;
        RECT 25.800 38.695 25.970 38.865 ;
        RECT 25.800 38.335 25.970 38.505 ;
        RECT 25.800 33.945 25.970 34.115 ;
        RECT 25.800 33.585 25.970 33.755 ;
        RECT 25.800 33.225 25.970 33.395 ;
        RECT 25.800 32.865 25.970 33.035 ;
        RECT 25.800 28.475 25.970 28.645 ;
        RECT 25.800 28.115 25.970 28.285 ;
        RECT 25.800 27.755 25.970 27.925 ;
        RECT 25.800 27.395 25.970 27.565 ;
        RECT 25.800 23.005 25.970 23.175 ;
        RECT 25.800 22.645 25.970 22.815 ;
        RECT 25.800 22.285 25.970 22.455 ;
        RECT 25.800 21.925 25.970 22.095 ;
        RECT 25.800 17.535 25.970 17.705 ;
        RECT 31.090 39.055 31.260 39.225 ;
        RECT 31.090 38.695 31.260 38.865 ;
        RECT 36.380 39.055 36.550 39.225 ;
        RECT 31.090 38.335 31.260 38.505 ;
        RECT 31.090 33.945 31.260 34.115 ;
        RECT 31.090 33.585 31.260 33.755 ;
        RECT 31.090 33.225 31.260 33.395 ;
        RECT 31.090 32.865 31.260 33.035 ;
        RECT 31.090 28.475 31.260 28.645 ;
        RECT 31.090 28.115 31.260 28.285 ;
        RECT 31.090 27.755 31.260 27.925 ;
        RECT 31.090 27.395 31.260 27.565 ;
        RECT 31.090 23.005 31.260 23.175 ;
        RECT 31.090 22.645 31.260 22.815 ;
        RECT 31.090 22.285 31.260 22.455 ;
        RECT 31.090 21.925 31.260 22.095 ;
        RECT 9.930 17.175 10.100 17.345 ;
        RECT 9.930 16.815 10.100 16.985 ;
        RECT 15.220 17.175 15.390 17.345 ;
        RECT 9.930 16.455 10.100 16.625 ;
        RECT 15.220 16.815 15.390 16.985 ;
        RECT 20.510 17.175 20.680 17.345 ;
        RECT 15.220 16.455 15.390 16.625 ;
        RECT -97.130 15.015 -96.960 15.185 ;
        RECT -97.130 14.655 -96.960 14.825 ;
        RECT -97.130 14.295 -96.960 14.465 ;
        RECT -97.130 13.935 -96.960 14.105 ;
        RECT -94.550 15.015 -94.380 15.185 ;
        RECT -94.550 14.655 -94.380 14.825 ;
        RECT -94.550 14.295 -94.380 14.465 ;
        RECT -94.550 13.935 -94.380 14.105 ;
        RECT -91.970 15.015 -91.800 15.185 ;
        RECT -91.970 14.655 -91.800 14.825 ;
        RECT -91.970 14.295 -91.800 14.465 ;
        RECT -91.970 13.935 -91.800 14.105 ;
        RECT -89.390 15.015 -89.220 15.185 ;
        RECT -89.390 14.655 -89.220 14.825 ;
        RECT -89.390 14.295 -89.220 14.465 ;
        RECT -89.390 13.935 -89.220 14.105 ;
        RECT -86.810 15.015 -86.640 15.185 ;
        RECT -86.810 14.655 -86.640 14.825 ;
        RECT -86.810 14.295 -86.640 14.465 ;
        RECT -86.810 13.935 -86.640 14.105 ;
        RECT -84.230 15.015 -84.060 15.185 ;
        RECT -84.230 14.655 -84.060 14.825 ;
        RECT -84.230 14.295 -84.060 14.465 ;
        RECT -84.230 13.935 -84.060 14.105 ;
        RECT -81.650 15.015 -81.480 15.185 ;
        RECT -81.650 14.655 -81.480 14.825 ;
        RECT -81.650 14.295 -81.480 14.465 ;
        RECT -81.650 13.935 -81.480 14.105 ;
        RECT -79.070 15.015 -78.900 15.185 ;
        RECT -79.070 14.655 -78.900 14.825 ;
        RECT -79.070 14.295 -78.900 14.465 ;
        RECT -79.070 13.935 -78.900 14.105 ;
        RECT -76.490 15.015 -76.320 15.185 ;
        RECT -76.490 14.655 -76.320 14.825 ;
        RECT -76.490 14.295 -76.320 14.465 ;
        RECT -76.490 13.935 -76.320 14.105 ;
        RECT -73.910 15.015 -73.740 15.185 ;
        RECT -73.910 14.655 -73.740 14.825 ;
        RECT -73.910 14.295 -73.740 14.465 ;
        RECT -73.910 13.935 -73.740 14.105 ;
        RECT -71.330 15.015 -71.160 15.185 ;
        RECT -71.330 14.655 -71.160 14.825 ;
        RECT -71.330 14.295 -71.160 14.465 ;
        RECT -71.330 13.935 -71.160 14.105 ;
        RECT 20.510 16.815 20.680 16.985 ;
        RECT 31.090 17.535 31.260 17.705 ;
        RECT 36.380 38.695 36.550 38.865 ;
        RECT 36.380 38.335 36.550 38.505 ;
        RECT 36.380 33.945 36.550 34.115 ;
        RECT 36.380 33.585 36.550 33.755 ;
        RECT 36.380 33.225 36.550 33.395 ;
        RECT 36.380 32.865 36.550 33.035 ;
        RECT 36.380 28.475 36.550 28.645 ;
        RECT 36.380 28.115 36.550 28.285 ;
        RECT 36.380 27.755 36.550 27.925 ;
        RECT 36.380 27.395 36.550 27.565 ;
        RECT 42.410 68.995 42.580 69.165 ;
        RECT 42.410 68.635 42.580 68.805 ;
        RECT 47.700 68.995 47.870 69.165 ;
        RECT 52.990 68.995 53.160 69.165 ;
        RECT 58.280 68.995 58.450 69.165 ;
        RECT 63.570 68.995 63.740 69.165 ;
        RECT 42.410 68.275 42.580 68.445 ;
        RECT 42.410 67.915 42.580 68.085 ;
        RECT 42.410 63.525 42.580 63.695 ;
        RECT 42.410 63.165 42.580 63.335 ;
        RECT 42.410 62.805 42.580 62.975 ;
        RECT 42.410 62.445 42.580 62.615 ;
        RECT 42.410 58.055 42.580 58.225 ;
        RECT 42.410 57.695 42.580 57.865 ;
        RECT 42.410 57.335 42.580 57.505 ;
        RECT 42.410 56.975 42.580 57.145 ;
        RECT 42.410 52.585 42.580 52.755 ;
        RECT 42.410 52.225 42.580 52.395 ;
        RECT 42.410 51.865 42.580 52.035 ;
        RECT 42.410 51.505 42.580 51.675 ;
        RECT 42.410 47.115 42.580 47.285 ;
        RECT 47.700 68.635 47.870 68.805 ;
        RECT 47.700 68.275 47.870 68.445 ;
        RECT 47.700 67.915 47.870 68.085 ;
        RECT 47.700 63.525 47.870 63.695 ;
        RECT 47.700 63.165 47.870 63.335 ;
        RECT 47.700 62.805 47.870 62.975 ;
        RECT 47.700 62.445 47.870 62.615 ;
        RECT 47.700 58.055 47.870 58.225 ;
        RECT 47.700 57.695 47.870 57.865 ;
        RECT 47.700 57.335 47.870 57.505 ;
        RECT 47.700 56.975 47.870 57.145 ;
        RECT 47.700 52.585 47.870 52.755 ;
        RECT 47.700 52.225 47.870 52.395 ;
        RECT 47.700 51.865 47.870 52.035 ;
        RECT 47.700 51.505 47.870 51.675 ;
        RECT 47.700 47.115 47.870 47.285 ;
        RECT 52.990 68.635 53.160 68.805 ;
        RECT 52.990 68.275 53.160 68.445 ;
        RECT 52.990 67.915 53.160 68.085 ;
        RECT 52.990 63.525 53.160 63.695 ;
        RECT 52.990 63.165 53.160 63.335 ;
        RECT 52.990 62.805 53.160 62.975 ;
        RECT 52.990 62.445 53.160 62.615 ;
        RECT 52.990 58.055 53.160 58.225 ;
        RECT 52.990 57.695 53.160 57.865 ;
        RECT 52.990 57.335 53.160 57.505 ;
        RECT 52.990 56.975 53.160 57.145 ;
        RECT 52.990 52.585 53.160 52.755 ;
        RECT 52.990 52.225 53.160 52.395 ;
        RECT 52.990 51.865 53.160 52.035 ;
        RECT 52.990 51.505 53.160 51.675 ;
        RECT 52.990 47.115 53.160 47.285 ;
        RECT 68.860 68.995 69.030 69.165 ;
        RECT 58.280 68.635 58.450 68.805 ;
        RECT 58.280 68.275 58.450 68.445 ;
        RECT 58.280 67.915 58.450 68.085 ;
        RECT 58.280 63.525 58.450 63.695 ;
        RECT 58.280 63.165 58.450 63.335 ;
        RECT 58.280 62.805 58.450 62.975 ;
        RECT 58.280 62.445 58.450 62.615 ;
        RECT 58.280 58.055 58.450 58.225 ;
        RECT 58.280 57.695 58.450 57.865 ;
        RECT 58.280 57.335 58.450 57.505 ;
        RECT 58.280 56.975 58.450 57.145 ;
        RECT 58.280 52.585 58.450 52.755 ;
        RECT 58.280 52.225 58.450 52.395 ;
        RECT 58.280 51.865 58.450 52.035 ;
        RECT 58.280 51.505 58.450 51.675 ;
        RECT 58.280 47.115 58.450 47.285 ;
        RECT 63.570 68.635 63.740 68.805 ;
        RECT 63.570 68.275 63.740 68.445 ;
        RECT 63.570 67.915 63.740 68.085 ;
        RECT 63.570 63.525 63.740 63.695 ;
        RECT 63.570 63.165 63.740 63.335 ;
        RECT 63.570 62.805 63.740 62.975 ;
        RECT 63.570 62.445 63.740 62.615 ;
        RECT 63.570 58.055 63.740 58.225 ;
        RECT 63.570 57.695 63.740 57.865 ;
        RECT 63.570 57.335 63.740 57.505 ;
        RECT 63.570 56.975 63.740 57.145 ;
        RECT 63.570 52.585 63.740 52.755 ;
        RECT 63.570 52.225 63.740 52.395 ;
        RECT 63.570 51.865 63.740 52.035 ;
        RECT 63.570 51.505 63.740 51.675 ;
        RECT 42.410 46.755 42.580 46.925 ;
        RECT 42.410 46.395 42.580 46.565 ;
        RECT 47.700 46.755 47.870 46.925 ;
        RECT 42.410 46.035 42.580 46.205 ;
        RECT 47.700 46.395 47.870 46.565 ;
        RECT 52.990 46.755 53.160 46.925 ;
        RECT 47.700 46.035 47.870 46.205 ;
        RECT 52.990 46.395 53.160 46.565 ;
        RECT 63.570 47.115 63.740 47.285 ;
        RECT 68.860 68.635 69.030 68.805 ;
        RECT 68.860 68.275 69.030 68.445 ;
        RECT 68.860 67.915 69.030 68.085 ;
        RECT 68.860 63.525 69.030 63.695 ;
        RECT 68.860 63.165 69.030 63.335 ;
        RECT 68.860 62.805 69.030 62.975 ;
        RECT 68.860 62.445 69.030 62.615 ;
        RECT 68.860 58.055 69.030 58.225 ;
        RECT 68.860 57.695 69.030 57.865 ;
        RECT 68.860 57.335 69.030 57.505 ;
        RECT 68.860 56.975 69.030 57.145 ;
        RECT 68.860 52.585 69.030 52.755 ;
        RECT 68.860 52.225 69.030 52.395 ;
        RECT 68.860 51.865 69.030 52.035 ;
        RECT 68.860 51.505 69.030 51.675 ;
        RECT 58.280 46.755 58.450 46.925 ;
        RECT 58.280 46.395 58.450 46.565 ;
        RECT 68.860 47.115 69.030 47.285 ;
        RECT 63.570 46.755 63.740 46.925 ;
        RECT 63.570 46.395 63.740 46.565 ;
        RECT 68.860 46.755 69.030 46.925 ;
        RECT 52.990 46.035 53.160 46.205 ;
        RECT 58.280 46.035 58.450 46.205 ;
        RECT 63.570 46.035 63.740 46.205 ;
        RECT 68.860 46.395 69.030 46.565 ;
        RECT 68.860 46.035 69.030 46.205 ;
        RECT 74.890 98.315 75.060 98.485 ;
        RECT 74.890 97.955 75.060 98.125 ;
        RECT 80.180 98.315 80.350 98.485 ;
        RECT 85.470 98.315 85.640 98.485 ;
        RECT 90.760 98.315 90.930 98.485 ;
        RECT 96.050 98.315 96.220 98.485 ;
        RECT 74.890 97.595 75.060 97.765 ;
        RECT 74.890 97.235 75.060 97.405 ;
        RECT 74.890 92.845 75.060 93.015 ;
        RECT 74.890 92.485 75.060 92.655 ;
        RECT 74.890 92.125 75.060 92.295 ;
        RECT 74.890 91.765 75.060 91.935 ;
        RECT 74.890 87.375 75.060 87.545 ;
        RECT 74.890 87.015 75.060 87.185 ;
        RECT 74.890 86.655 75.060 86.825 ;
        RECT 74.890 86.295 75.060 86.465 ;
        RECT 74.890 81.905 75.060 82.075 ;
        RECT 74.890 81.545 75.060 81.715 ;
        RECT 74.890 81.185 75.060 81.355 ;
        RECT 74.890 80.825 75.060 80.995 ;
        RECT 74.890 76.435 75.060 76.605 ;
        RECT 80.180 97.955 80.350 98.125 ;
        RECT 80.180 97.595 80.350 97.765 ;
        RECT 80.180 97.235 80.350 97.405 ;
        RECT 80.180 92.845 80.350 93.015 ;
        RECT 80.180 92.485 80.350 92.655 ;
        RECT 80.180 92.125 80.350 92.295 ;
        RECT 80.180 91.765 80.350 91.935 ;
        RECT 80.180 87.375 80.350 87.545 ;
        RECT 80.180 87.015 80.350 87.185 ;
        RECT 80.180 86.655 80.350 86.825 ;
        RECT 80.180 86.295 80.350 86.465 ;
        RECT 80.180 81.905 80.350 82.075 ;
        RECT 80.180 81.545 80.350 81.715 ;
        RECT 80.180 81.185 80.350 81.355 ;
        RECT 80.180 80.825 80.350 80.995 ;
        RECT 80.180 76.435 80.350 76.605 ;
        RECT 85.470 97.955 85.640 98.125 ;
        RECT 85.470 97.595 85.640 97.765 ;
        RECT 85.470 97.235 85.640 97.405 ;
        RECT 85.470 92.845 85.640 93.015 ;
        RECT 85.470 92.485 85.640 92.655 ;
        RECT 85.470 92.125 85.640 92.295 ;
        RECT 85.470 91.765 85.640 91.935 ;
        RECT 85.470 87.375 85.640 87.545 ;
        RECT 85.470 87.015 85.640 87.185 ;
        RECT 85.470 86.655 85.640 86.825 ;
        RECT 85.470 86.295 85.640 86.465 ;
        RECT 85.470 81.905 85.640 82.075 ;
        RECT 85.470 81.545 85.640 81.715 ;
        RECT 85.470 81.185 85.640 81.355 ;
        RECT 85.470 80.825 85.640 80.995 ;
        RECT 85.470 76.435 85.640 76.605 ;
        RECT 101.340 98.315 101.510 98.485 ;
        RECT 90.760 97.955 90.930 98.125 ;
        RECT 90.760 97.595 90.930 97.765 ;
        RECT 90.760 97.235 90.930 97.405 ;
        RECT 90.760 92.845 90.930 93.015 ;
        RECT 90.760 92.485 90.930 92.655 ;
        RECT 90.760 92.125 90.930 92.295 ;
        RECT 90.760 91.765 90.930 91.935 ;
        RECT 90.760 87.375 90.930 87.545 ;
        RECT 90.760 87.015 90.930 87.185 ;
        RECT 90.760 86.655 90.930 86.825 ;
        RECT 90.760 86.295 90.930 86.465 ;
        RECT 90.760 81.905 90.930 82.075 ;
        RECT 90.760 81.545 90.930 81.715 ;
        RECT 90.760 81.185 90.930 81.355 ;
        RECT 90.760 80.825 90.930 80.995 ;
        RECT 90.760 76.435 90.930 76.605 ;
        RECT 96.050 97.955 96.220 98.125 ;
        RECT 96.050 97.595 96.220 97.765 ;
        RECT 96.050 97.235 96.220 97.405 ;
        RECT 96.050 92.845 96.220 93.015 ;
        RECT 96.050 92.485 96.220 92.655 ;
        RECT 96.050 92.125 96.220 92.295 ;
        RECT 96.050 91.765 96.220 91.935 ;
        RECT 96.050 87.375 96.220 87.545 ;
        RECT 96.050 87.015 96.220 87.185 ;
        RECT 96.050 86.655 96.220 86.825 ;
        RECT 96.050 86.295 96.220 86.465 ;
        RECT 96.050 81.905 96.220 82.075 ;
        RECT 96.050 81.545 96.220 81.715 ;
        RECT 96.050 81.185 96.220 81.355 ;
        RECT 96.050 80.825 96.220 80.995 ;
        RECT 74.890 76.075 75.060 76.245 ;
        RECT 74.890 75.715 75.060 75.885 ;
        RECT 80.180 76.075 80.350 76.245 ;
        RECT 74.890 75.355 75.060 75.525 ;
        RECT 80.180 75.715 80.350 75.885 ;
        RECT 85.470 76.075 85.640 76.245 ;
        RECT 80.180 75.355 80.350 75.525 ;
        RECT 85.470 75.715 85.640 75.885 ;
        RECT 96.050 76.435 96.220 76.605 ;
        RECT 101.340 97.955 101.510 98.125 ;
        RECT 101.340 97.595 101.510 97.765 ;
        RECT 101.340 97.235 101.510 97.405 ;
        RECT 101.340 92.845 101.510 93.015 ;
        RECT 101.340 92.485 101.510 92.655 ;
        RECT 101.340 92.125 101.510 92.295 ;
        RECT 101.340 91.765 101.510 91.935 ;
        RECT 101.340 87.375 101.510 87.545 ;
        RECT 101.340 87.015 101.510 87.185 ;
        RECT 101.340 86.655 101.510 86.825 ;
        RECT 101.340 86.295 101.510 86.465 ;
        RECT 101.340 81.905 101.510 82.075 ;
        RECT 101.340 81.545 101.510 81.715 ;
        RECT 101.340 81.185 101.510 81.355 ;
        RECT 101.340 80.825 101.510 80.995 ;
        RECT 90.760 76.075 90.930 76.245 ;
        RECT 90.760 75.715 90.930 75.885 ;
        RECT 96.050 76.075 96.220 76.245 ;
        RECT 96.050 75.715 96.220 75.885 ;
        RECT 85.470 75.355 85.640 75.525 ;
        RECT 90.760 75.355 90.930 75.525 ;
        RECT 96.050 75.355 96.220 75.525 ;
        RECT 101.340 76.435 101.510 76.605 ;
        RECT 101.340 76.075 101.510 76.245 ;
        RECT 101.340 75.715 101.510 75.885 ;
        RECT 101.340 75.355 101.510 75.525 ;
        RECT 104.330 90.645 104.500 90.815 ;
        RECT 104.330 90.285 104.500 90.455 ;
        RECT 104.330 89.925 104.500 90.095 ;
        RECT 104.330 89.565 104.500 89.735 ;
        RECT 104.330 89.205 104.500 89.375 ;
        RECT 104.330 88.845 104.500 89.015 ;
        RECT 104.330 88.485 104.500 88.655 ;
        RECT 104.330 88.125 104.500 88.295 ;
        RECT 104.330 87.765 104.500 87.935 ;
        RECT 104.330 87.405 104.500 87.575 ;
        RECT 104.330 87.045 104.500 87.215 ;
        RECT 104.330 86.685 104.500 86.855 ;
        RECT 104.330 86.325 104.500 86.495 ;
        RECT 104.330 85.965 104.500 86.135 ;
        RECT 104.330 85.605 104.500 85.775 ;
        RECT 104.330 85.245 104.500 85.415 ;
        RECT 104.330 84.885 104.500 85.055 ;
        RECT 71.930 61.445 72.100 61.615 ;
        RECT 71.930 61.085 72.100 61.255 ;
        RECT 71.930 60.725 72.100 60.895 ;
        RECT 71.930 60.365 72.100 60.535 ;
        RECT 71.930 60.005 72.100 60.175 ;
        RECT 71.930 59.645 72.100 59.815 ;
        RECT 71.930 59.285 72.100 59.455 ;
        RECT 71.930 58.925 72.100 59.095 ;
        RECT 71.930 58.565 72.100 58.735 ;
        RECT 71.930 58.205 72.100 58.375 ;
        RECT 71.930 57.845 72.100 58.015 ;
        RECT 71.930 57.485 72.100 57.655 ;
        RECT 71.930 57.125 72.100 57.295 ;
        RECT 71.930 56.765 72.100 56.935 ;
        RECT 71.930 56.405 72.100 56.575 ;
        RECT 71.930 56.045 72.100 56.215 ;
        RECT 71.930 55.685 72.100 55.855 ;
        RECT 42.500 39.455 42.670 39.625 ;
        RECT 42.500 39.095 42.670 39.265 ;
        RECT 47.790 39.455 47.960 39.625 ;
        RECT 53.080 39.455 53.250 39.625 ;
        RECT 58.370 39.455 58.540 39.625 ;
        RECT 63.660 39.455 63.830 39.625 ;
        RECT 42.500 38.735 42.670 38.905 ;
        RECT 39.490 31.865 39.660 32.035 ;
        RECT 39.490 31.505 39.660 31.675 ;
        RECT 39.490 31.145 39.660 31.315 ;
        RECT 39.490 30.785 39.660 30.955 ;
        RECT 39.490 30.425 39.660 30.595 ;
        RECT 39.490 30.065 39.660 30.235 ;
        RECT 39.490 29.705 39.660 29.875 ;
        RECT 39.490 29.345 39.660 29.515 ;
        RECT 39.490 28.985 39.660 29.155 ;
        RECT 39.490 28.625 39.660 28.795 ;
        RECT 39.490 28.265 39.660 28.435 ;
        RECT 39.490 27.905 39.660 28.075 ;
        RECT 39.490 27.545 39.660 27.715 ;
        RECT 39.490 27.185 39.660 27.355 ;
        RECT 39.490 26.825 39.660 26.995 ;
        RECT 39.490 26.465 39.660 26.635 ;
        RECT 39.490 26.105 39.660 26.275 ;
        RECT 42.500 38.375 42.670 38.545 ;
        RECT 47.790 39.095 47.960 39.265 ;
        RECT 47.790 38.735 47.960 38.905 ;
        RECT 47.790 38.375 47.960 38.545 ;
        RECT 42.500 33.985 42.670 34.155 ;
        RECT 42.500 33.625 42.670 33.795 ;
        RECT 42.500 33.265 42.670 33.435 ;
        RECT 42.500 32.905 42.670 33.075 ;
        RECT 47.790 33.985 47.960 34.155 ;
        RECT 47.790 33.625 47.960 33.795 ;
        RECT 47.790 33.265 47.960 33.435 ;
        RECT 47.790 32.905 47.960 33.075 ;
        RECT 42.500 28.515 42.670 28.685 ;
        RECT 42.500 28.155 42.670 28.325 ;
        RECT 42.500 27.795 42.670 27.965 ;
        RECT 42.500 27.435 42.670 27.605 ;
        RECT 47.790 28.515 47.960 28.685 ;
        RECT 47.790 28.155 47.960 28.325 ;
        RECT 47.790 27.795 47.960 27.965 ;
        RECT 47.790 27.435 47.960 27.605 ;
        RECT 36.380 23.005 36.550 23.175 ;
        RECT 36.380 22.645 36.550 22.815 ;
        RECT 36.380 22.285 36.550 22.455 ;
        RECT 36.380 21.925 36.550 22.095 ;
        RECT 25.800 17.175 25.970 17.345 ;
        RECT 25.800 16.815 25.970 16.985 ;
        RECT 36.380 17.535 36.550 17.705 ;
        RECT 42.500 23.045 42.670 23.215 ;
        RECT 42.500 22.685 42.670 22.855 ;
        RECT 42.500 22.325 42.670 22.495 ;
        RECT 42.500 21.965 42.670 22.135 ;
        RECT 47.790 23.045 47.960 23.215 ;
        RECT 47.790 22.685 47.960 22.855 ;
        RECT 47.790 22.325 47.960 22.495 ;
        RECT 47.790 21.965 47.960 22.135 ;
        RECT 42.500 17.575 42.670 17.745 ;
        RECT 31.090 17.175 31.260 17.345 ;
        RECT 31.090 16.815 31.260 16.985 ;
        RECT 36.380 17.175 36.550 17.345 ;
        RECT 20.510 16.455 20.680 16.625 ;
        RECT 25.800 16.455 25.970 16.625 ;
        RECT 31.090 16.455 31.260 16.625 ;
        RECT 36.380 16.815 36.550 16.985 ;
        RECT 47.790 17.575 47.960 17.745 ;
        RECT 53.080 39.095 53.250 39.265 ;
        RECT 53.080 38.735 53.250 38.905 ;
        RECT 53.080 38.375 53.250 38.545 ;
        RECT 53.080 33.985 53.250 34.155 ;
        RECT 53.080 33.625 53.250 33.795 ;
        RECT 53.080 33.265 53.250 33.435 ;
        RECT 53.080 32.905 53.250 33.075 ;
        RECT 53.080 28.515 53.250 28.685 ;
        RECT 53.080 28.155 53.250 28.325 ;
        RECT 53.080 27.795 53.250 27.965 ;
        RECT 53.080 27.435 53.250 27.605 ;
        RECT 53.080 23.045 53.250 23.215 ;
        RECT 53.080 22.685 53.250 22.855 ;
        RECT 53.080 22.325 53.250 22.495 ;
        RECT 53.080 21.965 53.250 22.135 ;
        RECT 53.080 17.575 53.250 17.745 ;
        RECT 68.950 39.455 69.120 39.625 ;
        RECT 58.370 39.095 58.540 39.265 ;
        RECT 58.370 38.735 58.540 38.905 ;
        RECT 58.370 38.375 58.540 38.545 ;
        RECT 58.370 33.985 58.540 34.155 ;
        RECT 58.370 33.625 58.540 33.795 ;
        RECT 58.370 33.265 58.540 33.435 ;
        RECT 58.370 32.905 58.540 33.075 ;
        RECT 58.370 28.515 58.540 28.685 ;
        RECT 58.370 28.155 58.540 28.325 ;
        RECT 58.370 27.795 58.540 27.965 ;
        RECT 58.370 27.435 58.540 27.605 ;
        RECT 58.370 23.045 58.540 23.215 ;
        RECT 58.370 22.685 58.540 22.855 ;
        RECT 58.370 22.325 58.540 22.495 ;
        RECT 58.370 21.965 58.540 22.135 ;
        RECT 58.370 17.575 58.540 17.745 ;
        RECT 63.660 39.095 63.830 39.265 ;
        RECT 63.660 38.735 63.830 38.905 ;
        RECT 63.660 38.375 63.830 38.545 ;
        RECT 63.660 33.985 63.830 34.155 ;
        RECT 63.660 33.625 63.830 33.795 ;
        RECT 63.660 33.265 63.830 33.435 ;
        RECT 63.660 32.905 63.830 33.075 ;
        RECT 63.660 28.515 63.830 28.685 ;
        RECT 63.660 28.155 63.830 28.325 ;
        RECT 63.660 27.795 63.830 27.965 ;
        RECT 63.660 27.435 63.830 27.605 ;
        RECT 63.660 23.045 63.830 23.215 ;
        RECT 63.660 22.685 63.830 22.855 ;
        RECT 63.660 22.325 63.830 22.495 ;
        RECT 63.660 21.965 63.830 22.135 ;
        RECT 42.500 17.215 42.670 17.385 ;
        RECT 42.500 16.855 42.670 17.025 ;
        RECT 47.790 17.215 47.960 17.385 ;
        RECT 36.380 16.455 36.550 16.625 ;
        RECT 42.500 16.495 42.670 16.665 ;
        RECT 47.790 16.855 47.960 17.025 ;
        RECT 53.080 17.215 53.250 17.385 ;
        RECT 47.790 16.495 47.960 16.665 ;
        RECT 53.080 16.855 53.250 17.025 ;
        RECT 63.660 17.575 63.830 17.745 ;
        RECT 68.950 39.095 69.120 39.265 ;
        RECT 68.950 38.735 69.120 38.905 ;
        RECT 68.950 38.375 69.120 38.545 ;
        RECT 68.950 33.985 69.120 34.155 ;
        RECT 68.950 33.625 69.120 33.795 ;
        RECT 68.950 33.265 69.120 33.435 ;
        RECT 68.950 32.905 69.120 33.075 ;
        RECT 68.950 28.515 69.120 28.685 ;
        RECT 68.950 28.155 69.120 28.325 ;
        RECT 68.950 27.795 69.120 27.965 ;
        RECT 68.950 27.435 69.120 27.605 ;
        RECT 68.950 23.045 69.120 23.215 ;
        RECT 68.950 22.685 69.120 22.855 ;
        RECT 68.950 22.325 69.120 22.495 ;
        RECT 68.950 21.965 69.120 22.135 ;
        RECT 58.370 17.215 58.540 17.385 ;
        RECT 58.370 16.855 58.540 17.025 ;
        RECT 68.950 17.575 69.120 17.745 ;
        RECT 74.940 69.035 75.110 69.205 ;
        RECT 74.940 68.675 75.110 68.845 ;
        RECT 80.230 69.035 80.400 69.205 ;
        RECT 85.520 69.035 85.690 69.205 ;
        RECT 90.810 69.035 90.980 69.205 ;
        RECT 96.100 69.035 96.270 69.205 ;
        RECT 74.940 68.315 75.110 68.485 ;
        RECT 74.940 67.955 75.110 68.125 ;
        RECT 74.940 63.565 75.110 63.735 ;
        RECT 74.940 63.205 75.110 63.375 ;
        RECT 74.940 62.845 75.110 63.015 ;
        RECT 74.940 62.485 75.110 62.655 ;
        RECT 74.940 58.095 75.110 58.265 ;
        RECT 74.940 57.735 75.110 57.905 ;
        RECT 74.940 57.375 75.110 57.545 ;
        RECT 74.940 57.015 75.110 57.185 ;
        RECT 74.940 52.625 75.110 52.795 ;
        RECT 74.940 52.265 75.110 52.435 ;
        RECT 74.940 51.905 75.110 52.075 ;
        RECT 74.940 51.545 75.110 51.715 ;
        RECT 74.940 47.155 75.110 47.325 ;
        RECT 80.230 68.675 80.400 68.845 ;
        RECT 80.230 68.315 80.400 68.485 ;
        RECT 80.230 67.955 80.400 68.125 ;
        RECT 80.230 63.565 80.400 63.735 ;
        RECT 80.230 63.205 80.400 63.375 ;
        RECT 80.230 62.845 80.400 63.015 ;
        RECT 80.230 62.485 80.400 62.655 ;
        RECT 80.230 58.095 80.400 58.265 ;
        RECT 80.230 57.735 80.400 57.905 ;
        RECT 80.230 57.375 80.400 57.545 ;
        RECT 80.230 57.015 80.400 57.185 ;
        RECT 80.230 52.625 80.400 52.795 ;
        RECT 80.230 52.265 80.400 52.435 ;
        RECT 80.230 51.905 80.400 52.075 ;
        RECT 80.230 51.545 80.400 51.715 ;
        RECT 80.230 47.155 80.400 47.325 ;
        RECT 85.520 68.675 85.690 68.845 ;
        RECT 85.520 68.315 85.690 68.485 ;
        RECT 85.520 67.955 85.690 68.125 ;
        RECT 85.520 63.565 85.690 63.735 ;
        RECT 85.520 63.205 85.690 63.375 ;
        RECT 85.520 62.845 85.690 63.015 ;
        RECT 85.520 62.485 85.690 62.655 ;
        RECT 85.520 58.095 85.690 58.265 ;
        RECT 85.520 57.735 85.690 57.905 ;
        RECT 85.520 57.375 85.690 57.545 ;
        RECT 85.520 57.015 85.690 57.185 ;
        RECT 85.520 52.625 85.690 52.795 ;
        RECT 85.520 52.265 85.690 52.435 ;
        RECT 85.520 51.905 85.690 52.075 ;
        RECT 85.520 51.545 85.690 51.715 ;
        RECT 85.520 47.155 85.690 47.325 ;
        RECT 101.390 69.035 101.560 69.205 ;
        RECT 90.810 68.675 90.980 68.845 ;
        RECT 90.810 68.315 90.980 68.485 ;
        RECT 90.810 67.955 90.980 68.125 ;
        RECT 90.810 63.565 90.980 63.735 ;
        RECT 90.810 63.205 90.980 63.375 ;
        RECT 90.810 62.845 90.980 63.015 ;
        RECT 90.810 62.485 90.980 62.655 ;
        RECT 90.810 58.095 90.980 58.265 ;
        RECT 90.810 57.735 90.980 57.905 ;
        RECT 90.810 57.375 90.980 57.545 ;
        RECT 90.810 57.015 90.980 57.185 ;
        RECT 90.810 52.625 90.980 52.795 ;
        RECT 90.810 52.265 90.980 52.435 ;
        RECT 90.810 51.905 90.980 52.075 ;
        RECT 90.810 51.545 90.980 51.715 ;
        RECT 90.810 47.155 90.980 47.325 ;
        RECT 96.100 68.675 96.270 68.845 ;
        RECT 96.100 68.315 96.270 68.485 ;
        RECT 96.100 67.955 96.270 68.125 ;
        RECT 96.100 63.565 96.270 63.735 ;
        RECT 96.100 63.205 96.270 63.375 ;
        RECT 96.100 62.845 96.270 63.015 ;
        RECT 96.100 62.485 96.270 62.655 ;
        RECT 96.100 58.095 96.270 58.265 ;
        RECT 96.100 57.735 96.270 57.905 ;
        RECT 96.100 57.375 96.270 57.545 ;
        RECT 96.100 57.015 96.270 57.185 ;
        RECT 96.100 52.625 96.270 52.795 ;
        RECT 96.100 52.265 96.270 52.435 ;
        RECT 96.100 51.905 96.270 52.075 ;
        RECT 96.100 51.545 96.270 51.715 ;
        RECT 74.940 46.795 75.110 46.965 ;
        RECT 74.940 46.435 75.110 46.605 ;
        RECT 80.230 46.795 80.400 46.965 ;
        RECT 74.940 46.075 75.110 46.245 ;
        RECT 80.230 46.435 80.400 46.605 ;
        RECT 85.520 46.795 85.690 46.965 ;
        RECT 80.230 46.075 80.400 46.245 ;
        RECT 85.520 46.435 85.690 46.605 ;
        RECT 96.100 47.155 96.270 47.325 ;
        RECT 101.390 68.675 101.560 68.845 ;
        RECT 101.390 68.315 101.560 68.485 ;
        RECT 101.390 67.955 101.560 68.125 ;
        RECT 101.390 63.565 101.560 63.735 ;
        RECT 101.390 63.205 101.560 63.375 ;
        RECT 101.390 62.845 101.560 63.015 ;
        RECT 101.390 62.485 101.560 62.655 ;
        RECT 101.390 58.095 101.560 58.265 ;
        RECT 101.390 57.735 101.560 57.905 ;
        RECT 101.390 57.375 101.560 57.545 ;
        RECT 101.390 57.015 101.560 57.185 ;
        RECT 101.390 52.625 101.560 52.795 ;
        RECT 101.390 52.265 101.560 52.435 ;
        RECT 101.390 51.905 101.560 52.075 ;
        RECT 101.390 51.545 101.560 51.715 ;
        RECT 90.810 46.795 90.980 46.965 ;
        RECT 90.810 46.435 90.980 46.605 ;
        RECT 96.100 46.795 96.270 46.965 ;
        RECT 96.100 46.435 96.270 46.605 ;
        RECT 85.520 46.075 85.690 46.245 ;
        RECT 90.810 46.075 90.980 46.245 ;
        RECT 96.100 46.075 96.270 46.245 ;
        RECT 101.390 47.155 101.560 47.325 ;
        RECT 101.390 46.795 101.560 46.965 ;
        RECT 101.390 46.435 101.560 46.605 ;
        RECT 101.390 46.075 101.560 46.245 ;
        RECT 104.380 61.365 104.550 61.535 ;
        RECT 104.380 61.005 104.550 61.175 ;
        RECT 104.380 60.645 104.550 60.815 ;
        RECT 104.380 60.285 104.550 60.455 ;
        RECT 104.380 59.925 104.550 60.095 ;
        RECT 104.380 59.565 104.550 59.735 ;
        RECT 104.380 59.205 104.550 59.375 ;
        RECT 104.380 58.845 104.550 59.015 ;
        RECT 104.380 58.485 104.550 58.655 ;
        RECT 104.380 58.125 104.550 58.295 ;
        RECT 104.380 57.765 104.550 57.935 ;
        RECT 104.380 57.405 104.550 57.575 ;
        RECT 104.380 57.045 104.550 57.215 ;
        RECT 104.380 56.685 104.550 56.855 ;
        RECT 104.380 56.325 104.550 56.495 ;
        RECT 104.380 55.965 104.550 56.135 ;
        RECT 104.380 55.605 104.550 55.775 ;
        RECT 75.030 39.495 75.200 39.665 ;
        RECT 72.020 31.905 72.190 32.075 ;
        RECT 72.020 31.545 72.190 31.715 ;
        RECT 72.020 31.185 72.190 31.355 ;
        RECT 72.020 30.825 72.190 30.995 ;
        RECT 72.020 30.465 72.190 30.635 ;
        RECT 72.020 30.105 72.190 30.275 ;
        RECT 72.020 29.745 72.190 29.915 ;
        RECT 72.020 29.385 72.190 29.555 ;
        RECT 72.020 29.025 72.190 29.195 ;
        RECT 72.020 28.665 72.190 28.835 ;
        RECT 72.020 28.305 72.190 28.475 ;
        RECT 72.020 27.945 72.190 28.115 ;
        RECT 72.020 27.585 72.190 27.755 ;
        RECT 72.020 27.225 72.190 27.395 ;
        RECT 72.020 26.865 72.190 27.035 ;
        RECT 72.020 26.505 72.190 26.675 ;
        RECT 72.020 26.145 72.190 26.315 ;
        RECT 63.660 17.215 63.830 17.385 ;
        RECT 63.660 16.855 63.830 17.025 ;
        RECT 68.950 17.215 69.120 17.385 ;
        RECT 53.080 16.495 53.250 16.665 ;
        RECT 58.370 16.495 58.540 16.665 ;
        RECT 63.660 16.495 63.830 16.665 ;
        RECT 68.950 16.855 69.120 17.025 ;
        RECT 75.030 39.135 75.200 39.305 ;
        RECT 80.320 39.495 80.490 39.665 ;
        RECT 85.610 39.495 85.780 39.665 ;
        RECT 90.900 39.495 91.070 39.665 ;
        RECT 96.190 39.495 96.360 39.665 ;
        RECT 75.030 38.775 75.200 38.945 ;
        RECT 75.030 38.415 75.200 38.585 ;
        RECT 80.320 39.135 80.490 39.305 ;
        RECT 80.320 38.775 80.490 38.945 ;
        RECT 80.320 38.415 80.490 38.585 ;
        RECT 75.030 34.025 75.200 34.195 ;
        RECT 75.030 33.665 75.200 33.835 ;
        RECT 75.030 33.305 75.200 33.475 ;
        RECT 75.030 32.945 75.200 33.115 ;
        RECT 80.320 34.025 80.490 34.195 ;
        RECT 80.320 33.665 80.490 33.835 ;
        RECT 80.320 33.305 80.490 33.475 ;
        RECT 80.320 32.945 80.490 33.115 ;
        RECT 75.030 28.555 75.200 28.725 ;
        RECT 75.030 28.195 75.200 28.365 ;
        RECT 75.030 27.835 75.200 28.005 ;
        RECT 75.030 27.475 75.200 27.645 ;
        RECT 80.320 28.555 80.490 28.725 ;
        RECT 80.320 28.195 80.490 28.365 ;
        RECT 80.320 27.835 80.490 28.005 ;
        RECT 80.320 27.475 80.490 27.645 ;
        RECT 75.030 23.085 75.200 23.255 ;
        RECT 75.030 22.725 75.200 22.895 ;
        RECT 75.030 22.365 75.200 22.535 ;
        RECT 75.030 22.005 75.200 22.175 ;
        RECT 80.320 23.085 80.490 23.255 ;
        RECT 80.320 22.725 80.490 22.895 ;
        RECT 80.320 22.365 80.490 22.535 ;
        RECT 80.320 22.005 80.490 22.175 ;
        RECT 75.030 17.615 75.200 17.785 ;
        RECT 80.320 17.615 80.490 17.785 ;
        RECT 85.610 39.135 85.780 39.305 ;
        RECT 85.610 38.775 85.780 38.945 ;
        RECT 85.610 38.415 85.780 38.585 ;
        RECT 85.610 34.025 85.780 34.195 ;
        RECT 85.610 33.665 85.780 33.835 ;
        RECT 85.610 33.305 85.780 33.475 ;
        RECT 85.610 32.945 85.780 33.115 ;
        RECT 85.610 28.555 85.780 28.725 ;
        RECT 85.610 28.195 85.780 28.365 ;
        RECT 85.610 27.835 85.780 28.005 ;
        RECT 85.610 27.475 85.780 27.645 ;
        RECT 85.610 23.085 85.780 23.255 ;
        RECT 85.610 22.725 85.780 22.895 ;
        RECT 85.610 22.365 85.780 22.535 ;
        RECT 85.610 22.005 85.780 22.175 ;
        RECT 85.610 17.615 85.780 17.785 ;
        RECT 101.480 39.495 101.650 39.665 ;
        RECT 90.900 39.135 91.070 39.305 ;
        RECT 90.900 38.775 91.070 38.945 ;
        RECT 90.900 38.415 91.070 38.585 ;
        RECT 90.900 34.025 91.070 34.195 ;
        RECT 90.900 33.665 91.070 33.835 ;
        RECT 90.900 33.305 91.070 33.475 ;
        RECT 90.900 32.945 91.070 33.115 ;
        RECT 90.900 28.555 91.070 28.725 ;
        RECT 90.900 28.195 91.070 28.365 ;
        RECT 90.900 27.835 91.070 28.005 ;
        RECT 90.900 27.475 91.070 27.645 ;
        RECT 90.900 23.085 91.070 23.255 ;
        RECT 90.900 22.725 91.070 22.895 ;
        RECT 90.900 22.365 91.070 22.535 ;
        RECT 90.900 22.005 91.070 22.175 ;
        RECT 90.900 17.615 91.070 17.785 ;
        RECT 96.190 39.135 96.360 39.305 ;
        RECT 101.480 39.135 101.650 39.305 ;
        RECT 96.190 38.775 96.360 38.945 ;
        RECT 96.190 38.415 96.360 38.585 ;
        RECT 96.190 34.025 96.360 34.195 ;
        RECT 96.190 33.665 96.360 33.835 ;
        RECT 96.190 33.305 96.360 33.475 ;
        RECT 96.190 32.945 96.360 33.115 ;
        RECT 96.190 28.555 96.360 28.725 ;
        RECT 96.190 28.195 96.360 28.365 ;
        RECT 96.190 27.835 96.360 28.005 ;
        RECT 96.190 27.475 96.360 27.645 ;
        RECT 96.190 23.085 96.360 23.255 ;
        RECT 96.190 22.725 96.360 22.895 ;
        RECT 96.190 22.365 96.360 22.535 ;
        RECT 96.190 22.005 96.360 22.175 ;
        RECT 75.030 17.255 75.200 17.425 ;
        RECT 75.030 16.895 75.200 17.065 ;
        RECT 80.320 17.255 80.490 17.425 ;
        RECT 68.950 16.495 69.120 16.665 ;
        RECT 75.030 16.535 75.200 16.705 ;
        RECT 80.320 16.895 80.490 17.065 ;
        RECT 85.610 17.255 85.780 17.425 ;
        RECT 80.320 16.535 80.490 16.705 ;
        RECT 85.610 16.895 85.780 17.065 ;
        RECT 96.190 17.615 96.360 17.785 ;
        RECT 101.480 38.775 101.650 38.945 ;
        RECT 101.480 38.415 101.650 38.585 ;
        RECT 101.480 34.025 101.650 34.195 ;
        RECT 101.480 33.665 101.650 33.835 ;
        RECT 101.480 33.305 101.650 33.475 ;
        RECT 101.480 32.945 101.650 33.115 ;
        RECT 101.480 28.555 101.650 28.725 ;
        RECT 101.480 28.195 101.650 28.365 ;
        RECT 101.480 27.835 101.650 28.005 ;
        RECT 101.480 27.475 101.650 27.645 ;
        RECT 101.480 23.085 101.650 23.255 ;
        RECT 101.480 22.725 101.650 22.895 ;
        RECT 101.480 22.365 101.650 22.535 ;
        RECT 101.480 22.005 101.650 22.175 ;
        RECT 104.470 31.825 104.640 31.995 ;
        RECT 104.470 31.465 104.640 31.635 ;
        RECT 104.470 31.105 104.640 31.275 ;
        RECT 104.470 30.745 104.640 30.915 ;
        RECT 104.470 30.385 104.640 30.555 ;
        RECT 104.470 30.025 104.640 30.195 ;
        RECT 104.470 29.665 104.640 29.835 ;
        RECT 104.470 29.305 104.640 29.475 ;
        RECT 104.470 28.945 104.640 29.115 ;
        RECT 104.470 28.585 104.640 28.755 ;
        RECT 104.470 28.225 104.640 28.395 ;
        RECT 104.470 27.865 104.640 28.035 ;
        RECT 104.470 27.505 104.640 27.675 ;
        RECT 104.470 27.145 104.640 27.315 ;
        RECT 104.470 26.785 104.640 26.955 ;
        RECT 104.470 26.425 104.640 26.595 ;
        RECT 104.470 26.065 104.640 26.235 ;
        RECT 136.940 207.475 137.110 207.645 ;
        RECT 136.940 207.115 137.110 207.285 ;
        RECT 136.940 206.755 137.110 206.925 ;
        RECT 136.940 206.395 137.110 206.565 ;
        RECT 136.940 206.035 137.110 206.205 ;
        RECT 136.940 205.675 137.110 205.845 ;
        RECT 136.940 205.315 137.110 205.485 ;
        RECT 136.940 204.955 137.110 205.125 ;
        RECT 136.940 204.595 137.110 204.765 ;
        RECT 136.940 204.235 137.110 204.405 ;
        RECT 136.940 203.875 137.110 204.045 ;
        RECT 136.940 203.515 137.110 203.685 ;
        RECT 136.940 203.155 137.110 203.325 ;
        RECT 136.940 202.795 137.110 202.965 ;
        RECT 136.940 202.435 137.110 202.605 ;
        RECT 136.940 202.075 137.110 202.245 ;
        RECT 136.940 201.715 137.110 201.885 ;
        RECT 136.940 178.395 137.110 178.565 ;
        RECT 136.940 178.035 137.110 178.205 ;
        RECT 136.940 177.675 137.110 177.845 ;
        RECT 136.940 177.315 137.110 177.485 ;
        RECT 136.940 176.955 137.110 177.125 ;
        RECT 136.940 176.595 137.110 176.765 ;
        RECT 136.940 176.235 137.110 176.405 ;
        RECT 136.940 175.875 137.110 176.045 ;
        RECT 136.940 175.515 137.110 175.685 ;
        RECT 136.940 175.155 137.110 175.325 ;
        RECT 136.940 174.795 137.110 174.965 ;
        RECT 136.940 174.435 137.110 174.605 ;
        RECT 136.940 174.075 137.110 174.245 ;
        RECT 136.940 173.715 137.110 173.885 ;
        RECT 136.940 173.355 137.110 173.525 ;
        RECT 136.940 172.995 137.110 173.165 ;
        RECT 136.940 172.635 137.110 172.805 ;
        RECT 136.940 149.225 137.110 149.395 ;
        RECT 136.940 148.865 137.110 149.035 ;
        RECT 136.940 148.505 137.110 148.675 ;
        RECT 136.940 148.145 137.110 148.315 ;
        RECT 136.940 147.785 137.110 147.955 ;
        RECT 136.940 147.425 137.110 147.595 ;
        RECT 136.940 147.065 137.110 147.235 ;
        RECT 136.940 146.705 137.110 146.875 ;
        RECT 136.940 146.345 137.110 146.515 ;
        RECT 136.940 145.985 137.110 146.155 ;
        RECT 136.940 145.625 137.110 145.795 ;
        RECT 136.940 145.265 137.110 145.435 ;
        RECT 136.940 144.905 137.110 145.075 ;
        RECT 136.940 144.545 137.110 144.715 ;
        RECT 136.940 144.185 137.110 144.355 ;
        RECT 136.940 143.825 137.110 143.995 ;
        RECT 136.940 143.465 137.110 143.635 ;
        RECT 136.940 120.045 137.110 120.215 ;
        RECT 136.940 119.685 137.110 119.855 ;
        RECT 136.940 119.325 137.110 119.495 ;
        RECT 136.940 118.965 137.110 119.135 ;
        RECT 136.940 118.605 137.110 118.775 ;
        RECT 136.940 118.245 137.110 118.415 ;
        RECT 136.940 117.885 137.110 118.055 ;
        RECT 136.940 117.525 137.110 117.695 ;
        RECT 136.940 117.165 137.110 117.335 ;
        RECT 136.940 116.805 137.110 116.975 ;
        RECT 136.940 116.445 137.110 116.615 ;
        RECT 136.940 116.085 137.110 116.255 ;
        RECT 136.940 115.725 137.110 115.895 ;
        RECT 136.940 115.365 137.110 115.535 ;
        RECT 136.940 115.005 137.110 115.175 ;
        RECT 136.940 114.645 137.110 114.815 ;
        RECT 136.940 114.285 137.110 114.455 ;
        RECT 136.940 90.725 137.110 90.895 ;
        RECT 136.940 90.365 137.110 90.535 ;
        RECT 136.940 90.005 137.110 90.175 ;
        RECT 136.940 89.645 137.110 89.815 ;
        RECT 136.940 89.285 137.110 89.455 ;
        RECT 136.940 88.925 137.110 89.095 ;
        RECT 136.940 88.565 137.110 88.735 ;
        RECT 136.940 88.205 137.110 88.375 ;
        RECT 136.940 87.845 137.110 88.015 ;
        RECT 136.940 87.485 137.110 87.655 ;
        RECT 136.940 87.125 137.110 87.295 ;
        RECT 136.940 86.765 137.110 86.935 ;
        RECT 136.940 86.405 137.110 86.575 ;
        RECT 136.940 86.045 137.110 86.215 ;
        RECT 136.940 85.685 137.110 85.855 ;
        RECT 136.940 85.325 137.110 85.495 ;
        RECT 136.940 84.965 137.110 85.135 ;
        RECT 136.990 61.445 137.160 61.615 ;
        RECT 136.990 61.085 137.160 61.255 ;
        RECT 136.990 60.725 137.160 60.895 ;
        RECT 136.990 60.365 137.160 60.535 ;
        RECT 136.990 60.005 137.160 60.175 ;
        RECT 136.990 59.645 137.160 59.815 ;
        RECT 136.990 59.285 137.160 59.455 ;
        RECT 136.990 58.925 137.160 59.095 ;
        RECT 136.990 58.565 137.160 58.735 ;
        RECT 136.990 58.205 137.160 58.375 ;
        RECT 136.990 57.845 137.160 58.015 ;
        RECT 136.990 57.485 137.160 57.655 ;
        RECT 136.990 57.125 137.160 57.295 ;
        RECT 136.990 56.765 137.160 56.935 ;
        RECT 136.990 56.405 137.160 56.575 ;
        RECT 136.990 56.045 137.160 56.215 ;
        RECT 136.990 55.685 137.160 55.855 ;
        RECT 137.080 31.905 137.250 32.075 ;
        RECT 137.080 31.545 137.250 31.715 ;
        RECT 137.080 31.185 137.250 31.355 ;
        RECT 137.080 30.825 137.250 30.995 ;
        RECT 137.080 30.465 137.250 30.635 ;
        RECT 137.080 30.105 137.250 30.275 ;
        RECT 137.080 29.745 137.250 29.915 ;
        RECT 137.080 29.385 137.250 29.555 ;
        RECT 137.080 29.025 137.250 29.195 ;
        RECT 137.080 28.665 137.250 28.835 ;
        RECT 137.080 28.305 137.250 28.475 ;
        RECT 137.080 27.945 137.250 28.115 ;
        RECT 137.080 27.585 137.250 27.755 ;
        RECT 137.080 27.225 137.250 27.395 ;
        RECT 137.080 26.865 137.250 27.035 ;
        RECT 137.080 26.505 137.250 26.675 ;
        RECT 137.080 26.145 137.250 26.315 ;
        RECT 90.900 17.255 91.070 17.425 ;
        RECT 90.900 16.895 91.070 17.065 ;
        RECT 101.480 17.615 101.650 17.785 ;
        RECT 204.950 214.015 205.120 214.185 ;
        RECT 210.240 214.735 210.410 214.905 ;
        RECT 210.240 214.375 210.410 214.545 ;
        RECT 210.240 214.015 210.410 214.185 ;
        RECT 169.490 207.505 169.660 207.675 ;
        RECT 169.490 207.145 169.660 207.315 ;
        RECT 169.490 206.785 169.660 206.955 ;
        RECT 169.490 206.425 169.660 206.595 ;
        RECT 169.490 206.065 169.660 206.235 ;
        RECT 169.490 205.705 169.660 205.875 ;
        RECT 169.490 205.345 169.660 205.515 ;
        RECT 169.490 204.985 169.660 205.155 ;
        RECT 169.490 204.625 169.660 204.795 ;
        RECT 169.490 204.265 169.660 204.435 ;
        RECT 169.490 203.905 169.660 204.075 ;
        RECT 169.490 203.545 169.660 203.715 ;
        RECT 169.490 203.185 169.660 203.355 ;
        RECT 169.490 202.825 169.660 202.995 ;
        RECT 169.490 202.465 169.660 202.635 ;
        RECT 169.490 202.105 169.660 202.275 ;
        RECT 169.490 201.745 169.660 201.915 ;
        RECT 169.490 178.425 169.660 178.595 ;
        RECT 169.490 178.065 169.660 178.235 ;
        RECT 169.490 177.705 169.660 177.875 ;
        RECT 169.490 177.345 169.660 177.515 ;
        RECT 169.490 176.985 169.660 177.155 ;
        RECT 169.490 176.625 169.660 176.795 ;
        RECT 169.490 176.265 169.660 176.435 ;
        RECT 169.490 175.905 169.660 176.075 ;
        RECT 169.490 175.545 169.660 175.715 ;
        RECT 169.490 175.185 169.660 175.355 ;
        RECT 169.490 174.825 169.660 174.995 ;
        RECT 169.490 174.465 169.660 174.635 ;
        RECT 169.490 174.105 169.660 174.275 ;
        RECT 169.490 173.745 169.660 173.915 ;
        RECT 169.490 173.385 169.660 173.555 ;
        RECT 169.490 173.025 169.660 173.195 ;
        RECT 169.490 172.665 169.660 172.835 ;
        RECT 169.490 149.255 169.660 149.425 ;
        RECT 169.490 148.895 169.660 149.065 ;
        RECT 169.490 148.535 169.660 148.705 ;
        RECT 169.490 148.175 169.660 148.345 ;
        RECT 169.490 147.815 169.660 147.985 ;
        RECT 169.490 147.455 169.660 147.625 ;
        RECT 169.490 147.095 169.660 147.265 ;
        RECT 169.490 146.735 169.660 146.905 ;
        RECT 169.490 146.375 169.660 146.545 ;
        RECT 169.490 146.015 169.660 146.185 ;
        RECT 169.490 145.655 169.660 145.825 ;
        RECT 169.490 145.295 169.660 145.465 ;
        RECT 169.490 144.935 169.660 145.105 ;
        RECT 169.490 144.575 169.660 144.745 ;
        RECT 169.490 144.215 169.660 144.385 ;
        RECT 169.490 143.855 169.660 144.025 ;
        RECT 169.490 143.495 169.660 143.665 ;
        RECT 169.490 120.075 169.660 120.245 ;
        RECT 169.490 119.715 169.660 119.885 ;
        RECT 169.490 119.355 169.660 119.525 ;
        RECT 169.490 118.995 169.660 119.165 ;
        RECT 169.490 118.635 169.660 118.805 ;
        RECT 169.490 118.275 169.660 118.445 ;
        RECT 169.490 117.915 169.660 118.085 ;
        RECT 169.490 117.555 169.660 117.725 ;
        RECT 169.490 117.195 169.660 117.365 ;
        RECT 169.490 116.835 169.660 117.005 ;
        RECT 169.490 116.475 169.660 116.645 ;
        RECT 169.490 116.115 169.660 116.285 ;
        RECT 169.490 115.755 169.660 115.925 ;
        RECT 169.490 115.395 169.660 115.565 ;
        RECT 169.490 115.035 169.660 115.205 ;
        RECT 169.490 114.675 169.660 114.845 ;
        RECT 169.490 114.315 169.660 114.485 ;
        RECT 169.490 90.755 169.660 90.925 ;
        RECT 169.490 90.395 169.660 90.565 ;
        RECT 169.490 90.035 169.660 90.205 ;
        RECT 169.490 89.675 169.660 89.845 ;
        RECT 169.490 89.315 169.660 89.485 ;
        RECT 169.490 88.955 169.660 89.125 ;
        RECT 169.490 88.595 169.660 88.765 ;
        RECT 169.490 88.235 169.660 88.405 ;
        RECT 169.490 87.875 169.660 88.045 ;
        RECT 169.490 87.515 169.660 87.685 ;
        RECT 169.490 87.155 169.660 87.325 ;
        RECT 169.490 86.795 169.660 86.965 ;
        RECT 169.490 86.435 169.660 86.605 ;
        RECT 169.490 86.075 169.660 86.245 ;
        RECT 169.490 85.715 169.660 85.885 ;
        RECT 169.490 85.355 169.660 85.525 ;
        RECT 169.490 84.995 169.660 85.165 ;
        RECT 169.540 61.475 169.710 61.645 ;
        RECT 169.540 61.115 169.710 61.285 ;
        RECT 169.540 60.755 169.710 60.925 ;
        RECT 169.540 60.395 169.710 60.565 ;
        RECT 169.540 60.035 169.710 60.205 ;
        RECT 169.540 59.675 169.710 59.845 ;
        RECT 169.540 59.315 169.710 59.485 ;
        RECT 169.540 58.955 169.710 59.125 ;
        RECT 169.540 58.595 169.710 58.765 ;
        RECT 169.540 58.235 169.710 58.405 ;
        RECT 169.540 57.875 169.710 58.045 ;
        RECT 169.540 57.515 169.710 57.685 ;
        RECT 169.540 57.155 169.710 57.325 ;
        RECT 169.540 56.795 169.710 56.965 ;
        RECT 169.540 56.435 169.710 56.605 ;
        RECT 169.540 56.075 169.710 56.245 ;
        RECT 169.540 55.715 169.710 55.885 ;
        RECT 169.630 31.935 169.800 32.105 ;
        RECT 169.630 31.575 169.800 31.745 ;
        RECT 169.630 31.215 169.800 31.385 ;
        RECT 169.630 30.855 169.800 31.025 ;
        RECT 169.630 30.495 169.800 30.665 ;
        RECT 169.630 30.135 169.800 30.305 ;
        RECT 169.630 29.775 169.800 29.945 ;
        RECT 169.630 29.415 169.800 29.585 ;
        RECT 169.630 29.055 169.800 29.225 ;
        RECT 169.630 28.695 169.800 28.865 ;
        RECT 169.630 28.335 169.800 28.505 ;
        RECT 169.630 27.975 169.800 28.145 ;
        RECT 201.940 207.505 202.110 207.675 ;
        RECT 201.940 207.145 202.110 207.315 ;
        RECT 201.940 206.785 202.110 206.955 ;
        RECT 201.940 206.425 202.110 206.595 ;
        RECT 201.940 206.065 202.110 206.235 ;
        RECT 201.940 205.705 202.110 205.875 ;
        RECT 201.940 205.345 202.110 205.515 ;
        RECT 201.940 204.985 202.110 205.155 ;
        RECT 201.940 204.625 202.110 204.795 ;
        RECT 201.940 204.265 202.110 204.435 ;
        RECT 201.940 203.905 202.110 204.075 ;
        RECT 201.940 203.545 202.110 203.715 ;
        RECT 201.940 203.185 202.110 203.355 ;
        RECT 201.940 202.825 202.110 202.995 ;
        RECT 201.940 202.465 202.110 202.635 ;
        RECT 201.940 202.105 202.110 202.275 ;
        RECT 201.940 201.745 202.110 201.915 ;
        RECT 204.950 209.625 205.120 209.795 ;
        RECT 204.950 209.265 205.120 209.435 ;
        RECT 204.950 208.905 205.120 209.075 ;
        RECT 204.950 208.545 205.120 208.715 ;
        RECT 210.240 209.625 210.410 209.795 ;
        RECT 210.240 209.265 210.410 209.435 ;
        RECT 210.240 208.905 210.410 209.075 ;
        RECT 210.240 208.545 210.410 208.715 ;
        RECT 204.950 204.155 205.120 204.325 ;
        RECT 204.950 203.795 205.120 203.965 ;
        RECT 204.950 203.435 205.120 203.605 ;
        RECT 204.950 203.075 205.120 203.245 ;
        RECT 210.240 204.155 210.410 204.325 ;
        RECT 210.240 203.795 210.410 203.965 ;
        RECT 210.240 203.435 210.410 203.605 ;
        RECT 210.240 203.075 210.410 203.245 ;
        RECT 204.950 198.685 205.120 198.855 ;
        RECT 204.950 198.325 205.120 198.495 ;
        RECT 204.950 197.965 205.120 198.135 ;
        RECT 204.950 197.605 205.120 197.775 ;
        RECT 210.240 198.685 210.410 198.855 ;
        RECT 210.240 198.325 210.410 198.495 ;
        RECT 210.240 197.965 210.410 198.135 ;
        RECT 210.240 197.605 210.410 197.775 ;
        RECT 204.950 193.215 205.120 193.385 ;
        RECT 210.240 193.215 210.410 193.385 ;
        RECT 215.530 214.735 215.700 214.905 ;
        RECT 215.530 214.375 215.700 214.545 ;
        RECT 215.530 214.015 215.700 214.185 ;
        RECT 215.530 209.625 215.700 209.795 ;
        RECT 215.530 209.265 215.700 209.435 ;
        RECT 215.530 208.905 215.700 209.075 ;
        RECT 215.530 208.545 215.700 208.715 ;
        RECT 215.530 204.155 215.700 204.325 ;
        RECT 215.530 203.795 215.700 203.965 ;
        RECT 215.530 203.435 215.700 203.605 ;
        RECT 215.530 203.075 215.700 203.245 ;
        RECT 215.530 198.685 215.700 198.855 ;
        RECT 215.530 198.325 215.700 198.495 ;
        RECT 215.530 197.965 215.700 198.135 ;
        RECT 215.530 197.605 215.700 197.775 ;
        RECT 215.530 193.215 215.700 193.385 ;
        RECT 231.400 215.095 231.570 215.265 ;
        RECT 220.820 214.735 220.990 214.905 ;
        RECT 220.820 214.375 220.990 214.545 ;
        RECT 220.820 214.015 220.990 214.185 ;
        RECT 220.820 209.625 220.990 209.795 ;
        RECT 220.820 209.265 220.990 209.435 ;
        RECT 220.820 208.905 220.990 209.075 ;
        RECT 220.820 208.545 220.990 208.715 ;
        RECT 220.820 204.155 220.990 204.325 ;
        RECT 220.820 203.795 220.990 203.965 ;
        RECT 220.820 203.435 220.990 203.605 ;
        RECT 220.820 203.075 220.990 203.245 ;
        RECT 220.820 198.685 220.990 198.855 ;
        RECT 220.820 198.325 220.990 198.495 ;
        RECT 220.820 197.965 220.990 198.135 ;
        RECT 220.820 197.605 220.990 197.775 ;
        RECT 220.820 193.215 220.990 193.385 ;
        RECT 226.110 214.735 226.280 214.905 ;
        RECT 226.110 214.375 226.280 214.545 ;
        RECT 226.110 214.015 226.280 214.185 ;
        RECT 231.400 214.735 231.570 214.905 ;
        RECT 231.400 214.375 231.570 214.545 ;
        RECT 231.400 214.015 231.570 214.185 ;
        RECT 237.890 215.205 238.060 215.375 ;
        RECT 237.890 214.845 238.060 215.015 ;
        RECT 243.180 215.205 243.350 215.375 ;
        RECT 248.470 215.205 248.640 215.375 ;
        RECT 253.760 215.205 253.930 215.375 ;
        RECT 259.050 215.205 259.220 215.375 ;
        RECT 237.890 214.485 238.060 214.655 ;
        RECT 237.890 214.125 238.060 214.295 ;
        RECT 243.180 214.845 243.350 215.015 ;
        RECT 243.180 214.485 243.350 214.655 ;
        RECT 243.180 214.125 243.350 214.295 ;
        RECT 226.110 209.625 226.280 209.795 ;
        RECT 226.110 209.265 226.280 209.435 ;
        RECT 226.110 208.905 226.280 209.075 ;
        RECT 226.110 208.545 226.280 208.715 ;
        RECT 226.110 204.155 226.280 204.325 ;
        RECT 226.110 203.795 226.280 203.965 ;
        RECT 226.110 203.435 226.280 203.605 ;
        RECT 226.110 203.075 226.280 203.245 ;
        RECT 226.110 198.685 226.280 198.855 ;
        RECT 226.110 198.325 226.280 198.495 ;
        RECT 226.110 197.965 226.280 198.135 ;
        RECT 226.110 197.605 226.280 197.775 ;
        RECT 204.950 192.855 205.120 193.025 ;
        RECT 204.950 192.495 205.120 192.665 ;
        RECT 210.240 192.855 210.410 193.025 ;
        RECT 204.950 192.135 205.120 192.305 ;
        RECT 210.240 192.495 210.410 192.665 ;
        RECT 215.530 192.855 215.700 193.025 ;
        RECT 210.240 192.135 210.410 192.305 ;
        RECT 215.530 192.495 215.700 192.665 ;
        RECT 226.110 193.215 226.280 193.385 ;
        RECT 231.400 209.625 231.570 209.795 ;
        RECT 231.400 209.265 231.570 209.435 ;
        RECT 231.400 208.905 231.570 209.075 ;
        RECT 231.400 208.545 231.570 208.715 ;
        RECT 231.400 204.155 231.570 204.325 ;
        RECT 231.400 203.795 231.570 203.965 ;
        RECT 231.400 203.435 231.570 203.605 ;
        RECT 231.400 203.075 231.570 203.245 ;
        RECT 231.400 198.685 231.570 198.855 ;
        RECT 231.400 198.325 231.570 198.495 ;
        RECT 231.400 197.965 231.570 198.135 ;
        RECT 231.400 197.605 231.570 197.775 ;
        RECT 220.820 192.855 220.990 193.025 ;
        RECT 220.820 192.495 220.990 192.665 ;
        RECT 231.400 193.215 231.570 193.385 ;
        RECT 234.880 207.615 235.050 207.785 ;
        RECT 234.880 207.255 235.050 207.425 ;
        RECT 234.880 206.895 235.050 207.065 ;
        RECT 234.880 206.535 235.050 206.705 ;
        RECT 234.880 206.175 235.050 206.345 ;
        RECT 234.880 205.815 235.050 205.985 ;
        RECT 234.880 205.455 235.050 205.625 ;
        RECT 234.880 205.095 235.050 205.265 ;
        RECT 234.880 204.735 235.050 204.905 ;
        RECT 234.880 204.375 235.050 204.545 ;
        RECT 234.880 204.015 235.050 204.185 ;
        RECT 234.880 203.655 235.050 203.825 ;
        RECT 234.880 203.295 235.050 203.465 ;
        RECT 234.880 202.935 235.050 203.105 ;
        RECT 234.880 202.575 235.050 202.745 ;
        RECT 234.880 202.215 235.050 202.385 ;
        RECT 234.880 201.855 235.050 202.025 ;
        RECT 226.110 192.855 226.280 193.025 ;
        RECT 226.110 192.495 226.280 192.665 ;
        RECT 231.400 192.855 231.570 193.025 ;
        RECT 215.530 192.135 215.700 192.305 ;
        RECT 220.820 192.135 220.990 192.305 ;
        RECT 226.110 192.135 226.280 192.305 ;
        RECT 231.400 192.495 231.570 192.665 ;
        RECT 231.400 192.135 231.570 192.305 ;
        RECT 201.940 178.425 202.110 178.595 ;
        RECT 201.940 178.065 202.110 178.235 ;
        RECT 201.940 177.705 202.110 177.875 ;
        RECT 201.940 177.345 202.110 177.515 ;
        RECT 201.940 176.985 202.110 177.155 ;
        RECT 201.940 176.625 202.110 176.795 ;
        RECT 201.940 176.265 202.110 176.435 ;
        RECT 201.940 175.905 202.110 176.075 ;
        RECT 201.940 175.545 202.110 175.715 ;
        RECT 201.940 175.185 202.110 175.355 ;
        RECT 201.940 174.825 202.110 174.995 ;
        RECT 201.940 174.465 202.110 174.635 ;
        RECT 201.940 174.105 202.110 174.275 ;
        RECT 201.940 173.745 202.110 173.915 ;
        RECT 201.940 173.385 202.110 173.555 ;
        RECT 201.940 173.025 202.110 173.195 ;
        RECT 201.940 172.665 202.110 172.835 ;
        RECT 204.950 186.015 205.120 186.185 ;
        RECT 204.950 185.655 205.120 185.825 ;
        RECT 210.240 186.015 210.410 186.185 ;
        RECT 215.530 186.015 215.700 186.185 ;
        RECT 220.820 186.015 220.990 186.185 ;
        RECT 226.110 186.015 226.280 186.185 ;
        RECT 204.950 185.295 205.120 185.465 ;
        RECT 204.950 184.935 205.120 185.105 ;
        RECT 210.240 185.655 210.410 185.825 ;
        RECT 210.240 185.295 210.410 185.465 ;
        RECT 210.240 184.935 210.410 185.105 ;
        RECT 204.950 180.545 205.120 180.715 ;
        RECT 204.950 180.185 205.120 180.355 ;
        RECT 204.950 179.825 205.120 179.995 ;
        RECT 204.950 179.465 205.120 179.635 ;
        RECT 210.240 180.545 210.410 180.715 ;
        RECT 210.240 180.185 210.410 180.355 ;
        RECT 210.240 179.825 210.410 179.995 ;
        RECT 210.240 179.465 210.410 179.635 ;
        RECT 204.950 175.075 205.120 175.245 ;
        RECT 204.950 174.715 205.120 174.885 ;
        RECT 204.950 174.355 205.120 174.525 ;
        RECT 204.950 173.995 205.120 174.165 ;
        RECT 210.240 175.075 210.410 175.245 ;
        RECT 210.240 174.715 210.410 174.885 ;
        RECT 210.240 174.355 210.410 174.525 ;
        RECT 210.240 173.995 210.410 174.165 ;
        RECT 204.950 169.605 205.120 169.775 ;
        RECT 204.950 169.245 205.120 169.415 ;
        RECT 204.950 168.885 205.120 169.055 ;
        RECT 204.950 168.525 205.120 168.695 ;
        RECT 210.240 169.605 210.410 169.775 ;
        RECT 210.240 169.245 210.410 169.415 ;
        RECT 210.240 168.885 210.410 169.055 ;
        RECT 210.240 168.525 210.410 168.695 ;
        RECT 204.950 164.135 205.120 164.305 ;
        RECT 210.240 164.135 210.410 164.305 ;
        RECT 215.530 185.655 215.700 185.825 ;
        RECT 215.530 185.295 215.700 185.465 ;
        RECT 215.530 184.935 215.700 185.105 ;
        RECT 215.530 180.545 215.700 180.715 ;
        RECT 215.530 180.185 215.700 180.355 ;
        RECT 215.530 179.825 215.700 179.995 ;
        RECT 215.530 179.465 215.700 179.635 ;
        RECT 215.530 175.075 215.700 175.245 ;
        RECT 215.530 174.715 215.700 174.885 ;
        RECT 215.530 174.355 215.700 174.525 ;
        RECT 215.530 173.995 215.700 174.165 ;
        RECT 215.530 169.605 215.700 169.775 ;
        RECT 215.530 169.245 215.700 169.415 ;
        RECT 215.530 168.885 215.700 169.055 ;
        RECT 215.530 168.525 215.700 168.695 ;
        RECT 215.530 164.135 215.700 164.305 ;
        RECT 231.400 186.015 231.570 186.185 ;
        RECT 220.820 185.655 220.990 185.825 ;
        RECT 220.820 185.295 220.990 185.465 ;
        RECT 220.820 184.935 220.990 185.105 ;
        RECT 220.820 180.545 220.990 180.715 ;
        RECT 220.820 180.185 220.990 180.355 ;
        RECT 220.820 179.825 220.990 179.995 ;
        RECT 220.820 179.465 220.990 179.635 ;
        RECT 220.820 175.075 220.990 175.245 ;
        RECT 220.820 174.715 220.990 174.885 ;
        RECT 220.820 174.355 220.990 174.525 ;
        RECT 220.820 173.995 220.990 174.165 ;
        RECT 220.820 169.605 220.990 169.775 ;
        RECT 220.820 169.245 220.990 169.415 ;
        RECT 220.820 168.885 220.990 169.055 ;
        RECT 220.820 168.525 220.990 168.695 ;
        RECT 220.820 164.135 220.990 164.305 ;
        RECT 226.110 185.655 226.280 185.825 ;
        RECT 231.400 185.655 231.570 185.825 ;
        RECT 226.110 185.295 226.280 185.465 ;
        RECT 226.110 184.935 226.280 185.105 ;
        RECT 226.110 180.545 226.280 180.715 ;
        RECT 226.110 180.185 226.280 180.355 ;
        RECT 226.110 179.825 226.280 179.995 ;
        RECT 226.110 179.465 226.280 179.635 ;
        RECT 226.110 175.075 226.280 175.245 ;
        RECT 226.110 174.715 226.280 174.885 ;
        RECT 226.110 174.355 226.280 174.525 ;
        RECT 226.110 173.995 226.280 174.165 ;
        RECT 226.110 169.605 226.280 169.775 ;
        RECT 226.110 169.245 226.280 169.415 ;
        RECT 226.110 168.885 226.280 169.055 ;
        RECT 226.110 168.525 226.280 168.695 ;
        RECT 204.950 163.775 205.120 163.945 ;
        RECT 204.950 163.415 205.120 163.585 ;
        RECT 210.240 163.775 210.410 163.945 ;
        RECT 204.950 163.055 205.120 163.225 ;
        RECT 210.240 163.415 210.410 163.585 ;
        RECT 215.530 163.775 215.700 163.945 ;
        RECT 210.240 163.055 210.410 163.225 ;
        RECT 215.530 163.415 215.700 163.585 ;
        RECT 226.110 164.135 226.280 164.305 ;
        RECT 231.400 185.295 231.570 185.465 ;
        RECT 231.400 184.935 231.570 185.105 ;
        RECT 231.400 180.545 231.570 180.715 ;
        RECT 231.400 180.185 231.570 180.355 ;
        RECT 231.400 179.825 231.570 179.995 ;
        RECT 231.400 179.465 231.570 179.635 ;
        RECT 231.400 175.075 231.570 175.245 ;
        RECT 231.400 174.715 231.570 174.885 ;
        RECT 231.400 174.355 231.570 174.525 ;
        RECT 231.400 173.995 231.570 174.165 ;
        RECT 231.400 169.605 231.570 169.775 ;
        RECT 231.400 169.245 231.570 169.415 ;
        RECT 231.400 168.885 231.570 169.055 ;
        RECT 231.400 168.525 231.570 168.695 ;
        RECT 220.820 163.775 220.990 163.945 ;
        RECT 220.820 163.415 220.990 163.585 ;
        RECT 231.400 164.135 231.570 164.305 ;
        RECT 237.890 209.735 238.060 209.905 ;
        RECT 237.890 209.375 238.060 209.545 ;
        RECT 237.890 209.015 238.060 209.185 ;
        RECT 237.890 208.655 238.060 208.825 ;
        RECT 243.180 209.735 243.350 209.905 ;
        RECT 243.180 209.375 243.350 209.545 ;
        RECT 243.180 209.015 243.350 209.185 ;
        RECT 243.180 208.655 243.350 208.825 ;
        RECT 237.890 204.265 238.060 204.435 ;
        RECT 237.890 203.905 238.060 204.075 ;
        RECT 237.890 203.545 238.060 203.715 ;
        RECT 237.890 203.185 238.060 203.355 ;
        RECT 243.180 204.265 243.350 204.435 ;
        RECT 243.180 203.905 243.350 204.075 ;
        RECT 243.180 203.545 243.350 203.715 ;
        RECT 243.180 203.185 243.350 203.355 ;
        RECT 237.890 198.795 238.060 198.965 ;
        RECT 237.890 198.435 238.060 198.605 ;
        RECT 237.890 198.075 238.060 198.245 ;
        RECT 237.890 197.715 238.060 197.885 ;
        RECT 243.180 198.795 243.350 198.965 ;
        RECT 243.180 198.435 243.350 198.605 ;
        RECT 243.180 198.075 243.350 198.245 ;
        RECT 243.180 197.715 243.350 197.885 ;
        RECT 237.890 193.325 238.060 193.495 ;
        RECT 243.180 193.325 243.350 193.495 ;
        RECT 248.470 214.845 248.640 215.015 ;
        RECT 248.470 214.485 248.640 214.655 ;
        RECT 248.470 214.125 248.640 214.295 ;
        RECT 248.470 209.735 248.640 209.905 ;
        RECT 248.470 209.375 248.640 209.545 ;
        RECT 248.470 209.015 248.640 209.185 ;
        RECT 248.470 208.655 248.640 208.825 ;
        RECT 248.470 204.265 248.640 204.435 ;
        RECT 248.470 203.905 248.640 204.075 ;
        RECT 248.470 203.545 248.640 203.715 ;
        RECT 248.470 203.185 248.640 203.355 ;
        RECT 248.470 198.795 248.640 198.965 ;
        RECT 248.470 198.435 248.640 198.605 ;
        RECT 248.470 198.075 248.640 198.245 ;
        RECT 248.470 197.715 248.640 197.885 ;
        RECT 248.470 193.325 248.640 193.495 ;
        RECT 264.340 215.205 264.510 215.375 ;
        RECT 253.760 214.845 253.930 215.015 ;
        RECT 253.760 214.485 253.930 214.655 ;
        RECT 253.760 214.125 253.930 214.295 ;
        RECT 253.760 209.735 253.930 209.905 ;
        RECT 253.760 209.375 253.930 209.545 ;
        RECT 253.760 209.015 253.930 209.185 ;
        RECT 253.760 208.655 253.930 208.825 ;
        RECT 253.760 204.265 253.930 204.435 ;
        RECT 253.760 203.905 253.930 204.075 ;
        RECT 253.760 203.545 253.930 203.715 ;
        RECT 253.760 203.185 253.930 203.355 ;
        RECT 253.760 198.795 253.930 198.965 ;
        RECT 253.760 198.435 253.930 198.605 ;
        RECT 253.760 198.075 253.930 198.245 ;
        RECT 253.760 197.715 253.930 197.885 ;
        RECT 253.760 193.325 253.930 193.495 ;
        RECT 259.050 214.845 259.220 215.015 ;
        RECT 259.050 214.485 259.220 214.655 ;
        RECT 259.050 214.125 259.220 214.295 ;
        RECT 264.340 214.845 264.510 215.015 ;
        RECT 264.340 214.485 264.510 214.655 ;
        RECT 264.340 214.125 264.510 214.295 ;
        RECT 270.460 215.275 270.630 215.445 ;
        RECT 270.460 214.915 270.630 215.085 ;
        RECT 275.750 215.275 275.920 215.445 ;
        RECT 281.040 215.275 281.210 215.445 ;
        RECT 286.330 215.275 286.500 215.445 ;
        RECT 291.620 215.275 291.790 215.445 ;
        RECT 270.460 214.555 270.630 214.725 ;
        RECT 270.460 214.195 270.630 214.365 ;
        RECT 275.750 214.915 275.920 215.085 ;
        RECT 275.750 214.555 275.920 214.725 ;
        RECT 275.750 214.195 275.920 214.365 ;
        RECT 259.050 209.735 259.220 209.905 ;
        RECT 259.050 209.375 259.220 209.545 ;
        RECT 259.050 209.015 259.220 209.185 ;
        RECT 259.050 208.655 259.220 208.825 ;
        RECT 259.050 204.265 259.220 204.435 ;
        RECT 259.050 203.905 259.220 204.075 ;
        RECT 259.050 203.545 259.220 203.715 ;
        RECT 259.050 203.185 259.220 203.355 ;
        RECT 259.050 198.795 259.220 198.965 ;
        RECT 259.050 198.435 259.220 198.605 ;
        RECT 259.050 198.075 259.220 198.245 ;
        RECT 259.050 197.715 259.220 197.885 ;
        RECT 237.890 192.965 238.060 193.135 ;
        RECT 237.890 192.605 238.060 192.775 ;
        RECT 243.180 192.965 243.350 193.135 ;
        RECT 237.890 192.245 238.060 192.415 ;
        RECT 243.180 192.605 243.350 192.775 ;
        RECT 248.470 192.965 248.640 193.135 ;
        RECT 243.180 192.245 243.350 192.415 ;
        RECT 248.470 192.605 248.640 192.775 ;
        RECT 259.050 193.325 259.220 193.495 ;
        RECT 264.340 209.735 264.510 209.905 ;
        RECT 264.340 209.375 264.510 209.545 ;
        RECT 264.340 209.015 264.510 209.185 ;
        RECT 264.340 208.655 264.510 208.825 ;
        RECT 264.340 204.265 264.510 204.435 ;
        RECT 264.340 203.905 264.510 204.075 ;
        RECT 264.340 203.545 264.510 203.715 ;
        RECT 264.340 203.185 264.510 203.355 ;
        RECT 264.340 198.795 264.510 198.965 ;
        RECT 264.340 198.435 264.510 198.605 ;
        RECT 264.340 198.075 264.510 198.245 ;
        RECT 264.340 197.715 264.510 197.885 ;
        RECT 253.760 192.965 253.930 193.135 ;
        RECT 253.760 192.605 253.930 192.775 ;
        RECT 264.340 193.325 264.510 193.495 ;
        RECT 267.450 207.685 267.620 207.855 ;
        RECT 267.450 207.325 267.620 207.495 ;
        RECT 267.450 206.965 267.620 207.135 ;
        RECT 267.450 206.605 267.620 206.775 ;
        RECT 267.450 206.245 267.620 206.415 ;
        RECT 267.450 205.885 267.620 206.055 ;
        RECT 267.450 205.525 267.620 205.695 ;
        RECT 267.450 205.165 267.620 205.335 ;
        RECT 267.450 204.805 267.620 204.975 ;
        RECT 267.450 204.445 267.620 204.615 ;
        RECT 267.450 204.085 267.620 204.255 ;
        RECT 267.450 203.725 267.620 203.895 ;
        RECT 267.450 203.365 267.620 203.535 ;
        RECT 267.450 203.005 267.620 203.175 ;
        RECT 267.450 202.645 267.620 202.815 ;
        RECT 267.450 202.285 267.620 202.455 ;
        RECT 267.450 201.925 267.620 202.095 ;
        RECT 259.050 192.965 259.220 193.135 ;
        RECT 259.050 192.605 259.220 192.775 ;
        RECT 264.340 192.965 264.510 193.135 ;
        RECT 248.470 192.245 248.640 192.415 ;
        RECT 253.760 192.245 253.930 192.415 ;
        RECT 259.050 192.245 259.220 192.415 ;
        RECT 264.340 192.605 264.510 192.775 ;
        RECT 264.340 192.245 264.510 192.415 ;
        RECT 237.890 186.125 238.060 186.295 ;
        RECT 243.180 186.125 243.350 186.295 ;
        RECT 234.880 178.535 235.050 178.705 ;
        RECT 234.880 178.175 235.050 178.345 ;
        RECT 234.880 177.815 235.050 177.985 ;
        RECT 234.880 177.455 235.050 177.625 ;
        RECT 234.880 177.095 235.050 177.265 ;
        RECT 234.880 176.735 235.050 176.905 ;
        RECT 234.880 176.375 235.050 176.545 ;
        RECT 234.880 176.015 235.050 176.185 ;
        RECT 234.880 175.655 235.050 175.825 ;
        RECT 234.880 175.295 235.050 175.465 ;
        RECT 234.880 174.935 235.050 175.105 ;
        RECT 234.880 174.575 235.050 174.745 ;
        RECT 234.880 174.215 235.050 174.385 ;
        RECT 234.880 173.855 235.050 174.025 ;
        RECT 234.880 173.495 235.050 173.665 ;
        RECT 234.880 173.135 235.050 173.305 ;
        RECT 234.880 172.775 235.050 172.945 ;
        RECT 226.110 163.775 226.280 163.945 ;
        RECT 226.110 163.415 226.280 163.585 ;
        RECT 231.400 163.775 231.570 163.945 ;
        RECT 215.530 163.055 215.700 163.225 ;
        RECT 220.820 163.055 220.990 163.225 ;
        RECT 226.110 163.055 226.280 163.225 ;
        RECT 231.400 163.415 231.570 163.585 ;
        RECT 231.400 163.055 231.570 163.225 ;
        RECT 204.950 156.845 205.120 157.015 ;
        RECT 201.940 149.255 202.110 149.425 ;
        RECT 201.940 148.895 202.110 149.065 ;
        RECT 201.940 148.535 202.110 148.705 ;
        RECT 201.940 148.175 202.110 148.345 ;
        RECT 201.940 147.815 202.110 147.985 ;
        RECT 201.940 147.455 202.110 147.625 ;
        RECT 201.940 147.095 202.110 147.265 ;
        RECT 201.940 146.735 202.110 146.905 ;
        RECT 201.940 146.375 202.110 146.545 ;
        RECT 201.940 146.015 202.110 146.185 ;
        RECT 201.940 145.655 202.110 145.825 ;
        RECT 201.940 145.295 202.110 145.465 ;
        RECT 201.940 144.935 202.110 145.105 ;
        RECT 201.940 144.575 202.110 144.745 ;
        RECT 201.940 144.215 202.110 144.385 ;
        RECT 201.940 143.855 202.110 144.025 ;
        RECT 201.940 143.495 202.110 143.665 ;
        RECT 204.950 156.485 205.120 156.655 ;
        RECT 210.240 156.845 210.410 157.015 ;
        RECT 215.530 156.845 215.700 157.015 ;
        RECT 220.820 156.845 220.990 157.015 ;
        RECT 226.110 156.845 226.280 157.015 ;
        RECT 204.950 156.125 205.120 156.295 ;
        RECT 204.950 155.765 205.120 155.935 ;
        RECT 210.240 156.485 210.410 156.655 ;
        RECT 210.240 156.125 210.410 156.295 ;
        RECT 210.240 155.765 210.410 155.935 ;
        RECT 204.950 151.375 205.120 151.545 ;
        RECT 204.950 151.015 205.120 151.185 ;
        RECT 204.950 150.655 205.120 150.825 ;
        RECT 204.950 150.295 205.120 150.465 ;
        RECT 210.240 151.375 210.410 151.545 ;
        RECT 210.240 151.015 210.410 151.185 ;
        RECT 210.240 150.655 210.410 150.825 ;
        RECT 210.240 150.295 210.410 150.465 ;
        RECT 204.950 145.905 205.120 146.075 ;
        RECT 204.950 145.545 205.120 145.715 ;
        RECT 204.950 145.185 205.120 145.355 ;
        RECT 204.950 144.825 205.120 144.995 ;
        RECT 210.240 145.905 210.410 146.075 ;
        RECT 210.240 145.545 210.410 145.715 ;
        RECT 210.240 145.185 210.410 145.355 ;
        RECT 210.240 144.825 210.410 144.995 ;
        RECT 204.950 140.435 205.120 140.605 ;
        RECT 204.950 140.075 205.120 140.245 ;
        RECT 204.950 139.715 205.120 139.885 ;
        RECT 204.950 139.355 205.120 139.525 ;
        RECT 210.240 140.435 210.410 140.605 ;
        RECT 210.240 140.075 210.410 140.245 ;
        RECT 210.240 139.715 210.410 139.885 ;
        RECT 210.240 139.355 210.410 139.525 ;
        RECT 204.950 134.965 205.120 135.135 ;
        RECT 210.240 134.965 210.410 135.135 ;
        RECT 215.530 156.485 215.700 156.655 ;
        RECT 215.530 156.125 215.700 156.295 ;
        RECT 215.530 155.765 215.700 155.935 ;
        RECT 215.530 151.375 215.700 151.545 ;
        RECT 215.530 151.015 215.700 151.185 ;
        RECT 215.530 150.655 215.700 150.825 ;
        RECT 215.530 150.295 215.700 150.465 ;
        RECT 215.530 145.905 215.700 146.075 ;
        RECT 215.530 145.545 215.700 145.715 ;
        RECT 215.530 145.185 215.700 145.355 ;
        RECT 215.530 144.825 215.700 144.995 ;
        RECT 215.530 140.435 215.700 140.605 ;
        RECT 215.530 140.075 215.700 140.245 ;
        RECT 215.530 139.715 215.700 139.885 ;
        RECT 215.530 139.355 215.700 139.525 ;
        RECT 215.530 134.965 215.700 135.135 ;
        RECT 231.400 156.845 231.570 157.015 ;
        RECT 220.820 156.485 220.990 156.655 ;
        RECT 220.820 156.125 220.990 156.295 ;
        RECT 220.820 155.765 220.990 155.935 ;
        RECT 220.820 151.375 220.990 151.545 ;
        RECT 220.820 151.015 220.990 151.185 ;
        RECT 220.820 150.655 220.990 150.825 ;
        RECT 220.820 150.295 220.990 150.465 ;
        RECT 220.820 145.905 220.990 146.075 ;
        RECT 220.820 145.545 220.990 145.715 ;
        RECT 220.820 145.185 220.990 145.355 ;
        RECT 220.820 144.825 220.990 144.995 ;
        RECT 220.820 140.435 220.990 140.605 ;
        RECT 220.820 140.075 220.990 140.245 ;
        RECT 220.820 139.715 220.990 139.885 ;
        RECT 220.820 139.355 220.990 139.525 ;
        RECT 220.820 134.965 220.990 135.135 ;
        RECT 226.110 156.485 226.280 156.655 ;
        RECT 226.110 156.125 226.280 156.295 ;
        RECT 231.400 156.485 231.570 156.655 ;
        RECT 226.110 155.765 226.280 155.935 ;
        RECT 226.110 151.375 226.280 151.545 ;
        RECT 226.110 151.015 226.280 151.185 ;
        RECT 226.110 150.655 226.280 150.825 ;
        RECT 226.110 150.295 226.280 150.465 ;
        RECT 226.110 145.905 226.280 146.075 ;
        RECT 226.110 145.545 226.280 145.715 ;
        RECT 226.110 145.185 226.280 145.355 ;
        RECT 226.110 144.825 226.280 144.995 ;
        RECT 226.110 140.435 226.280 140.605 ;
        RECT 226.110 140.075 226.280 140.245 ;
        RECT 226.110 139.715 226.280 139.885 ;
        RECT 226.110 139.355 226.280 139.525 ;
        RECT 204.950 134.605 205.120 134.775 ;
        RECT 204.950 134.245 205.120 134.415 ;
        RECT 210.240 134.605 210.410 134.775 ;
        RECT 210.240 134.245 210.410 134.415 ;
        RECT 215.530 134.605 215.700 134.775 ;
        RECT 204.950 133.885 205.120 134.055 ;
        RECT 210.240 133.885 210.410 134.055 ;
        RECT 215.530 134.245 215.700 134.415 ;
        RECT 226.110 134.965 226.280 135.135 ;
        RECT 231.400 156.125 231.570 156.295 ;
        RECT 231.400 155.765 231.570 155.935 ;
        RECT 231.400 151.375 231.570 151.545 ;
        RECT 231.400 151.015 231.570 151.185 ;
        RECT 231.400 150.655 231.570 150.825 ;
        RECT 231.400 150.295 231.570 150.465 ;
        RECT 231.400 145.905 231.570 146.075 ;
        RECT 231.400 145.545 231.570 145.715 ;
        RECT 231.400 145.185 231.570 145.355 ;
        RECT 231.400 144.825 231.570 144.995 ;
        RECT 231.400 140.435 231.570 140.605 ;
        RECT 231.400 140.075 231.570 140.245 ;
        RECT 231.400 139.715 231.570 139.885 ;
        RECT 231.400 139.355 231.570 139.525 ;
        RECT 220.820 134.605 220.990 134.775 ;
        RECT 220.820 134.245 220.990 134.415 ;
        RECT 231.400 134.965 231.570 135.135 ;
        RECT 237.890 185.765 238.060 185.935 ;
        RECT 248.470 186.125 248.640 186.295 ;
        RECT 253.760 186.125 253.930 186.295 ;
        RECT 259.050 186.125 259.220 186.295 ;
        RECT 237.890 185.405 238.060 185.575 ;
        RECT 237.890 185.045 238.060 185.215 ;
        RECT 243.180 185.765 243.350 185.935 ;
        RECT 243.180 185.405 243.350 185.575 ;
        RECT 243.180 185.045 243.350 185.215 ;
        RECT 237.890 180.655 238.060 180.825 ;
        RECT 237.890 180.295 238.060 180.465 ;
        RECT 237.890 179.935 238.060 180.105 ;
        RECT 237.890 179.575 238.060 179.745 ;
        RECT 243.180 180.655 243.350 180.825 ;
        RECT 243.180 180.295 243.350 180.465 ;
        RECT 243.180 179.935 243.350 180.105 ;
        RECT 243.180 179.575 243.350 179.745 ;
        RECT 237.890 175.185 238.060 175.355 ;
        RECT 237.890 174.825 238.060 174.995 ;
        RECT 237.890 174.465 238.060 174.635 ;
        RECT 237.890 174.105 238.060 174.275 ;
        RECT 243.180 175.185 243.350 175.355 ;
        RECT 243.180 174.825 243.350 174.995 ;
        RECT 243.180 174.465 243.350 174.635 ;
        RECT 243.180 174.105 243.350 174.275 ;
        RECT 237.890 169.715 238.060 169.885 ;
        RECT 237.890 169.355 238.060 169.525 ;
        RECT 237.890 168.995 238.060 169.165 ;
        RECT 237.890 168.635 238.060 168.805 ;
        RECT 243.180 169.715 243.350 169.885 ;
        RECT 243.180 169.355 243.350 169.525 ;
        RECT 243.180 168.995 243.350 169.165 ;
        RECT 243.180 168.635 243.350 168.805 ;
        RECT 237.890 164.245 238.060 164.415 ;
        RECT 243.180 164.245 243.350 164.415 ;
        RECT 248.470 185.765 248.640 185.935 ;
        RECT 248.470 185.405 248.640 185.575 ;
        RECT 248.470 185.045 248.640 185.215 ;
        RECT 248.470 180.655 248.640 180.825 ;
        RECT 248.470 180.295 248.640 180.465 ;
        RECT 248.470 179.935 248.640 180.105 ;
        RECT 248.470 179.575 248.640 179.745 ;
        RECT 248.470 175.185 248.640 175.355 ;
        RECT 248.470 174.825 248.640 174.995 ;
        RECT 248.470 174.465 248.640 174.635 ;
        RECT 248.470 174.105 248.640 174.275 ;
        RECT 248.470 169.715 248.640 169.885 ;
        RECT 248.470 169.355 248.640 169.525 ;
        RECT 248.470 168.995 248.640 169.165 ;
        RECT 248.470 168.635 248.640 168.805 ;
        RECT 248.470 164.245 248.640 164.415 ;
        RECT 264.340 186.125 264.510 186.295 ;
        RECT 253.760 185.765 253.930 185.935 ;
        RECT 253.760 185.405 253.930 185.575 ;
        RECT 253.760 185.045 253.930 185.215 ;
        RECT 253.760 180.655 253.930 180.825 ;
        RECT 253.760 180.295 253.930 180.465 ;
        RECT 253.760 179.935 253.930 180.105 ;
        RECT 253.760 179.575 253.930 179.745 ;
        RECT 253.760 175.185 253.930 175.355 ;
        RECT 253.760 174.825 253.930 174.995 ;
        RECT 253.760 174.465 253.930 174.635 ;
        RECT 253.760 174.105 253.930 174.275 ;
        RECT 253.760 169.715 253.930 169.885 ;
        RECT 253.760 169.355 253.930 169.525 ;
        RECT 253.760 168.995 253.930 169.165 ;
        RECT 253.760 168.635 253.930 168.805 ;
        RECT 253.760 164.245 253.930 164.415 ;
        RECT 259.050 185.765 259.220 185.935 ;
        RECT 259.050 185.405 259.220 185.575 ;
        RECT 259.050 185.045 259.220 185.215 ;
        RECT 259.050 180.655 259.220 180.825 ;
        RECT 259.050 180.295 259.220 180.465 ;
        RECT 259.050 179.935 259.220 180.105 ;
        RECT 259.050 179.575 259.220 179.745 ;
        RECT 259.050 175.185 259.220 175.355 ;
        RECT 259.050 174.825 259.220 174.995 ;
        RECT 259.050 174.465 259.220 174.635 ;
        RECT 259.050 174.105 259.220 174.275 ;
        RECT 259.050 169.715 259.220 169.885 ;
        RECT 259.050 169.355 259.220 169.525 ;
        RECT 259.050 168.995 259.220 169.165 ;
        RECT 259.050 168.635 259.220 168.805 ;
        RECT 237.890 163.885 238.060 164.055 ;
        RECT 237.890 163.525 238.060 163.695 ;
        RECT 243.180 163.885 243.350 164.055 ;
        RECT 237.890 163.165 238.060 163.335 ;
        RECT 243.180 163.525 243.350 163.695 ;
        RECT 248.470 163.885 248.640 164.055 ;
        RECT 243.180 163.165 243.350 163.335 ;
        RECT 248.470 163.525 248.640 163.695 ;
        RECT 259.050 164.245 259.220 164.415 ;
        RECT 264.340 185.765 264.510 185.935 ;
        RECT 264.340 185.405 264.510 185.575 ;
        RECT 264.340 185.045 264.510 185.215 ;
        RECT 264.340 180.655 264.510 180.825 ;
        RECT 264.340 180.295 264.510 180.465 ;
        RECT 264.340 179.935 264.510 180.105 ;
        RECT 264.340 179.575 264.510 179.745 ;
        RECT 264.340 175.185 264.510 175.355 ;
        RECT 264.340 174.825 264.510 174.995 ;
        RECT 264.340 174.465 264.510 174.635 ;
        RECT 264.340 174.105 264.510 174.275 ;
        RECT 264.340 169.715 264.510 169.885 ;
        RECT 264.340 169.355 264.510 169.525 ;
        RECT 264.340 168.995 264.510 169.165 ;
        RECT 264.340 168.635 264.510 168.805 ;
        RECT 253.760 163.885 253.930 164.055 ;
        RECT 253.760 163.525 253.930 163.695 ;
        RECT 264.340 164.245 264.510 164.415 ;
        RECT 270.460 209.805 270.630 209.975 ;
        RECT 270.460 209.445 270.630 209.615 ;
        RECT 270.460 209.085 270.630 209.255 ;
        RECT 270.460 208.725 270.630 208.895 ;
        RECT 275.750 209.805 275.920 209.975 ;
        RECT 275.750 209.445 275.920 209.615 ;
        RECT 275.750 209.085 275.920 209.255 ;
        RECT 275.750 208.725 275.920 208.895 ;
        RECT 270.460 204.335 270.630 204.505 ;
        RECT 270.460 203.975 270.630 204.145 ;
        RECT 270.460 203.615 270.630 203.785 ;
        RECT 270.460 203.255 270.630 203.425 ;
        RECT 275.750 204.335 275.920 204.505 ;
        RECT 275.750 203.975 275.920 204.145 ;
        RECT 275.750 203.615 275.920 203.785 ;
        RECT 275.750 203.255 275.920 203.425 ;
        RECT 270.460 198.865 270.630 199.035 ;
        RECT 270.460 198.505 270.630 198.675 ;
        RECT 270.460 198.145 270.630 198.315 ;
        RECT 270.460 197.785 270.630 197.955 ;
        RECT 275.750 198.865 275.920 199.035 ;
        RECT 275.750 198.505 275.920 198.675 ;
        RECT 275.750 198.145 275.920 198.315 ;
        RECT 275.750 197.785 275.920 197.955 ;
        RECT 270.460 193.395 270.630 193.565 ;
        RECT 275.750 193.395 275.920 193.565 ;
        RECT 281.040 214.915 281.210 215.085 ;
        RECT 281.040 214.555 281.210 214.725 ;
        RECT 281.040 214.195 281.210 214.365 ;
        RECT 281.040 209.805 281.210 209.975 ;
        RECT 281.040 209.445 281.210 209.615 ;
        RECT 281.040 209.085 281.210 209.255 ;
        RECT 281.040 208.725 281.210 208.895 ;
        RECT 281.040 204.335 281.210 204.505 ;
        RECT 281.040 203.975 281.210 204.145 ;
        RECT 281.040 203.615 281.210 203.785 ;
        RECT 281.040 203.255 281.210 203.425 ;
        RECT 281.040 198.865 281.210 199.035 ;
        RECT 281.040 198.505 281.210 198.675 ;
        RECT 281.040 198.145 281.210 198.315 ;
        RECT 281.040 197.785 281.210 197.955 ;
        RECT 281.040 193.395 281.210 193.565 ;
        RECT 296.910 215.275 297.080 215.445 ;
        RECT 286.330 214.915 286.500 215.085 ;
        RECT 286.330 214.555 286.500 214.725 ;
        RECT 286.330 214.195 286.500 214.365 ;
        RECT 286.330 209.805 286.500 209.975 ;
        RECT 286.330 209.445 286.500 209.615 ;
        RECT 286.330 209.085 286.500 209.255 ;
        RECT 286.330 208.725 286.500 208.895 ;
        RECT 286.330 204.335 286.500 204.505 ;
        RECT 286.330 203.975 286.500 204.145 ;
        RECT 286.330 203.615 286.500 203.785 ;
        RECT 286.330 203.255 286.500 203.425 ;
        RECT 286.330 198.865 286.500 199.035 ;
        RECT 286.330 198.505 286.500 198.675 ;
        RECT 286.330 198.145 286.500 198.315 ;
        RECT 286.330 197.785 286.500 197.955 ;
        RECT 286.330 193.395 286.500 193.565 ;
        RECT 291.620 214.915 291.790 215.085 ;
        RECT 291.620 214.555 291.790 214.725 ;
        RECT 291.620 214.195 291.790 214.365 ;
        RECT 296.910 214.915 297.080 215.085 ;
        RECT 312.540 215.205 312.710 215.375 ;
        RECT 315.830 215.205 316.000 215.375 ;
        RECT 319.120 215.205 319.290 215.375 ;
        RECT 312.540 214.845 312.710 215.015 ;
        RECT 315.830 214.845 316.000 215.015 ;
        RECT 296.910 214.555 297.080 214.725 ;
        RECT 291.620 209.805 291.790 209.975 ;
        RECT 291.620 209.445 291.790 209.615 ;
        RECT 291.620 209.085 291.790 209.255 ;
        RECT 291.620 208.725 291.790 208.895 ;
        RECT 291.620 204.335 291.790 204.505 ;
        RECT 291.620 203.975 291.790 204.145 ;
        RECT 291.620 203.615 291.790 203.785 ;
        RECT 291.620 203.255 291.790 203.425 ;
        RECT 291.620 198.865 291.790 199.035 ;
        RECT 291.620 198.505 291.790 198.675 ;
        RECT 291.620 198.145 291.790 198.315 ;
        RECT 291.620 197.785 291.790 197.955 ;
        RECT 270.460 193.035 270.630 193.205 ;
        RECT 275.750 193.035 275.920 193.205 ;
        RECT 270.460 192.675 270.630 192.845 ;
        RECT 270.460 192.315 270.630 192.485 ;
        RECT 275.750 192.675 275.920 192.845 ;
        RECT 281.040 193.035 281.210 193.205 ;
        RECT 275.750 192.315 275.920 192.485 ;
        RECT 281.040 192.675 281.210 192.845 ;
        RECT 291.620 193.395 291.790 193.565 ;
        RECT 296.910 214.195 297.080 214.365 ;
        RECT 296.910 209.805 297.080 209.975 ;
        RECT 311.120 212.415 311.290 212.585 ;
        RECT 311.120 212.055 311.290 212.225 ;
        RECT 311.120 211.695 311.290 211.865 ;
        RECT 311.120 211.335 311.290 211.505 ;
        RECT 311.120 210.975 311.290 211.145 ;
        RECT 311.120 210.615 311.290 210.785 ;
        RECT 311.120 210.255 311.290 210.425 ;
        RECT 311.120 209.895 311.290 210.065 ;
        RECT 296.910 209.445 297.080 209.615 ;
        RECT 296.910 209.085 297.080 209.255 ;
        RECT 296.910 208.725 297.080 208.895 ;
        RECT 296.910 204.335 297.080 204.505 ;
        RECT 296.910 203.975 297.080 204.145 ;
        RECT 296.910 203.615 297.080 203.785 ;
        RECT 296.910 203.255 297.080 203.425 ;
        RECT 297.895 201.075 299.145 208.805 ;
        RECT 311.120 209.535 311.290 209.705 ;
        RECT 311.120 209.175 311.290 209.345 ;
        RECT 311.120 208.815 311.290 208.985 ;
        RECT 311.120 208.455 311.290 208.625 ;
        RECT 311.120 208.095 311.290 208.265 ;
        RECT 311.120 207.735 311.290 207.905 ;
        RECT 311.120 207.375 311.290 207.545 ;
        RECT 311.120 207.015 311.290 207.185 ;
        RECT 311.120 206.655 311.290 206.825 ;
        RECT 311.120 206.295 311.290 206.465 ;
        RECT 311.120 205.935 311.290 206.105 ;
        RECT 311.120 205.575 311.290 205.745 ;
        RECT 311.120 205.215 311.290 205.385 ;
        RECT 312.540 211.735 312.710 211.905 ;
        RECT 312.540 211.375 312.710 211.545 ;
        RECT 312.540 208.265 312.710 208.435 ;
        RECT 312.540 207.905 312.710 208.075 ;
        RECT 312.540 204.795 312.710 204.965 ;
        RECT 312.540 204.435 312.710 204.605 ;
        RECT 312.540 201.325 312.710 201.495 ;
        RECT 315.830 211.735 316.000 211.905 ;
        RECT 315.830 211.375 316.000 211.545 ;
        RECT 315.830 208.265 316.000 208.435 ;
        RECT 315.830 207.905 316.000 208.075 ;
        RECT 315.830 204.795 316.000 204.965 ;
        RECT 315.830 204.435 316.000 204.605 ;
        RECT 312.540 200.965 312.710 201.135 ;
        RECT 315.830 201.325 316.000 201.495 ;
        RECT 319.120 214.845 319.290 215.015 ;
        RECT 322.410 215.205 322.580 215.375 ;
        RECT 322.410 214.845 322.580 215.015 ;
        RECT 319.120 211.735 319.290 211.905 ;
        RECT 319.120 211.375 319.290 211.545 ;
        RECT 319.120 208.265 319.290 208.435 ;
        RECT 319.120 207.905 319.290 208.075 ;
        RECT 319.120 204.795 319.290 204.965 ;
        RECT 319.120 204.435 319.290 204.605 ;
        RECT 325.700 215.205 325.870 215.375 ;
        RECT 328.990 215.205 329.160 215.375 ;
        RECT 334.800 215.215 334.970 215.385 ;
        RECT 341.380 215.215 341.550 215.385 ;
        RECT 358.320 217.375 358.850 217.905 ;
        RECT 325.700 214.845 325.870 215.015 ;
        RECT 328.990 214.845 329.160 215.015 ;
        RECT 322.410 211.735 322.580 211.905 ;
        RECT 322.410 211.375 322.580 211.545 ;
        RECT 322.410 208.265 322.580 208.435 ;
        RECT 322.410 207.905 322.580 208.075 ;
        RECT 322.410 204.795 322.580 204.965 ;
        RECT 322.410 204.435 322.580 204.605 ;
        RECT 325.700 211.735 325.870 211.905 ;
        RECT 325.700 211.375 325.870 211.545 ;
        RECT 325.700 208.265 325.870 208.435 ;
        RECT 325.700 207.905 325.870 208.075 ;
        RECT 325.700 204.795 325.870 204.965 ;
        RECT 325.700 204.435 325.870 204.605 ;
        RECT 315.830 200.965 316.000 201.135 ;
        RECT 319.120 201.325 319.290 201.495 ;
        RECT 319.120 200.965 319.290 201.135 ;
        RECT 322.410 201.325 322.580 201.495 ;
        RECT 322.410 200.965 322.580 201.135 ;
        RECT 325.700 201.325 325.870 201.495 ;
        RECT 334.800 214.855 334.970 215.025 ;
        RECT 330.090 212.425 330.260 212.595 ;
        RECT 328.990 211.735 329.160 211.905 ;
        RECT 328.990 211.375 329.160 211.545 ;
        RECT 328.990 208.265 329.160 208.435 ;
        RECT 328.990 207.905 329.160 208.075 ;
        RECT 328.990 204.795 329.160 204.965 ;
        RECT 328.990 204.435 329.160 204.605 ;
        RECT 330.090 212.065 330.260 212.235 ;
        RECT 330.090 211.705 330.260 211.875 ;
        RECT 330.090 211.345 330.260 211.515 ;
        RECT 330.090 210.985 330.260 211.155 ;
        RECT 330.090 210.625 330.260 210.795 ;
        RECT 330.090 210.265 330.260 210.435 ;
        RECT 330.090 209.905 330.260 210.075 ;
        RECT 330.090 209.545 330.260 209.715 ;
        RECT 330.090 209.185 330.260 209.355 ;
        RECT 330.090 208.825 330.260 208.995 ;
        RECT 330.090 208.465 330.260 208.635 ;
        RECT 330.090 208.105 330.260 208.275 ;
        RECT 330.090 207.745 330.260 207.915 ;
        RECT 330.090 207.385 330.260 207.555 ;
        RECT 330.090 207.025 330.260 207.195 ;
        RECT 330.090 206.665 330.260 206.835 ;
        RECT 330.090 206.305 330.260 206.475 ;
        RECT 330.090 205.945 330.260 206.115 ;
        RECT 330.090 205.585 330.260 205.755 ;
        RECT 330.090 205.225 330.260 205.395 ;
        RECT 334.800 211.745 334.970 211.915 ;
        RECT 334.800 211.385 334.970 211.555 ;
        RECT 334.800 208.275 334.970 208.445 ;
        RECT 334.800 207.915 334.970 208.085 ;
        RECT 334.800 204.805 334.970 204.975 ;
        RECT 334.800 204.445 334.970 204.615 ;
        RECT 325.700 200.965 325.870 201.135 ;
        RECT 328.990 201.325 329.160 201.495 ;
        RECT 341.380 214.855 341.550 215.025 ;
        RECT 347.960 215.215 348.130 215.385 ;
        RECT 347.960 214.855 348.130 215.025 ;
        RECT 350.550 215.285 350.720 215.455 ;
        RECT 353.840 215.285 354.010 215.455 ;
        RECT 357.130 215.285 357.300 215.455 ;
        RECT 350.550 214.925 350.720 215.095 ;
        RECT 353.840 214.925 354.010 215.095 ;
        RECT 341.380 211.745 341.550 211.915 ;
        RECT 341.380 211.385 341.550 211.555 ;
        RECT 347.960 211.745 348.130 211.915 ;
        RECT 347.960 211.385 348.130 211.555 ;
        RECT 349.130 212.495 349.300 212.665 ;
        RECT 349.130 212.135 349.300 212.305 ;
        RECT 349.130 211.775 349.300 211.945 ;
        RECT 349.130 211.415 349.300 211.585 ;
        RECT 349.130 211.055 349.300 211.225 ;
        RECT 349.130 210.695 349.300 210.865 ;
        RECT 349.130 210.335 349.300 210.505 ;
        RECT 349.130 209.975 349.300 210.145 ;
        RECT 349.130 209.615 349.300 209.785 ;
        RECT 349.130 209.255 349.300 209.425 ;
        RECT 341.380 208.275 341.550 208.445 ;
        RECT 341.380 207.915 341.550 208.085 ;
        RECT 341.380 204.805 341.550 204.975 ;
        RECT 341.380 204.445 341.550 204.615 ;
        RECT 347.960 208.275 348.130 208.445 ;
        RECT 347.960 207.915 348.130 208.085 ;
        RECT 347.960 204.805 348.130 204.975 ;
        RECT 347.960 204.445 348.130 204.615 ;
        RECT 334.800 201.335 334.970 201.505 ;
        RECT 328.990 200.965 329.160 201.135 ;
        RECT 334.800 200.975 334.970 201.145 ;
        RECT 341.380 201.335 341.550 201.505 ;
        RECT 349.130 208.895 349.300 209.065 ;
        RECT 349.130 208.535 349.300 208.705 ;
        RECT 349.130 208.175 349.300 208.345 ;
        RECT 349.130 207.815 349.300 207.985 ;
        RECT 349.130 207.455 349.300 207.625 ;
        RECT 349.130 207.095 349.300 207.265 ;
        RECT 349.130 206.735 349.300 206.905 ;
        RECT 349.130 206.375 349.300 206.545 ;
        RECT 349.130 206.015 349.300 206.185 ;
        RECT 349.130 205.655 349.300 205.825 ;
        RECT 349.130 205.295 349.300 205.465 ;
        RECT 350.550 211.815 350.720 211.985 ;
        RECT 350.550 211.455 350.720 211.625 ;
        RECT 350.550 208.345 350.720 208.515 ;
        RECT 350.550 207.985 350.720 208.155 ;
        RECT 350.550 204.875 350.720 205.045 ;
        RECT 350.550 204.515 350.720 204.685 ;
        RECT 341.380 200.975 341.550 201.145 ;
        RECT 347.960 201.335 348.130 201.505 ;
        RECT 350.550 201.405 350.720 201.575 ;
        RECT 353.840 211.815 354.010 211.985 ;
        RECT 353.840 211.455 354.010 211.625 ;
        RECT 353.840 208.345 354.010 208.515 ;
        RECT 353.840 207.985 354.010 208.155 ;
        RECT 353.840 204.875 354.010 205.045 ;
        RECT 353.840 204.515 354.010 204.685 ;
        RECT 347.960 200.975 348.130 201.145 ;
        RECT 350.550 201.045 350.720 201.215 ;
        RECT 353.840 201.405 354.010 201.575 ;
        RECT 357.130 214.925 357.300 215.095 ;
        RECT 360.420 215.285 360.590 215.455 ;
        RECT 360.420 214.925 360.590 215.095 ;
        RECT 357.130 211.815 357.300 211.985 ;
        RECT 357.130 211.455 357.300 211.625 ;
        RECT 357.130 208.345 357.300 208.515 ;
        RECT 357.130 207.985 357.300 208.155 ;
        RECT 357.130 204.875 357.300 205.045 ;
        RECT 357.130 204.515 357.300 204.685 ;
        RECT 363.710 215.285 363.880 215.455 ;
        RECT 367.000 215.285 367.170 215.455 ;
        RECT 363.710 214.925 363.880 215.095 ;
        RECT 367.000 214.925 367.170 215.095 ;
        RECT 360.420 211.815 360.590 211.985 ;
        RECT 360.420 211.455 360.590 211.625 ;
        RECT 360.420 208.345 360.590 208.515 ;
        RECT 360.420 207.985 360.590 208.155 ;
        RECT 360.420 204.875 360.590 205.045 ;
        RECT 360.420 204.515 360.590 204.685 ;
        RECT 363.710 211.815 363.880 211.985 ;
        RECT 363.710 211.455 363.880 211.625 ;
        RECT 363.710 208.345 363.880 208.515 ;
        RECT 363.710 207.985 363.880 208.155 ;
        RECT 363.710 204.875 363.880 205.045 ;
        RECT 363.710 204.515 363.880 204.685 ;
        RECT 353.840 201.045 354.010 201.215 ;
        RECT 357.130 201.405 357.300 201.575 ;
        RECT 357.130 201.045 357.300 201.215 ;
        RECT 360.420 201.405 360.590 201.575 ;
        RECT 360.420 201.045 360.590 201.215 ;
        RECT 363.710 201.405 363.880 201.575 ;
        RECT 367.000 211.815 367.170 211.985 ;
        RECT 367.000 211.455 367.170 211.625 ;
        RECT 367.000 208.345 367.170 208.515 ;
        RECT 367.000 207.985 367.170 208.155 ;
        RECT 367.000 204.875 367.170 205.045 ;
        RECT 367.000 204.515 367.170 204.685 ;
        RECT 368.360 204.850 369.250 214.380 ;
        RECT 363.710 201.045 363.880 201.215 ;
        RECT 367.000 201.405 367.170 201.575 ;
        RECT 367.000 201.045 367.170 201.215 ;
        RECT 296.910 198.865 297.080 199.035 ;
        RECT 296.910 198.505 297.080 198.675 ;
        RECT 296.910 198.145 297.080 198.315 ;
        RECT 296.910 197.785 297.080 197.955 ;
        RECT 392.915 197.220 393.085 197.390 ;
        RECT 393.275 197.220 393.445 197.390 ;
        RECT 393.635 197.220 393.805 197.390 ;
        RECT 425.475 197.255 425.645 197.425 ;
        RECT 425.835 197.255 426.005 197.425 ;
        RECT 426.195 197.255 426.365 197.425 ;
        RECT 286.330 193.035 286.500 193.205 ;
        RECT 286.330 192.675 286.500 192.845 ;
        RECT 296.910 193.395 297.080 193.565 ;
        RECT 385.850 195.135 386.020 195.305 ;
        RECT 389.140 195.135 389.310 195.305 ;
        RECT 291.620 193.035 291.790 193.205 ;
        RECT 291.620 192.675 291.790 192.845 ;
        RECT 296.910 193.035 297.080 193.205 ;
        RECT 281.040 192.315 281.210 192.485 ;
        RECT 286.330 192.315 286.500 192.485 ;
        RECT 291.620 192.315 291.790 192.485 ;
        RECT 296.910 192.675 297.080 192.845 ;
        RECT 296.910 192.315 297.080 192.485 ;
        RECT 267.450 178.605 267.620 178.775 ;
        RECT 267.450 178.245 267.620 178.415 ;
        RECT 267.450 177.885 267.620 178.055 ;
        RECT 267.450 177.525 267.620 177.695 ;
        RECT 267.450 177.165 267.620 177.335 ;
        RECT 267.450 176.805 267.620 176.975 ;
        RECT 267.450 176.445 267.620 176.615 ;
        RECT 267.450 176.085 267.620 176.255 ;
        RECT 267.450 175.725 267.620 175.895 ;
        RECT 267.450 175.365 267.620 175.535 ;
        RECT 267.450 175.005 267.620 175.175 ;
        RECT 267.450 174.645 267.620 174.815 ;
        RECT 267.450 174.285 267.620 174.455 ;
        RECT 267.450 173.925 267.620 174.095 ;
        RECT 267.450 173.565 267.620 173.735 ;
        RECT 267.450 173.205 267.620 173.375 ;
        RECT 267.450 172.845 267.620 173.015 ;
        RECT 259.050 163.885 259.220 164.055 ;
        RECT 259.050 163.525 259.220 163.695 ;
        RECT 264.340 163.885 264.510 164.055 ;
        RECT 248.470 163.165 248.640 163.335 ;
        RECT 253.760 163.165 253.930 163.335 ;
        RECT 264.340 163.525 264.510 163.695 ;
        RECT 259.050 163.165 259.220 163.335 ;
        RECT 264.340 163.165 264.510 163.335 ;
        RECT 237.890 156.955 238.060 157.125 ;
        RECT 243.180 156.955 243.350 157.125 ;
        RECT 234.880 149.365 235.050 149.535 ;
        RECT 234.880 149.005 235.050 149.175 ;
        RECT 234.880 148.645 235.050 148.815 ;
        RECT 234.880 148.285 235.050 148.455 ;
        RECT 234.880 147.925 235.050 148.095 ;
        RECT 234.880 147.565 235.050 147.735 ;
        RECT 234.880 147.205 235.050 147.375 ;
        RECT 234.880 146.845 235.050 147.015 ;
        RECT 234.880 146.485 235.050 146.655 ;
        RECT 234.880 146.125 235.050 146.295 ;
        RECT 234.880 145.765 235.050 145.935 ;
        RECT 234.880 145.405 235.050 145.575 ;
        RECT 234.880 145.045 235.050 145.215 ;
        RECT 234.880 144.685 235.050 144.855 ;
        RECT 234.880 144.325 235.050 144.495 ;
        RECT 234.880 143.965 235.050 144.135 ;
        RECT 234.880 143.605 235.050 143.775 ;
        RECT 226.110 134.605 226.280 134.775 ;
        RECT 226.110 134.245 226.280 134.415 ;
        RECT 231.400 134.605 231.570 134.775 ;
        RECT 215.530 133.885 215.700 134.055 ;
        RECT 220.820 133.885 220.990 134.055 ;
        RECT 226.110 133.885 226.280 134.055 ;
        RECT 231.400 134.245 231.570 134.415 ;
        RECT 231.400 133.885 231.570 134.055 ;
        RECT 204.950 127.665 205.120 127.835 ;
        RECT 204.950 127.305 205.120 127.475 ;
        RECT 210.240 127.665 210.410 127.835 ;
        RECT 215.530 127.665 215.700 127.835 ;
        RECT 220.820 127.665 220.990 127.835 ;
        RECT 226.110 127.665 226.280 127.835 ;
        RECT 210.240 127.305 210.410 127.475 ;
        RECT 201.940 120.075 202.110 120.245 ;
        RECT 201.940 119.715 202.110 119.885 ;
        RECT 201.940 119.355 202.110 119.525 ;
        RECT 201.940 118.995 202.110 119.165 ;
        RECT 201.940 118.635 202.110 118.805 ;
        RECT 201.940 118.275 202.110 118.445 ;
        RECT 201.940 117.915 202.110 118.085 ;
        RECT 201.940 117.555 202.110 117.725 ;
        RECT 201.940 117.195 202.110 117.365 ;
        RECT 201.940 116.835 202.110 117.005 ;
        RECT 201.940 116.475 202.110 116.645 ;
        RECT 201.940 116.115 202.110 116.285 ;
        RECT 201.940 115.755 202.110 115.925 ;
        RECT 201.940 115.395 202.110 115.565 ;
        RECT 201.940 115.035 202.110 115.205 ;
        RECT 201.940 114.675 202.110 114.845 ;
        RECT 201.940 114.315 202.110 114.485 ;
        RECT 204.950 126.945 205.120 127.115 ;
        RECT 204.950 126.585 205.120 126.755 ;
        RECT 210.240 126.945 210.410 127.115 ;
        RECT 210.240 126.585 210.410 126.755 ;
        RECT 204.950 122.195 205.120 122.365 ;
        RECT 204.950 121.835 205.120 122.005 ;
        RECT 204.950 121.475 205.120 121.645 ;
        RECT 204.950 121.115 205.120 121.285 ;
        RECT 210.240 122.195 210.410 122.365 ;
        RECT 210.240 121.835 210.410 122.005 ;
        RECT 210.240 121.475 210.410 121.645 ;
        RECT 210.240 121.115 210.410 121.285 ;
        RECT 204.950 116.725 205.120 116.895 ;
        RECT 204.950 116.365 205.120 116.535 ;
        RECT 204.950 116.005 205.120 116.175 ;
        RECT 204.950 115.645 205.120 115.815 ;
        RECT 210.240 116.725 210.410 116.895 ;
        RECT 210.240 116.365 210.410 116.535 ;
        RECT 210.240 116.005 210.410 116.175 ;
        RECT 210.240 115.645 210.410 115.815 ;
        RECT 204.950 111.255 205.120 111.425 ;
        RECT 204.950 110.895 205.120 111.065 ;
        RECT 204.950 110.535 205.120 110.705 ;
        RECT 204.950 110.175 205.120 110.345 ;
        RECT 210.240 111.255 210.410 111.425 ;
        RECT 210.240 110.895 210.410 111.065 ;
        RECT 210.240 110.535 210.410 110.705 ;
        RECT 210.240 110.175 210.410 110.345 ;
        RECT 204.950 105.785 205.120 105.955 ;
        RECT 210.240 105.785 210.410 105.955 ;
        RECT 215.530 127.305 215.700 127.475 ;
        RECT 215.530 126.945 215.700 127.115 ;
        RECT 215.530 126.585 215.700 126.755 ;
        RECT 215.530 122.195 215.700 122.365 ;
        RECT 215.530 121.835 215.700 122.005 ;
        RECT 215.530 121.475 215.700 121.645 ;
        RECT 215.530 121.115 215.700 121.285 ;
        RECT 215.530 116.725 215.700 116.895 ;
        RECT 215.530 116.365 215.700 116.535 ;
        RECT 215.530 116.005 215.700 116.175 ;
        RECT 215.530 115.645 215.700 115.815 ;
        RECT 215.530 111.255 215.700 111.425 ;
        RECT 215.530 110.895 215.700 111.065 ;
        RECT 215.530 110.535 215.700 110.705 ;
        RECT 215.530 110.175 215.700 110.345 ;
        RECT 215.530 105.785 215.700 105.955 ;
        RECT 231.400 127.665 231.570 127.835 ;
        RECT 220.820 127.305 220.990 127.475 ;
        RECT 220.820 126.945 220.990 127.115 ;
        RECT 220.820 126.585 220.990 126.755 ;
        RECT 220.820 122.195 220.990 122.365 ;
        RECT 220.820 121.835 220.990 122.005 ;
        RECT 220.820 121.475 220.990 121.645 ;
        RECT 220.820 121.115 220.990 121.285 ;
        RECT 220.820 116.725 220.990 116.895 ;
        RECT 220.820 116.365 220.990 116.535 ;
        RECT 220.820 116.005 220.990 116.175 ;
        RECT 220.820 115.645 220.990 115.815 ;
        RECT 220.820 111.255 220.990 111.425 ;
        RECT 220.820 110.895 220.990 111.065 ;
        RECT 220.820 110.535 220.990 110.705 ;
        RECT 220.820 110.175 220.990 110.345 ;
        RECT 220.820 105.785 220.990 105.955 ;
        RECT 226.110 127.305 226.280 127.475 ;
        RECT 226.110 126.945 226.280 127.115 ;
        RECT 226.110 126.585 226.280 126.755 ;
        RECT 226.110 122.195 226.280 122.365 ;
        RECT 226.110 121.835 226.280 122.005 ;
        RECT 226.110 121.475 226.280 121.645 ;
        RECT 226.110 121.115 226.280 121.285 ;
        RECT 226.110 116.725 226.280 116.895 ;
        RECT 226.110 116.365 226.280 116.535 ;
        RECT 226.110 116.005 226.280 116.175 ;
        RECT 226.110 115.645 226.280 115.815 ;
        RECT 226.110 111.255 226.280 111.425 ;
        RECT 226.110 110.895 226.280 111.065 ;
        RECT 226.110 110.535 226.280 110.705 ;
        RECT 226.110 110.175 226.280 110.345 ;
        RECT 204.950 105.425 205.120 105.595 ;
        RECT 204.950 105.065 205.120 105.235 ;
        RECT 210.240 105.425 210.410 105.595 ;
        RECT 204.950 104.705 205.120 104.875 ;
        RECT 210.240 105.065 210.410 105.235 ;
        RECT 215.530 105.425 215.700 105.595 ;
        RECT 210.240 104.705 210.410 104.875 ;
        RECT 215.530 105.065 215.700 105.235 ;
        RECT 226.110 105.785 226.280 105.955 ;
        RECT 231.400 127.305 231.570 127.475 ;
        RECT 231.400 126.945 231.570 127.115 ;
        RECT 231.400 126.585 231.570 126.755 ;
        RECT 231.400 122.195 231.570 122.365 ;
        RECT 231.400 121.835 231.570 122.005 ;
        RECT 231.400 121.475 231.570 121.645 ;
        RECT 231.400 121.115 231.570 121.285 ;
        RECT 231.400 116.725 231.570 116.895 ;
        RECT 231.400 116.365 231.570 116.535 ;
        RECT 231.400 116.005 231.570 116.175 ;
        RECT 231.400 115.645 231.570 115.815 ;
        RECT 231.400 111.255 231.570 111.425 ;
        RECT 231.400 110.895 231.570 111.065 ;
        RECT 231.400 110.535 231.570 110.705 ;
        RECT 231.400 110.175 231.570 110.345 ;
        RECT 220.820 105.425 220.990 105.595 ;
        RECT 220.820 105.065 220.990 105.235 ;
        RECT 231.400 105.785 231.570 105.955 ;
        RECT 237.890 156.595 238.060 156.765 ;
        RECT 248.470 156.955 248.640 157.125 ;
        RECT 253.760 156.955 253.930 157.125 ;
        RECT 259.050 156.955 259.220 157.125 ;
        RECT 237.890 156.235 238.060 156.405 ;
        RECT 237.890 155.875 238.060 156.045 ;
        RECT 243.180 156.595 243.350 156.765 ;
        RECT 243.180 156.235 243.350 156.405 ;
        RECT 243.180 155.875 243.350 156.045 ;
        RECT 237.890 151.485 238.060 151.655 ;
        RECT 237.890 151.125 238.060 151.295 ;
        RECT 237.890 150.765 238.060 150.935 ;
        RECT 237.890 150.405 238.060 150.575 ;
        RECT 243.180 151.485 243.350 151.655 ;
        RECT 243.180 151.125 243.350 151.295 ;
        RECT 243.180 150.765 243.350 150.935 ;
        RECT 243.180 150.405 243.350 150.575 ;
        RECT 237.890 146.015 238.060 146.185 ;
        RECT 237.890 145.655 238.060 145.825 ;
        RECT 237.890 145.295 238.060 145.465 ;
        RECT 237.890 144.935 238.060 145.105 ;
        RECT 243.180 146.015 243.350 146.185 ;
        RECT 243.180 145.655 243.350 145.825 ;
        RECT 243.180 145.295 243.350 145.465 ;
        RECT 243.180 144.935 243.350 145.105 ;
        RECT 237.890 140.545 238.060 140.715 ;
        RECT 237.890 140.185 238.060 140.355 ;
        RECT 237.890 139.825 238.060 139.995 ;
        RECT 237.890 139.465 238.060 139.635 ;
        RECT 243.180 140.545 243.350 140.715 ;
        RECT 243.180 140.185 243.350 140.355 ;
        RECT 243.180 139.825 243.350 139.995 ;
        RECT 243.180 139.465 243.350 139.635 ;
        RECT 237.890 135.075 238.060 135.245 ;
        RECT 243.180 135.075 243.350 135.245 ;
        RECT 248.470 156.595 248.640 156.765 ;
        RECT 248.470 156.235 248.640 156.405 ;
        RECT 248.470 155.875 248.640 156.045 ;
        RECT 248.470 151.485 248.640 151.655 ;
        RECT 248.470 151.125 248.640 151.295 ;
        RECT 248.470 150.765 248.640 150.935 ;
        RECT 248.470 150.405 248.640 150.575 ;
        RECT 248.470 146.015 248.640 146.185 ;
        RECT 248.470 145.655 248.640 145.825 ;
        RECT 248.470 145.295 248.640 145.465 ;
        RECT 248.470 144.935 248.640 145.105 ;
        RECT 248.470 140.545 248.640 140.715 ;
        RECT 248.470 140.185 248.640 140.355 ;
        RECT 248.470 139.825 248.640 139.995 ;
        RECT 248.470 139.465 248.640 139.635 ;
        RECT 248.470 135.075 248.640 135.245 ;
        RECT 264.340 156.955 264.510 157.125 ;
        RECT 253.760 156.595 253.930 156.765 ;
        RECT 253.760 156.235 253.930 156.405 ;
        RECT 253.760 155.875 253.930 156.045 ;
        RECT 253.760 151.485 253.930 151.655 ;
        RECT 253.760 151.125 253.930 151.295 ;
        RECT 253.760 150.765 253.930 150.935 ;
        RECT 253.760 150.405 253.930 150.575 ;
        RECT 253.760 146.015 253.930 146.185 ;
        RECT 253.760 145.655 253.930 145.825 ;
        RECT 253.760 145.295 253.930 145.465 ;
        RECT 253.760 144.935 253.930 145.105 ;
        RECT 253.760 140.545 253.930 140.715 ;
        RECT 253.760 140.185 253.930 140.355 ;
        RECT 253.760 139.825 253.930 139.995 ;
        RECT 253.760 139.465 253.930 139.635 ;
        RECT 253.760 135.075 253.930 135.245 ;
        RECT 259.050 156.595 259.220 156.765 ;
        RECT 259.050 156.235 259.220 156.405 ;
        RECT 259.050 155.875 259.220 156.045 ;
        RECT 259.050 151.485 259.220 151.655 ;
        RECT 259.050 151.125 259.220 151.295 ;
        RECT 259.050 150.765 259.220 150.935 ;
        RECT 259.050 150.405 259.220 150.575 ;
        RECT 259.050 146.015 259.220 146.185 ;
        RECT 259.050 145.655 259.220 145.825 ;
        RECT 259.050 145.295 259.220 145.465 ;
        RECT 259.050 144.935 259.220 145.105 ;
        RECT 259.050 140.545 259.220 140.715 ;
        RECT 259.050 140.185 259.220 140.355 ;
        RECT 259.050 139.825 259.220 139.995 ;
        RECT 259.050 139.465 259.220 139.635 ;
        RECT 237.890 134.715 238.060 134.885 ;
        RECT 237.890 134.355 238.060 134.525 ;
        RECT 243.180 134.715 243.350 134.885 ;
        RECT 237.890 133.995 238.060 134.165 ;
        RECT 243.180 134.355 243.350 134.525 ;
        RECT 248.470 134.715 248.640 134.885 ;
        RECT 243.180 133.995 243.350 134.165 ;
        RECT 248.470 134.355 248.640 134.525 ;
        RECT 259.050 135.075 259.220 135.245 ;
        RECT 264.340 156.595 264.510 156.765 ;
        RECT 264.340 156.235 264.510 156.405 ;
        RECT 264.340 155.875 264.510 156.045 ;
        RECT 264.340 151.485 264.510 151.655 ;
        RECT 264.340 151.125 264.510 151.295 ;
        RECT 264.340 150.765 264.510 150.935 ;
        RECT 264.340 150.405 264.510 150.575 ;
        RECT 264.340 146.015 264.510 146.185 ;
        RECT 264.340 145.655 264.510 145.825 ;
        RECT 264.340 145.295 264.510 145.465 ;
        RECT 264.340 144.935 264.510 145.105 ;
        RECT 264.340 140.545 264.510 140.715 ;
        RECT 264.340 140.185 264.510 140.355 ;
        RECT 264.340 139.825 264.510 139.995 ;
        RECT 264.340 139.465 264.510 139.635 ;
        RECT 253.760 134.715 253.930 134.885 ;
        RECT 253.760 134.355 253.930 134.525 ;
        RECT 264.340 135.075 264.510 135.245 ;
        RECT 270.460 186.195 270.630 186.365 ;
        RECT 270.460 185.835 270.630 186.005 ;
        RECT 275.750 186.195 275.920 186.365 ;
        RECT 281.040 186.195 281.210 186.365 ;
        RECT 286.330 186.195 286.500 186.365 ;
        RECT 291.620 186.195 291.790 186.365 ;
        RECT 270.460 185.475 270.630 185.645 ;
        RECT 270.460 185.115 270.630 185.285 ;
        RECT 275.750 185.835 275.920 186.005 ;
        RECT 275.750 185.475 275.920 185.645 ;
        RECT 275.750 185.115 275.920 185.285 ;
        RECT 270.460 180.725 270.630 180.895 ;
        RECT 270.460 180.365 270.630 180.535 ;
        RECT 270.460 180.005 270.630 180.175 ;
        RECT 270.460 179.645 270.630 179.815 ;
        RECT 275.750 180.725 275.920 180.895 ;
        RECT 275.750 180.365 275.920 180.535 ;
        RECT 275.750 180.005 275.920 180.175 ;
        RECT 275.750 179.645 275.920 179.815 ;
        RECT 270.460 175.255 270.630 175.425 ;
        RECT 270.460 174.895 270.630 175.065 ;
        RECT 270.460 174.535 270.630 174.705 ;
        RECT 270.460 174.175 270.630 174.345 ;
        RECT 275.750 175.255 275.920 175.425 ;
        RECT 275.750 174.895 275.920 175.065 ;
        RECT 275.750 174.535 275.920 174.705 ;
        RECT 275.750 174.175 275.920 174.345 ;
        RECT 270.460 169.785 270.630 169.955 ;
        RECT 270.460 169.425 270.630 169.595 ;
        RECT 270.460 169.065 270.630 169.235 ;
        RECT 270.460 168.705 270.630 168.875 ;
        RECT 275.750 169.785 275.920 169.955 ;
        RECT 275.750 169.425 275.920 169.595 ;
        RECT 275.750 169.065 275.920 169.235 ;
        RECT 275.750 168.705 275.920 168.875 ;
        RECT 270.460 164.315 270.630 164.485 ;
        RECT 275.750 164.315 275.920 164.485 ;
        RECT 281.040 185.835 281.210 186.005 ;
        RECT 281.040 185.475 281.210 185.645 ;
        RECT 281.040 185.115 281.210 185.285 ;
        RECT 281.040 180.725 281.210 180.895 ;
        RECT 281.040 180.365 281.210 180.535 ;
        RECT 281.040 180.005 281.210 180.175 ;
        RECT 281.040 179.645 281.210 179.815 ;
        RECT 281.040 175.255 281.210 175.425 ;
        RECT 281.040 174.895 281.210 175.065 ;
        RECT 281.040 174.535 281.210 174.705 ;
        RECT 281.040 174.175 281.210 174.345 ;
        RECT 281.040 169.785 281.210 169.955 ;
        RECT 281.040 169.425 281.210 169.595 ;
        RECT 281.040 169.065 281.210 169.235 ;
        RECT 281.040 168.705 281.210 168.875 ;
        RECT 281.040 164.315 281.210 164.485 ;
        RECT 296.910 186.195 297.080 186.365 ;
        RECT 286.330 185.835 286.500 186.005 ;
        RECT 286.330 185.475 286.500 185.645 ;
        RECT 286.330 185.115 286.500 185.285 ;
        RECT 286.330 180.725 286.500 180.895 ;
        RECT 286.330 180.365 286.500 180.535 ;
        RECT 286.330 180.005 286.500 180.175 ;
        RECT 286.330 179.645 286.500 179.815 ;
        RECT 286.330 175.255 286.500 175.425 ;
        RECT 286.330 174.895 286.500 175.065 ;
        RECT 286.330 174.535 286.500 174.705 ;
        RECT 286.330 174.175 286.500 174.345 ;
        RECT 286.330 169.785 286.500 169.955 ;
        RECT 286.330 169.425 286.500 169.595 ;
        RECT 286.330 169.065 286.500 169.235 ;
        RECT 286.330 168.705 286.500 168.875 ;
        RECT 286.330 164.315 286.500 164.485 ;
        RECT 291.620 185.835 291.790 186.005 ;
        RECT 296.910 185.835 297.080 186.005 ;
        RECT 291.620 185.475 291.790 185.645 ;
        RECT 291.620 185.115 291.790 185.285 ;
        RECT 291.620 180.725 291.790 180.895 ;
        RECT 291.620 180.365 291.790 180.535 ;
        RECT 291.620 180.005 291.790 180.175 ;
        RECT 291.620 179.645 291.790 179.815 ;
        RECT 291.620 175.255 291.790 175.425 ;
        RECT 291.620 174.895 291.790 175.065 ;
        RECT 291.620 174.535 291.790 174.705 ;
        RECT 291.620 174.175 291.790 174.345 ;
        RECT 291.620 169.785 291.790 169.955 ;
        RECT 291.620 169.425 291.790 169.595 ;
        RECT 291.620 169.065 291.790 169.235 ;
        RECT 291.620 168.705 291.790 168.875 ;
        RECT 270.460 163.955 270.630 164.125 ;
        RECT 270.460 163.595 270.630 163.765 ;
        RECT 275.750 163.955 275.920 164.125 ;
        RECT 270.460 163.235 270.630 163.405 ;
        RECT 275.750 163.595 275.920 163.765 ;
        RECT 281.040 163.955 281.210 164.125 ;
        RECT 275.750 163.235 275.920 163.405 ;
        RECT 281.040 163.595 281.210 163.765 ;
        RECT 291.620 164.315 291.790 164.485 ;
        RECT 296.910 185.475 297.080 185.645 ;
        RECT 296.910 185.115 297.080 185.285 ;
        RECT 296.910 180.725 297.080 180.895 ;
        RECT 296.910 180.365 297.080 180.535 ;
        RECT 296.910 180.005 297.080 180.175 ;
        RECT 296.910 179.645 297.080 179.815 ;
        RECT 296.910 175.255 297.080 175.425 ;
        RECT 296.910 174.895 297.080 175.065 ;
        RECT 296.910 174.535 297.080 174.705 ;
        RECT 296.910 174.175 297.080 174.345 ;
        RECT 298.495 172.375 299.385 179.025 ;
        RECT 383.905 178.520 384.435 194.530 ;
        RECT 385.850 194.775 386.020 194.945 ;
        RECT 385.850 191.665 386.020 191.835 ;
        RECT 385.850 191.305 386.020 191.475 ;
        RECT 385.850 188.195 386.020 188.365 ;
        RECT 385.850 187.835 386.020 188.005 ;
        RECT 385.850 184.725 386.020 184.895 ;
        RECT 385.850 184.365 386.020 184.535 ;
        RECT 385.850 181.255 386.020 181.425 ;
        RECT 385.850 180.895 386.020 181.065 ;
        RECT 385.850 177.785 386.020 177.955 ;
        RECT 389.140 194.775 389.310 194.945 ;
        RECT 389.140 191.665 389.310 191.835 ;
        RECT 389.140 191.305 389.310 191.475 ;
        RECT 389.140 188.195 389.310 188.365 ;
        RECT 389.140 187.835 389.310 188.005 ;
        RECT 389.140 184.725 389.310 184.895 ;
        RECT 389.140 184.365 389.310 184.535 ;
        RECT 389.140 181.255 389.310 181.425 ;
        RECT 389.140 180.895 389.310 181.065 ;
        RECT 389.140 177.785 389.310 177.955 ;
        RECT 392.430 195.135 392.600 195.305 ;
        RECT 395.720 195.135 395.890 195.305 ;
        RECT 399.010 195.135 399.180 195.305 ;
        RECT 392.430 194.775 392.600 194.945 ;
        RECT 392.430 191.665 392.600 191.835 ;
        RECT 392.430 191.305 392.600 191.475 ;
        RECT 392.430 188.195 392.600 188.365 ;
        RECT 392.430 187.835 392.600 188.005 ;
        RECT 392.430 184.725 392.600 184.895 ;
        RECT 392.430 184.365 392.600 184.535 ;
        RECT 392.430 181.255 392.600 181.425 ;
        RECT 392.430 180.895 392.600 181.065 ;
        RECT 392.430 177.785 392.600 177.955 ;
        RECT 395.720 194.775 395.890 194.945 ;
        RECT 399.010 194.775 399.180 194.945 ;
        RECT 395.720 191.665 395.890 191.835 ;
        RECT 395.720 191.305 395.890 191.475 ;
        RECT 395.720 188.195 395.890 188.365 ;
        RECT 395.720 187.835 395.890 188.005 ;
        RECT 395.720 184.725 395.890 184.895 ;
        RECT 395.720 184.365 395.890 184.535 ;
        RECT 395.720 181.255 395.890 181.425 ;
        RECT 395.720 180.895 395.890 181.065 ;
        RECT 395.720 177.785 395.890 177.955 ;
        RECT 399.010 191.665 399.180 191.835 ;
        RECT 399.010 191.305 399.180 191.475 ;
        RECT 399.010 188.195 399.180 188.365 ;
        RECT 399.010 187.835 399.180 188.005 ;
        RECT 399.010 184.725 399.180 184.895 ;
        RECT 399.010 184.365 399.180 184.535 ;
        RECT 399.010 181.255 399.180 181.425 ;
        RECT 399.010 180.895 399.180 181.065 ;
        RECT 399.010 177.785 399.180 177.955 ;
        RECT 400.535 178.490 401.065 194.500 ;
        RECT 385.850 177.425 386.020 177.595 ;
        RECT 389.140 177.425 389.310 177.595 ;
        RECT 392.430 177.425 392.600 177.595 ;
        RECT 395.720 177.425 395.890 177.595 ;
        RECT 405.770 195.105 405.940 195.275 ;
        RECT 405.770 194.745 405.940 194.915 ;
        RECT 405.770 191.635 405.940 191.805 ;
        RECT 405.770 191.275 405.940 191.445 ;
        RECT 405.770 188.165 405.940 188.335 ;
        RECT 405.770 187.805 405.940 187.975 ;
        RECT 405.770 184.695 405.940 184.865 ;
        RECT 405.770 184.335 405.940 184.505 ;
        RECT 405.770 181.225 405.940 181.395 ;
        RECT 405.770 180.865 405.940 181.035 ;
        RECT 405.770 177.755 405.940 177.925 ;
        RECT 412.350 195.105 412.520 195.275 ;
        RECT 412.350 194.745 412.520 194.915 ;
        RECT 412.350 191.635 412.520 191.805 ;
        RECT 412.350 191.275 412.520 191.445 ;
        RECT 412.350 188.165 412.520 188.335 ;
        RECT 412.350 187.805 412.520 187.975 ;
        RECT 412.350 184.695 412.520 184.865 ;
        RECT 412.350 184.335 412.520 184.505 ;
        RECT 412.350 181.225 412.520 181.395 ;
        RECT 412.350 180.865 412.520 181.035 ;
        RECT 412.350 177.755 412.520 177.925 ;
        RECT 419.030 195.105 419.200 195.275 ;
        RECT 422.320 195.105 422.490 195.275 ;
        RECT 417.085 178.490 417.615 194.500 ;
        RECT 399.010 177.425 399.180 177.595 ;
        RECT 405.770 177.395 405.940 177.565 ;
        RECT 419.030 194.745 419.200 194.915 ;
        RECT 419.030 191.635 419.200 191.805 ;
        RECT 419.030 191.275 419.200 191.445 ;
        RECT 419.030 188.165 419.200 188.335 ;
        RECT 419.030 187.805 419.200 187.975 ;
        RECT 419.030 184.695 419.200 184.865 ;
        RECT 419.030 184.335 419.200 184.505 ;
        RECT 419.030 181.225 419.200 181.395 ;
        RECT 419.030 180.865 419.200 181.035 ;
        RECT 419.030 177.755 419.200 177.925 ;
        RECT 422.320 194.745 422.490 194.915 ;
        RECT 422.320 191.635 422.490 191.805 ;
        RECT 422.320 191.275 422.490 191.445 ;
        RECT 422.320 188.165 422.490 188.335 ;
        RECT 422.320 187.805 422.490 187.975 ;
        RECT 422.320 184.695 422.490 184.865 ;
        RECT 422.320 184.335 422.490 184.505 ;
        RECT 422.320 181.225 422.490 181.395 ;
        RECT 422.320 180.865 422.490 181.035 ;
        RECT 422.320 177.755 422.490 177.925 ;
        RECT 425.610 195.105 425.780 195.275 ;
        RECT 428.900 195.105 429.070 195.275 ;
        RECT 432.190 195.105 432.360 195.275 ;
        RECT 425.610 194.745 425.780 194.915 ;
        RECT 425.610 191.635 425.780 191.805 ;
        RECT 425.610 191.275 425.780 191.445 ;
        RECT 425.610 188.165 425.780 188.335 ;
        RECT 425.610 187.805 425.780 187.975 ;
        RECT 425.610 184.695 425.780 184.865 ;
        RECT 425.610 184.335 425.780 184.505 ;
        RECT 425.610 181.225 425.780 181.395 ;
        RECT 425.610 180.865 425.780 181.035 ;
        RECT 425.610 177.755 425.780 177.925 ;
        RECT 428.900 194.745 429.070 194.915 ;
        RECT 432.190 194.745 432.360 194.915 ;
        RECT 428.900 191.635 429.070 191.805 ;
        RECT 428.900 191.275 429.070 191.445 ;
        RECT 428.900 188.165 429.070 188.335 ;
        RECT 428.900 187.805 429.070 187.975 ;
        RECT 428.900 184.695 429.070 184.865 ;
        RECT 428.900 184.335 429.070 184.505 ;
        RECT 428.900 181.225 429.070 181.395 ;
        RECT 428.900 180.865 429.070 181.035 ;
        RECT 428.900 177.755 429.070 177.925 ;
        RECT 432.190 191.635 432.360 191.805 ;
        RECT 432.190 191.275 432.360 191.445 ;
        RECT 432.190 188.165 432.360 188.335 ;
        RECT 432.190 187.805 432.360 187.975 ;
        RECT 432.190 184.695 432.360 184.865 ;
        RECT 432.190 184.335 432.360 184.505 ;
        RECT 432.190 181.225 432.360 181.395 ;
        RECT 432.190 180.865 432.360 181.035 ;
        RECT 432.190 177.755 432.360 177.925 ;
        RECT 433.960 178.425 434.490 194.795 ;
        RECT 412.350 177.395 412.520 177.565 ;
        RECT 419.030 177.395 419.200 177.565 ;
        RECT 422.320 177.395 422.490 177.565 ;
        RECT 425.610 177.395 425.780 177.565 ;
        RECT 428.900 177.395 429.070 177.565 ;
        RECT 432.190 177.395 432.360 177.565 ;
        RECT 296.910 169.785 297.080 169.955 ;
        RECT 296.910 169.425 297.080 169.595 ;
        RECT 296.910 169.065 297.080 169.235 ;
        RECT 296.910 168.705 297.080 168.875 ;
        RECT 286.330 163.955 286.500 164.125 ;
        RECT 286.330 163.595 286.500 163.765 ;
        RECT 296.910 164.315 297.080 164.485 ;
        RECT 291.620 163.955 291.790 164.125 ;
        RECT 291.620 163.595 291.790 163.765 ;
        RECT 296.910 163.955 297.080 164.125 ;
        RECT 281.040 163.235 281.210 163.405 ;
        RECT 286.330 163.235 286.500 163.405 ;
        RECT 296.910 163.595 297.080 163.765 ;
        RECT 291.620 163.235 291.790 163.405 ;
        RECT 296.910 163.235 297.080 163.405 ;
        RECT 270.460 157.025 270.630 157.195 ;
        RECT 275.750 157.025 275.920 157.195 ;
        RECT 267.450 149.435 267.620 149.605 ;
        RECT 267.450 149.075 267.620 149.245 ;
        RECT 267.450 148.715 267.620 148.885 ;
        RECT 267.450 148.355 267.620 148.525 ;
        RECT 267.450 147.995 267.620 148.165 ;
        RECT 267.450 147.635 267.620 147.805 ;
        RECT 267.450 147.275 267.620 147.445 ;
        RECT 267.450 146.915 267.620 147.085 ;
        RECT 267.450 146.555 267.620 146.725 ;
        RECT 267.450 146.195 267.620 146.365 ;
        RECT 267.450 145.835 267.620 146.005 ;
        RECT 267.450 145.475 267.620 145.645 ;
        RECT 267.450 145.115 267.620 145.285 ;
        RECT 267.450 144.755 267.620 144.925 ;
        RECT 267.450 144.395 267.620 144.565 ;
        RECT 267.450 144.035 267.620 144.205 ;
        RECT 267.450 143.675 267.620 143.845 ;
        RECT 259.050 134.715 259.220 134.885 ;
        RECT 259.050 134.355 259.220 134.525 ;
        RECT 264.340 134.715 264.510 134.885 ;
        RECT 248.470 133.995 248.640 134.165 ;
        RECT 253.760 133.995 253.930 134.165 ;
        RECT 264.340 134.355 264.510 134.525 ;
        RECT 259.050 133.995 259.220 134.165 ;
        RECT 264.340 133.995 264.510 134.165 ;
        RECT 234.880 120.185 235.050 120.355 ;
        RECT 234.880 119.825 235.050 119.995 ;
        RECT 234.880 119.465 235.050 119.635 ;
        RECT 234.880 119.105 235.050 119.275 ;
        RECT 234.880 118.745 235.050 118.915 ;
        RECT 234.880 118.385 235.050 118.555 ;
        RECT 234.880 118.025 235.050 118.195 ;
        RECT 234.880 117.665 235.050 117.835 ;
        RECT 234.880 117.305 235.050 117.475 ;
        RECT 234.880 116.945 235.050 117.115 ;
        RECT 234.880 116.585 235.050 116.755 ;
        RECT 234.880 116.225 235.050 116.395 ;
        RECT 234.880 115.865 235.050 116.035 ;
        RECT 234.880 115.505 235.050 115.675 ;
        RECT 234.880 115.145 235.050 115.315 ;
        RECT 234.880 114.785 235.050 114.955 ;
        RECT 234.880 114.425 235.050 114.595 ;
        RECT 226.110 105.425 226.280 105.595 ;
        RECT 226.110 105.065 226.280 105.235 ;
        RECT 231.400 105.425 231.570 105.595 ;
        RECT 215.530 104.705 215.700 104.875 ;
        RECT 220.820 104.705 220.990 104.875 ;
        RECT 231.400 105.065 231.570 105.235 ;
        RECT 226.110 104.705 226.280 104.875 ;
        RECT 231.400 104.705 231.570 104.875 ;
        RECT 201.940 90.755 202.110 90.925 ;
        RECT 201.940 90.395 202.110 90.565 ;
        RECT 201.940 90.035 202.110 90.205 ;
        RECT 201.940 89.675 202.110 89.845 ;
        RECT 201.940 89.315 202.110 89.485 ;
        RECT 201.940 88.955 202.110 89.125 ;
        RECT 201.940 88.595 202.110 88.765 ;
        RECT 201.940 88.235 202.110 88.405 ;
        RECT 201.940 87.875 202.110 88.045 ;
        RECT 201.940 87.515 202.110 87.685 ;
        RECT 201.940 87.155 202.110 87.325 ;
        RECT 201.940 86.795 202.110 86.965 ;
        RECT 201.940 86.435 202.110 86.605 ;
        RECT 201.940 86.075 202.110 86.245 ;
        RECT 201.940 85.715 202.110 85.885 ;
        RECT 201.940 85.355 202.110 85.525 ;
        RECT 201.940 84.995 202.110 85.165 ;
        RECT 204.950 98.345 205.120 98.515 ;
        RECT 204.950 97.985 205.120 98.155 ;
        RECT 210.240 98.345 210.410 98.515 ;
        RECT 215.530 98.345 215.700 98.515 ;
        RECT 220.820 98.345 220.990 98.515 ;
        RECT 226.110 98.345 226.280 98.515 ;
        RECT 204.950 97.625 205.120 97.795 ;
        RECT 204.950 97.265 205.120 97.435 ;
        RECT 210.240 97.985 210.410 98.155 ;
        RECT 210.240 97.625 210.410 97.795 ;
        RECT 210.240 97.265 210.410 97.435 ;
        RECT 204.950 92.875 205.120 93.045 ;
        RECT 204.950 92.515 205.120 92.685 ;
        RECT 204.950 92.155 205.120 92.325 ;
        RECT 204.950 91.795 205.120 91.965 ;
        RECT 210.240 92.875 210.410 93.045 ;
        RECT 210.240 92.515 210.410 92.685 ;
        RECT 210.240 92.155 210.410 92.325 ;
        RECT 210.240 91.795 210.410 91.965 ;
        RECT 204.950 87.405 205.120 87.575 ;
        RECT 204.950 87.045 205.120 87.215 ;
        RECT 204.950 86.685 205.120 86.855 ;
        RECT 204.950 86.325 205.120 86.495 ;
        RECT 210.240 87.405 210.410 87.575 ;
        RECT 210.240 87.045 210.410 87.215 ;
        RECT 210.240 86.685 210.410 86.855 ;
        RECT 210.240 86.325 210.410 86.495 ;
        RECT 204.950 81.935 205.120 82.105 ;
        RECT 204.950 81.575 205.120 81.745 ;
        RECT 204.950 81.215 205.120 81.385 ;
        RECT 204.950 80.855 205.120 81.025 ;
        RECT 210.240 81.935 210.410 82.105 ;
        RECT 210.240 81.575 210.410 81.745 ;
        RECT 210.240 81.215 210.410 81.385 ;
        RECT 210.240 80.855 210.410 81.025 ;
        RECT 204.950 76.465 205.120 76.635 ;
        RECT 210.240 76.465 210.410 76.635 ;
        RECT 215.530 97.985 215.700 98.155 ;
        RECT 215.530 97.625 215.700 97.795 ;
        RECT 215.530 97.265 215.700 97.435 ;
        RECT 215.530 92.875 215.700 93.045 ;
        RECT 215.530 92.515 215.700 92.685 ;
        RECT 215.530 92.155 215.700 92.325 ;
        RECT 215.530 91.795 215.700 91.965 ;
        RECT 215.530 87.405 215.700 87.575 ;
        RECT 215.530 87.045 215.700 87.215 ;
        RECT 215.530 86.685 215.700 86.855 ;
        RECT 215.530 86.325 215.700 86.495 ;
        RECT 215.530 81.935 215.700 82.105 ;
        RECT 215.530 81.575 215.700 81.745 ;
        RECT 215.530 81.215 215.700 81.385 ;
        RECT 215.530 80.855 215.700 81.025 ;
        RECT 215.530 76.465 215.700 76.635 ;
        RECT 231.400 98.345 231.570 98.515 ;
        RECT 220.820 97.985 220.990 98.155 ;
        RECT 220.820 97.625 220.990 97.795 ;
        RECT 220.820 97.265 220.990 97.435 ;
        RECT 220.820 92.875 220.990 93.045 ;
        RECT 220.820 92.515 220.990 92.685 ;
        RECT 220.820 92.155 220.990 92.325 ;
        RECT 220.820 91.795 220.990 91.965 ;
        RECT 220.820 87.405 220.990 87.575 ;
        RECT 220.820 87.045 220.990 87.215 ;
        RECT 220.820 86.685 220.990 86.855 ;
        RECT 220.820 86.325 220.990 86.495 ;
        RECT 220.820 81.935 220.990 82.105 ;
        RECT 220.820 81.575 220.990 81.745 ;
        RECT 220.820 81.215 220.990 81.385 ;
        RECT 220.820 80.855 220.990 81.025 ;
        RECT 220.820 76.465 220.990 76.635 ;
        RECT 226.110 97.985 226.280 98.155 ;
        RECT 226.110 97.625 226.280 97.795 ;
        RECT 226.110 97.265 226.280 97.435 ;
        RECT 226.110 92.875 226.280 93.045 ;
        RECT 226.110 92.515 226.280 92.685 ;
        RECT 226.110 92.155 226.280 92.325 ;
        RECT 226.110 91.795 226.280 91.965 ;
        RECT 226.110 87.405 226.280 87.575 ;
        RECT 226.110 87.045 226.280 87.215 ;
        RECT 226.110 86.685 226.280 86.855 ;
        RECT 226.110 86.325 226.280 86.495 ;
        RECT 226.110 81.935 226.280 82.105 ;
        RECT 226.110 81.575 226.280 81.745 ;
        RECT 226.110 81.215 226.280 81.385 ;
        RECT 226.110 80.855 226.280 81.025 ;
        RECT 204.950 76.105 205.120 76.275 ;
        RECT 204.950 75.745 205.120 75.915 ;
        RECT 210.240 76.105 210.410 76.275 ;
        RECT 204.950 75.385 205.120 75.555 ;
        RECT 210.240 75.745 210.410 75.915 ;
        RECT 215.530 76.105 215.700 76.275 ;
        RECT 210.240 75.385 210.410 75.555 ;
        RECT 215.530 75.745 215.700 75.915 ;
        RECT 226.110 76.465 226.280 76.635 ;
        RECT 231.400 97.985 231.570 98.155 ;
        RECT 231.400 97.625 231.570 97.795 ;
        RECT 231.400 97.265 231.570 97.435 ;
        RECT 231.400 92.875 231.570 93.045 ;
        RECT 231.400 92.515 231.570 92.685 ;
        RECT 231.400 92.155 231.570 92.325 ;
        RECT 231.400 91.795 231.570 91.965 ;
        RECT 231.400 87.405 231.570 87.575 ;
        RECT 231.400 87.045 231.570 87.215 ;
        RECT 231.400 86.685 231.570 86.855 ;
        RECT 231.400 86.325 231.570 86.495 ;
        RECT 231.400 81.935 231.570 82.105 ;
        RECT 231.400 81.575 231.570 81.745 ;
        RECT 231.400 81.215 231.570 81.385 ;
        RECT 231.400 80.855 231.570 81.025 ;
        RECT 220.820 76.105 220.990 76.275 ;
        RECT 220.820 75.745 220.990 75.915 ;
        RECT 231.400 76.465 231.570 76.635 ;
        RECT 237.890 127.775 238.060 127.945 ;
        RECT 237.890 127.415 238.060 127.585 ;
        RECT 243.180 127.775 243.350 127.945 ;
        RECT 248.470 127.775 248.640 127.945 ;
        RECT 253.760 127.775 253.930 127.945 ;
        RECT 259.050 127.775 259.220 127.945 ;
        RECT 237.890 127.055 238.060 127.225 ;
        RECT 237.890 126.695 238.060 126.865 ;
        RECT 243.180 127.415 243.350 127.585 ;
        RECT 243.180 127.055 243.350 127.225 ;
        RECT 243.180 126.695 243.350 126.865 ;
        RECT 237.890 122.305 238.060 122.475 ;
        RECT 237.890 121.945 238.060 122.115 ;
        RECT 237.890 121.585 238.060 121.755 ;
        RECT 237.890 121.225 238.060 121.395 ;
        RECT 243.180 122.305 243.350 122.475 ;
        RECT 243.180 121.945 243.350 122.115 ;
        RECT 243.180 121.585 243.350 121.755 ;
        RECT 243.180 121.225 243.350 121.395 ;
        RECT 237.890 116.835 238.060 117.005 ;
        RECT 237.890 116.475 238.060 116.645 ;
        RECT 237.890 116.115 238.060 116.285 ;
        RECT 237.890 115.755 238.060 115.925 ;
        RECT 243.180 116.835 243.350 117.005 ;
        RECT 243.180 116.475 243.350 116.645 ;
        RECT 243.180 116.115 243.350 116.285 ;
        RECT 243.180 115.755 243.350 115.925 ;
        RECT 237.890 111.365 238.060 111.535 ;
        RECT 237.890 111.005 238.060 111.175 ;
        RECT 237.890 110.645 238.060 110.815 ;
        RECT 237.890 110.285 238.060 110.455 ;
        RECT 243.180 111.365 243.350 111.535 ;
        RECT 243.180 111.005 243.350 111.175 ;
        RECT 243.180 110.645 243.350 110.815 ;
        RECT 243.180 110.285 243.350 110.455 ;
        RECT 237.890 105.895 238.060 106.065 ;
        RECT 243.180 105.895 243.350 106.065 ;
        RECT 248.470 127.415 248.640 127.585 ;
        RECT 248.470 127.055 248.640 127.225 ;
        RECT 248.470 126.695 248.640 126.865 ;
        RECT 248.470 122.305 248.640 122.475 ;
        RECT 248.470 121.945 248.640 122.115 ;
        RECT 248.470 121.585 248.640 121.755 ;
        RECT 248.470 121.225 248.640 121.395 ;
        RECT 248.470 116.835 248.640 117.005 ;
        RECT 248.470 116.475 248.640 116.645 ;
        RECT 248.470 116.115 248.640 116.285 ;
        RECT 248.470 115.755 248.640 115.925 ;
        RECT 248.470 111.365 248.640 111.535 ;
        RECT 248.470 111.005 248.640 111.175 ;
        RECT 248.470 110.645 248.640 110.815 ;
        RECT 248.470 110.285 248.640 110.455 ;
        RECT 248.470 105.895 248.640 106.065 ;
        RECT 264.340 127.775 264.510 127.945 ;
        RECT 253.760 127.415 253.930 127.585 ;
        RECT 253.760 127.055 253.930 127.225 ;
        RECT 253.760 126.695 253.930 126.865 ;
        RECT 253.760 122.305 253.930 122.475 ;
        RECT 253.760 121.945 253.930 122.115 ;
        RECT 253.760 121.585 253.930 121.755 ;
        RECT 253.760 121.225 253.930 121.395 ;
        RECT 253.760 116.835 253.930 117.005 ;
        RECT 253.760 116.475 253.930 116.645 ;
        RECT 253.760 116.115 253.930 116.285 ;
        RECT 253.760 115.755 253.930 115.925 ;
        RECT 253.760 111.365 253.930 111.535 ;
        RECT 253.760 111.005 253.930 111.175 ;
        RECT 253.760 110.645 253.930 110.815 ;
        RECT 253.760 110.285 253.930 110.455 ;
        RECT 253.760 105.895 253.930 106.065 ;
        RECT 259.050 127.415 259.220 127.585 ;
        RECT 259.050 127.055 259.220 127.225 ;
        RECT 259.050 126.695 259.220 126.865 ;
        RECT 259.050 122.305 259.220 122.475 ;
        RECT 259.050 121.945 259.220 122.115 ;
        RECT 259.050 121.585 259.220 121.755 ;
        RECT 259.050 121.225 259.220 121.395 ;
        RECT 259.050 116.835 259.220 117.005 ;
        RECT 259.050 116.475 259.220 116.645 ;
        RECT 259.050 116.115 259.220 116.285 ;
        RECT 259.050 115.755 259.220 115.925 ;
        RECT 259.050 111.365 259.220 111.535 ;
        RECT 259.050 111.005 259.220 111.175 ;
        RECT 259.050 110.645 259.220 110.815 ;
        RECT 259.050 110.285 259.220 110.455 ;
        RECT 237.890 105.535 238.060 105.705 ;
        RECT 243.180 105.535 243.350 105.705 ;
        RECT 237.890 105.175 238.060 105.345 ;
        RECT 237.890 104.815 238.060 104.985 ;
        RECT 243.180 105.175 243.350 105.345 ;
        RECT 248.470 105.535 248.640 105.705 ;
        RECT 243.180 104.815 243.350 104.985 ;
        RECT 248.470 105.175 248.640 105.345 ;
        RECT 259.050 105.895 259.220 106.065 ;
        RECT 264.340 127.415 264.510 127.585 ;
        RECT 264.340 127.055 264.510 127.225 ;
        RECT 264.340 126.695 264.510 126.865 ;
        RECT 264.340 122.305 264.510 122.475 ;
        RECT 264.340 121.945 264.510 122.115 ;
        RECT 264.340 121.585 264.510 121.755 ;
        RECT 264.340 121.225 264.510 121.395 ;
        RECT 264.340 116.835 264.510 117.005 ;
        RECT 264.340 116.475 264.510 116.645 ;
        RECT 264.340 116.115 264.510 116.285 ;
        RECT 264.340 115.755 264.510 115.925 ;
        RECT 264.340 111.365 264.510 111.535 ;
        RECT 264.340 111.005 264.510 111.175 ;
        RECT 264.340 110.645 264.510 110.815 ;
        RECT 264.340 110.285 264.510 110.455 ;
        RECT 253.760 105.535 253.930 105.705 ;
        RECT 253.760 105.175 253.930 105.345 ;
        RECT 264.340 105.895 264.510 106.065 ;
        RECT 270.460 156.665 270.630 156.835 ;
        RECT 281.040 157.025 281.210 157.195 ;
        RECT 286.330 157.025 286.500 157.195 ;
        RECT 291.620 157.025 291.790 157.195 ;
        RECT 270.460 156.305 270.630 156.475 ;
        RECT 270.460 155.945 270.630 156.115 ;
        RECT 275.750 156.665 275.920 156.835 ;
        RECT 275.750 156.305 275.920 156.475 ;
        RECT 275.750 155.945 275.920 156.115 ;
        RECT 270.460 151.555 270.630 151.725 ;
        RECT 270.460 151.195 270.630 151.365 ;
        RECT 270.460 150.835 270.630 151.005 ;
        RECT 270.460 150.475 270.630 150.645 ;
        RECT 275.750 151.555 275.920 151.725 ;
        RECT 275.750 151.195 275.920 151.365 ;
        RECT 275.750 150.835 275.920 151.005 ;
        RECT 275.750 150.475 275.920 150.645 ;
        RECT 270.460 146.085 270.630 146.255 ;
        RECT 270.460 145.725 270.630 145.895 ;
        RECT 270.460 145.365 270.630 145.535 ;
        RECT 270.460 145.005 270.630 145.175 ;
        RECT 275.750 146.085 275.920 146.255 ;
        RECT 275.750 145.725 275.920 145.895 ;
        RECT 275.750 145.365 275.920 145.535 ;
        RECT 275.750 145.005 275.920 145.175 ;
        RECT 270.460 140.615 270.630 140.785 ;
        RECT 270.460 140.255 270.630 140.425 ;
        RECT 270.460 139.895 270.630 140.065 ;
        RECT 270.460 139.535 270.630 139.705 ;
        RECT 275.750 140.615 275.920 140.785 ;
        RECT 275.750 140.255 275.920 140.425 ;
        RECT 275.750 139.895 275.920 140.065 ;
        RECT 275.750 139.535 275.920 139.705 ;
        RECT 270.460 135.145 270.630 135.315 ;
        RECT 275.750 135.145 275.920 135.315 ;
        RECT 281.040 156.665 281.210 156.835 ;
        RECT 281.040 156.305 281.210 156.475 ;
        RECT 281.040 155.945 281.210 156.115 ;
        RECT 281.040 151.555 281.210 151.725 ;
        RECT 281.040 151.195 281.210 151.365 ;
        RECT 281.040 150.835 281.210 151.005 ;
        RECT 281.040 150.475 281.210 150.645 ;
        RECT 281.040 146.085 281.210 146.255 ;
        RECT 281.040 145.725 281.210 145.895 ;
        RECT 281.040 145.365 281.210 145.535 ;
        RECT 281.040 145.005 281.210 145.175 ;
        RECT 281.040 140.615 281.210 140.785 ;
        RECT 281.040 140.255 281.210 140.425 ;
        RECT 281.040 139.895 281.210 140.065 ;
        RECT 281.040 139.535 281.210 139.705 ;
        RECT 281.040 135.145 281.210 135.315 ;
        RECT 296.910 157.025 297.080 157.195 ;
        RECT 286.330 156.665 286.500 156.835 ;
        RECT 286.330 156.305 286.500 156.475 ;
        RECT 286.330 155.945 286.500 156.115 ;
        RECT 286.330 151.555 286.500 151.725 ;
        RECT 286.330 151.195 286.500 151.365 ;
        RECT 286.330 150.835 286.500 151.005 ;
        RECT 286.330 150.475 286.500 150.645 ;
        RECT 286.330 146.085 286.500 146.255 ;
        RECT 286.330 145.725 286.500 145.895 ;
        RECT 286.330 145.365 286.500 145.535 ;
        RECT 286.330 145.005 286.500 145.175 ;
        RECT 286.330 140.615 286.500 140.785 ;
        RECT 286.330 140.255 286.500 140.425 ;
        RECT 286.330 139.895 286.500 140.065 ;
        RECT 286.330 139.535 286.500 139.705 ;
        RECT 286.330 135.145 286.500 135.315 ;
        RECT 291.620 156.665 291.790 156.835 ;
        RECT 291.620 156.305 291.790 156.475 ;
        RECT 291.620 155.945 291.790 156.115 ;
        RECT 291.620 151.555 291.790 151.725 ;
        RECT 291.620 151.195 291.790 151.365 ;
        RECT 291.620 150.835 291.790 151.005 ;
        RECT 291.620 150.475 291.790 150.645 ;
        RECT 291.620 146.085 291.790 146.255 ;
        RECT 291.620 145.725 291.790 145.895 ;
        RECT 291.620 145.365 291.790 145.535 ;
        RECT 291.620 145.005 291.790 145.175 ;
        RECT 291.620 140.615 291.790 140.785 ;
        RECT 291.620 140.255 291.790 140.425 ;
        RECT 291.620 139.895 291.790 140.065 ;
        RECT 291.620 139.535 291.790 139.705 ;
        RECT 270.460 134.785 270.630 134.955 ;
        RECT 270.460 134.425 270.630 134.595 ;
        RECT 275.750 134.785 275.920 134.955 ;
        RECT 270.460 134.065 270.630 134.235 ;
        RECT 275.750 134.425 275.920 134.595 ;
        RECT 281.040 134.785 281.210 134.955 ;
        RECT 275.750 134.065 275.920 134.235 ;
        RECT 281.040 134.425 281.210 134.595 ;
        RECT 291.620 135.145 291.790 135.315 ;
        RECT 296.910 156.665 297.080 156.835 ;
        RECT 296.910 156.305 297.080 156.475 ;
        RECT 296.910 155.945 297.080 156.115 ;
        RECT 296.910 151.555 297.080 151.725 ;
        RECT 296.910 151.195 297.080 151.365 ;
        RECT 296.910 150.835 297.080 151.005 ;
        RECT 296.910 150.475 297.080 150.645 ;
        RECT 296.910 146.085 297.080 146.255 ;
        RECT 296.910 145.725 297.080 145.895 ;
        RECT 296.910 145.365 297.080 145.535 ;
        RECT 296.910 145.005 297.080 145.175 ;
        RECT 296.910 140.615 297.080 140.785 ;
        RECT 298.235 142.300 299.845 149.310 ;
        RECT 296.910 140.255 297.080 140.425 ;
        RECT 296.910 139.895 297.080 140.065 ;
        RECT 296.910 139.535 297.080 139.705 ;
        RECT 286.330 134.785 286.500 134.955 ;
        RECT 286.330 134.425 286.500 134.595 ;
        RECT 296.910 135.145 297.080 135.315 ;
        RECT 291.620 134.785 291.790 134.955 ;
        RECT 291.620 134.425 291.790 134.595 ;
        RECT 296.910 134.785 297.080 134.955 ;
        RECT 281.040 134.065 281.210 134.235 ;
        RECT 286.330 134.065 286.500 134.235 ;
        RECT 296.910 134.425 297.080 134.595 ;
        RECT 291.620 134.065 291.790 134.235 ;
        RECT 296.910 134.065 297.080 134.235 ;
        RECT 267.450 120.255 267.620 120.425 ;
        RECT 267.450 119.895 267.620 120.065 ;
        RECT 267.450 119.535 267.620 119.705 ;
        RECT 267.450 119.175 267.620 119.345 ;
        RECT 267.450 118.815 267.620 118.985 ;
        RECT 267.450 118.455 267.620 118.625 ;
        RECT 267.450 118.095 267.620 118.265 ;
        RECT 267.450 117.735 267.620 117.905 ;
        RECT 267.450 117.375 267.620 117.545 ;
        RECT 267.450 117.015 267.620 117.185 ;
        RECT 267.450 116.655 267.620 116.825 ;
        RECT 267.450 116.295 267.620 116.465 ;
        RECT 267.450 115.935 267.620 116.105 ;
        RECT 267.450 115.575 267.620 115.745 ;
        RECT 267.450 115.215 267.620 115.385 ;
        RECT 267.450 114.855 267.620 115.025 ;
        RECT 267.450 114.495 267.620 114.665 ;
        RECT 259.050 105.535 259.220 105.705 ;
        RECT 259.050 105.175 259.220 105.345 ;
        RECT 264.340 105.535 264.510 105.705 ;
        RECT 248.470 104.815 248.640 104.985 ;
        RECT 253.760 104.815 253.930 104.985 ;
        RECT 259.050 104.815 259.220 104.985 ;
        RECT 264.340 105.175 264.510 105.345 ;
        RECT 264.340 104.815 264.510 104.985 ;
        RECT 237.890 98.455 238.060 98.625 ;
        RECT 243.180 98.455 243.350 98.625 ;
        RECT 234.880 90.865 235.050 91.035 ;
        RECT 234.880 90.505 235.050 90.675 ;
        RECT 234.880 90.145 235.050 90.315 ;
        RECT 234.880 89.785 235.050 89.955 ;
        RECT 234.880 89.425 235.050 89.595 ;
        RECT 234.880 89.065 235.050 89.235 ;
        RECT 234.880 88.705 235.050 88.875 ;
        RECT 234.880 88.345 235.050 88.515 ;
        RECT 234.880 87.985 235.050 88.155 ;
        RECT 234.880 87.625 235.050 87.795 ;
        RECT 234.880 87.265 235.050 87.435 ;
        RECT 234.880 86.905 235.050 87.075 ;
        RECT 234.880 86.545 235.050 86.715 ;
        RECT 234.880 86.185 235.050 86.355 ;
        RECT 234.880 85.825 235.050 85.995 ;
        RECT 234.880 85.465 235.050 85.635 ;
        RECT 234.880 85.105 235.050 85.275 ;
        RECT 226.110 76.105 226.280 76.275 ;
        RECT 226.110 75.745 226.280 75.915 ;
        RECT 231.400 76.105 231.570 76.275 ;
        RECT 215.530 75.385 215.700 75.555 ;
        RECT 220.820 75.385 220.990 75.555 ;
        RECT 226.110 75.385 226.280 75.555 ;
        RECT 231.400 75.745 231.570 75.915 ;
        RECT 231.400 75.385 231.570 75.555 ;
        RECT 201.990 61.475 202.160 61.645 ;
        RECT 201.990 61.115 202.160 61.285 ;
        RECT 201.990 60.755 202.160 60.925 ;
        RECT 201.990 60.395 202.160 60.565 ;
        RECT 201.990 60.035 202.160 60.205 ;
        RECT 201.990 59.675 202.160 59.845 ;
        RECT 201.990 59.315 202.160 59.485 ;
        RECT 201.990 58.955 202.160 59.125 ;
        RECT 201.990 58.595 202.160 58.765 ;
        RECT 201.990 58.235 202.160 58.405 ;
        RECT 201.990 57.875 202.160 58.045 ;
        RECT 201.990 57.515 202.160 57.685 ;
        RECT 201.990 57.155 202.160 57.325 ;
        RECT 201.990 56.795 202.160 56.965 ;
        RECT 201.990 56.435 202.160 56.605 ;
        RECT 201.990 56.075 202.160 56.245 ;
        RECT 201.990 55.715 202.160 55.885 ;
        RECT 205.000 69.065 205.170 69.235 ;
        RECT 205.000 68.705 205.170 68.875 ;
        RECT 210.290 69.065 210.460 69.235 ;
        RECT 215.580 69.065 215.750 69.235 ;
        RECT 220.870 69.065 221.040 69.235 ;
        RECT 226.160 69.065 226.330 69.235 ;
        RECT 205.000 68.345 205.170 68.515 ;
        RECT 205.000 67.985 205.170 68.155 ;
        RECT 210.290 68.705 210.460 68.875 ;
        RECT 210.290 68.345 210.460 68.515 ;
        RECT 210.290 67.985 210.460 68.155 ;
        RECT 205.000 63.595 205.170 63.765 ;
        RECT 205.000 63.235 205.170 63.405 ;
        RECT 205.000 62.875 205.170 63.045 ;
        RECT 205.000 62.515 205.170 62.685 ;
        RECT 210.290 63.595 210.460 63.765 ;
        RECT 210.290 63.235 210.460 63.405 ;
        RECT 210.290 62.875 210.460 63.045 ;
        RECT 210.290 62.515 210.460 62.685 ;
        RECT 205.000 58.125 205.170 58.295 ;
        RECT 205.000 57.765 205.170 57.935 ;
        RECT 205.000 57.405 205.170 57.575 ;
        RECT 205.000 57.045 205.170 57.215 ;
        RECT 210.290 58.125 210.460 58.295 ;
        RECT 210.290 57.765 210.460 57.935 ;
        RECT 210.290 57.405 210.460 57.575 ;
        RECT 210.290 57.045 210.460 57.215 ;
        RECT 205.000 52.655 205.170 52.825 ;
        RECT 205.000 52.295 205.170 52.465 ;
        RECT 205.000 51.935 205.170 52.105 ;
        RECT 205.000 51.575 205.170 51.745 ;
        RECT 210.290 52.655 210.460 52.825 ;
        RECT 210.290 52.295 210.460 52.465 ;
        RECT 210.290 51.935 210.460 52.105 ;
        RECT 210.290 51.575 210.460 51.745 ;
        RECT 205.000 47.185 205.170 47.355 ;
        RECT 210.290 47.185 210.460 47.355 ;
        RECT 215.580 68.705 215.750 68.875 ;
        RECT 215.580 68.345 215.750 68.515 ;
        RECT 215.580 67.985 215.750 68.155 ;
        RECT 215.580 63.595 215.750 63.765 ;
        RECT 215.580 63.235 215.750 63.405 ;
        RECT 215.580 62.875 215.750 63.045 ;
        RECT 215.580 62.515 215.750 62.685 ;
        RECT 215.580 58.125 215.750 58.295 ;
        RECT 215.580 57.765 215.750 57.935 ;
        RECT 215.580 57.405 215.750 57.575 ;
        RECT 215.580 57.045 215.750 57.215 ;
        RECT 215.580 52.655 215.750 52.825 ;
        RECT 215.580 52.295 215.750 52.465 ;
        RECT 215.580 51.935 215.750 52.105 ;
        RECT 215.580 51.575 215.750 51.745 ;
        RECT 215.580 47.185 215.750 47.355 ;
        RECT 231.450 69.065 231.620 69.235 ;
        RECT 220.870 68.705 221.040 68.875 ;
        RECT 220.870 68.345 221.040 68.515 ;
        RECT 220.870 67.985 221.040 68.155 ;
        RECT 220.870 63.595 221.040 63.765 ;
        RECT 220.870 63.235 221.040 63.405 ;
        RECT 220.870 62.875 221.040 63.045 ;
        RECT 220.870 62.515 221.040 62.685 ;
        RECT 220.870 58.125 221.040 58.295 ;
        RECT 220.870 57.765 221.040 57.935 ;
        RECT 220.870 57.405 221.040 57.575 ;
        RECT 220.870 57.045 221.040 57.215 ;
        RECT 220.870 52.655 221.040 52.825 ;
        RECT 220.870 52.295 221.040 52.465 ;
        RECT 220.870 51.935 221.040 52.105 ;
        RECT 220.870 51.575 221.040 51.745 ;
        RECT 220.870 47.185 221.040 47.355 ;
        RECT 226.160 68.705 226.330 68.875 ;
        RECT 226.160 68.345 226.330 68.515 ;
        RECT 231.450 68.705 231.620 68.875 ;
        RECT 231.450 68.345 231.620 68.515 ;
        RECT 226.160 67.985 226.330 68.155 ;
        RECT 226.160 63.595 226.330 63.765 ;
        RECT 226.160 63.235 226.330 63.405 ;
        RECT 226.160 62.875 226.330 63.045 ;
        RECT 226.160 62.515 226.330 62.685 ;
        RECT 226.160 58.125 226.330 58.295 ;
        RECT 226.160 57.765 226.330 57.935 ;
        RECT 226.160 57.405 226.330 57.575 ;
        RECT 226.160 57.045 226.330 57.215 ;
        RECT 226.160 52.655 226.330 52.825 ;
        RECT 226.160 52.295 226.330 52.465 ;
        RECT 226.160 51.935 226.330 52.105 ;
        RECT 226.160 51.575 226.330 51.745 ;
        RECT 205.000 46.825 205.170 46.995 ;
        RECT 205.000 46.465 205.170 46.635 ;
        RECT 210.290 46.825 210.460 46.995 ;
        RECT 205.000 46.105 205.170 46.275 ;
        RECT 210.290 46.465 210.460 46.635 ;
        RECT 215.580 46.825 215.750 46.995 ;
        RECT 210.290 46.105 210.460 46.275 ;
        RECT 215.580 46.465 215.750 46.635 ;
        RECT 226.160 47.185 226.330 47.355 ;
        RECT 231.450 67.985 231.620 68.155 ;
        RECT 231.450 63.595 231.620 63.765 ;
        RECT 231.450 63.235 231.620 63.405 ;
        RECT 231.450 62.875 231.620 63.045 ;
        RECT 231.450 62.515 231.620 62.685 ;
        RECT 231.450 58.125 231.620 58.295 ;
        RECT 231.450 57.765 231.620 57.935 ;
        RECT 231.450 57.405 231.620 57.575 ;
        RECT 231.450 57.045 231.620 57.215 ;
        RECT 231.450 52.655 231.620 52.825 ;
        RECT 231.450 52.295 231.620 52.465 ;
        RECT 231.450 51.935 231.620 52.105 ;
        RECT 231.450 51.575 231.620 51.745 ;
        RECT 220.870 46.825 221.040 46.995 ;
        RECT 220.870 46.465 221.040 46.635 ;
        RECT 231.450 47.185 231.620 47.355 ;
        RECT 237.890 98.095 238.060 98.265 ;
        RECT 248.470 98.455 248.640 98.625 ;
        RECT 253.760 98.455 253.930 98.625 ;
        RECT 259.050 98.455 259.220 98.625 ;
        RECT 237.890 97.735 238.060 97.905 ;
        RECT 237.890 97.375 238.060 97.545 ;
        RECT 243.180 98.095 243.350 98.265 ;
        RECT 243.180 97.735 243.350 97.905 ;
        RECT 243.180 97.375 243.350 97.545 ;
        RECT 237.890 92.985 238.060 93.155 ;
        RECT 237.890 92.625 238.060 92.795 ;
        RECT 237.890 92.265 238.060 92.435 ;
        RECT 237.890 91.905 238.060 92.075 ;
        RECT 243.180 92.985 243.350 93.155 ;
        RECT 243.180 92.625 243.350 92.795 ;
        RECT 243.180 92.265 243.350 92.435 ;
        RECT 243.180 91.905 243.350 92.075 ;
        RECT 237.890 87.515 238.060 87.685 ;
        RECT 237.890 87.155 238.060 87.325 ;
        RECT 237.890 86.795 238.060 86.965 ;
        RECT 237.890 86.435 238.060 86.605 ;
        RECT 243.180 87.515 243.350 87.685 ;
        RECT 243.180 87.155 243.350 87.325 ;
        RECT 243.180 86.795 243.350 86.965 ;
        RECT 243.180 86.435 243.350 86.605 ;
        RECT 237.890 82.045 238.060 82.215 ;
        RECT 237.890 81.685 238.060 81.855 ;
        RECT 237.890 81.325 238.060 81.495 ;
        RECT 237.890 80.965 238.060 81.135 ;
        RECT 243.180 82.045 243.350 82.215 ;
        RECT 243.180 81.685 243.350 81.855 ;
        RECT 243.180 81.325 243.350 81.495 ;
        RECT 243.180 80.965 243.350 81.135 ;
        RECT 237.890 76.575 238.060 76.745 ;
        RECT 243.180 76.575 243.350 76.745 ;
        RECT 248.470 98.095 248.640 98.265 ;
        RECT 248.470 97.735 248.640 97.905 ;
        RECT 248.470 97.375 248.640 97.545 ;
        RECT 248.470 92.985 248.640 93.155 ;
        RECT 248.470 92.625 248.640 92.795 ;
        RECT 248.470 92.265 248.640 92.435 ;
        RECT 248.470 91.905 248.640 92.075 ;
        RECT 248.470 87.515 248.640 87.685 ;
        RECT 248.470 87.155 248.640 87.325 ;
        RECT 248.470 86.795 248.640 86.965 ;
        RECT 248.470 86.435 248.640 86.605 ;
        RECT 248.470 82.045 248.640 82.215 ;
        RECT 248.470 81.685 248.640 81.855 ;
        RECT 248.470 81.325 248.640 81.495 ;
        RECT 248.470 80.965 248.640 81.135 ;
        RECT 248.470 76.575 248.640 76.745 ;
        RECT 264.340 98.455 264.510 98.625 ;
        RECT 253.760 98.095 253.930 98.265 ;
        RECT 253.760 97.735 253.930 97.905 ;
        RECT 253.760 97.375 253.930 97.545 ;
        RECT 253.760 92.985 253.930 93.155 ;
        RECT 253.760 92.625 253.930 92.795 ;
        RECT 253.760 92.265 253.930 92.435 ;
        RECT 253.760 91.905 253.930 92.075 ;
        RECT 253.760 87.515 253.930 87.685 ;
        RECT 253.760 87.155 253.930 87.325 ;
        RECT 253.760 86.795 253.930 86.965 ;
        RECT 253.760 86.435 253.930 86.605 ;
        RECT 253.760 82.045 253.930 82.215 ;
        RECT 253.760 81.685 253.930 81.855 ;
        RECT 253.760 81.325 253.930 81.495 ;
        RECT 253.760 80.965 253.930 81.135 ;
        RECT 253.760 76.575 253.930 76.745 ;
        RECT 259.050 98.095 259.220 98.265 ;
        RECT 259.050 97.735 259.220 97.905 ;
        RECT 259.050 97.375 259.220 97.545 ;
        RECT 259.050 92.985 259.220 93.155 ;
        RECT 259.050 92.625 259.220 92.795 ;
        RECT 259.050 92.265 259.220 92.435 ;
        RECT 259.050 91.905 259.220 92.075 ;
        RECT 259.050 87.515 259.220 87.685 ;
        RECT 259.050 87.155 259.220 87.325 ;
        RECT 259.050 86.795 259.220 86.965 ;
        RECT 259.050 86.435 259.220 86.605 ;
        RECT 259.050 82.045 259.220 82.215 ;
        RECT 259.050 81.685 259.220 81.855 ;
        RECT 259.050 81.325 259.220 81.495 ;
        RECT 259.050 80.965 259.220 81.135 ;
        RECT 237.890 76.215 238.060 76.385 ;
        RECT 237.890 75.855 238.060 76.025 ;
        RECT 243.180 76.215 243.350 76.385 ;
        RECT 237.890 75.495 238.060 75.665 ;
        RECT 243.180 75.855 243.350 76.025 ;
        RECT 248.470 76.215 248.640 76.385 ;
        RECT 243.180 75.495 243.350 75.665 ;
        RECT 248.470 75.855 248.640 76.025 ;
        RECT 259.050 76.575 259.220 76.745 ;
        RECT 264.340 98.095 264.510 98.265 ;
        RECT 264.340 97.735 264.510 97.905 ;
        RECT 264.340 97.375 264.510 97.545 ;
        RECT 264.340 92.985 264.510 93.155 ;
        RECT 264.340 92.625 264.510 92.795 ;
        RECT 264.340 92.265 264.510 92.435 ;
        RECT 264.340 91.905 264.510 92.075 ;
        RECT 264.340 87.515 264.510 87.685 ;
        RECT 264.340 87.155 264.510 87.325 ;
        RECT 264.340 86.795 264.510 86.965 ;
        RECT 264.340 86.435 264.510 86.605 ;
        RECT 264.340 82.045 264.510 82.215 ;
        RECT 264.340 81.685 264.510 81.855 ;
        RECT 264.340 81.325 264.510 81.495 ;
        RECT 264.340 80.965 264.510 81.135 ;
        RECT 253.760 76.215 253.930 76.385 ;
        RECT 253.760 75.855 253.930 76.025 ;
        RECT 259.050 76.215 259.220 76.385 ;
        RECT 259.050 75.855 259.220 76.025 ;
        RECT 248.470 75.495 248.640 75.665 ;
        RECT 253.760 75.495 253.930 75.665 ;
        RECT 259.050 75.495 259.220 75.665 ;
        RECT 264.340 76.575 264.510 76.745 ;
        RECT 270.460 127.845 270.630 128.015 ;
        RECT 270.460 127.485 270.630 127.655 ;
        RECT 275.750 127.845 275.920 128.015 ;
        RECT 281.040 127.845 281.210 128.015 ;
        RECT 286.330 127.845 286.500 128.015 ;
        RECT 291.620 127.845 291.790 128.015 ;
        RECT 270.460 127.125 270.630 127.295 ;
        RECT 270.460 126.765 270.630 126.935 ;
        RECT 275.750 127.485 275.920 127.655 ;
        RECT 275.750 127.125 275.920 127.295 ;
        RECT 275.750 126.765 275.920 126.935 ;
        RECT 270.460 122.375 270.630 122.545 ;
        RECT 270.460 122.015 270.630 122.185 ;
        RECT 270.460 121.655 270.630 121.825 ;
        RECT 270.460 121.295 270.630 121.465 ;
        RECT 275.750 122.375 275.920 122.545 ;
        RECT 275.750 122.015 275.920 122.185 ;
        RECT 275.750 121.655 275.920 121.825 ;
        RECT 275.750 121.295 275.920 121.465 ;
        RECT 270.460 116.905 270.630 117.075 ;
        RECT 270.460 116.545 270.630 116.715 ;
        RECT 270.460 116.185 270.630 116.355 ;
        RECT 270.460 115.825 270.630 115.995 ;
        RECT 275.750 116.905 275.920 117.075 ;
        RECT 275.750 116.545 275.920 116.715 ;
        RECT 275.750 116.185 275.920 116.355 ;
        RECT 275.750 115.825 275.920 115.995 ;
        RECT 270.460 111.435 270.630 111.605 ;
        RECT 270.460 111.075 270.630 111.245 ;
        RECT 270.460 110.715 270.630 110.885 ;
        RECT 270.460 110.355 270.630 110.525 ;
        RECT 275.750 111.435 275.920 111.605 ;
        RECT 275.750 111.075 275.920 111.245 ;
        RECT 275.750 110.715 275.920 110.885 ;
        RECT 275.750 110.355 275.920 110.525 ;
        RECT 270.460 105.965 270.630 106.135 ;
        RECT 275.750 105.965 275.920 106.135 ;
        RECT 281.040 127.485 281.210 127.655 ;
        RECT 281.040 127.125 281.210 127.295 ;
        RECT 281.040 126.765 281.210 126.935 ;
        RECT 281.040 122.375 281.210 122.545 ;
        RECT 281.040 122.015 281.210 122.185 ;
        RECT 281.040 121.655 281.210 121.825 ;
        RECT 281.040 121.295 281.210 121.465 ;
        RECT 281.040 116.905 281.210 117.075 ;
        RECT 281.040 116.545 281.210 116.715 ;
        RECT 281.040 116.185 281.210 116.355 ;
        RECT 281.040 115.825 281.210 115.995 ;
        RECT 281.040 111.435 281.210 111.605 ;
        RECT 281.040 111.075 281.210 111.245 ;
        RECT 281.040 110.715 281.210 110.885 ;
        RECT 281.040 110.355 281.210 110.525 ;
        RECT 281.040 105.965 281.210 106.135 ;
        RECT 338.535 131.240 338.705 131.410 ;
        RECT 338.895 131.240 339.065 131.410 ;
        RECT 339.255 131.240 339.425 131.410 ;
        RECT 339.615 131.240 339.785 131.410 ;
        RECT 339.975 131.240 340.145 131.410 ;
        RECT 340.335 131.240 340.505 131.410 ;
        RECT 340.695 131.240 340.865 131.410 ;
        RECT 470.330 131.065 470.500 131.235 ;
        RECT 470.690 131.065 470.860 131.235 ;
        RECT 471.050 131.065 471.220 131.235 ;
        RECT 471.410 131.065 471.580 131.235 ;
        RECT 471.770 131.065 471.940 131.235 ;
        RECT 296.910 127.845 297.080 128.015 ;
        RECT 286.330 127.485 286.500 127.655 ;
        RECT 286.330 127.125 286.500 127.295 ;
        RECT 286.330 126.765 286.500 126.935 ;
        RECT 286.330 122.375 286.500 122.545 ;
        RECT 286.330 122.015 286.500 122.185 ;
        RECT 286.330 121.655 286.500 121.825 ;
        RECT 286.330 121.295 286.500 121.465 ;
        RECT 286.330 116.905 286.500 117.075 ;
        RECT 286.330 116.545 286.500 116.715 ;
        RECT 286.330 116.185 286.500 116.355 ;
        RECT 286.330 115.825 286.500 115.995 ;
        RECT 286.330 111.435 286.500 111.605 ;
        RECT 286.330 111.075 286.500 111.245 ;
        RECT 286.330 110.715 286.500 110.885 ;
        RECT 286.330 110.355 286.500 110.525 ;
        RECT 286.330 105.965 286.500 106.135 ;
        RECT 291.620 127.485 291.790 127.655 ;
        RECT 291.620 127.125 291.790 127.295 ;
        RECT 291.620 126.765 291.790 126.935 ;
        RECT 291.620 122.375 291.790 122.545 ;
        RECT 291.620 122.015 291.790 122.185 ;
        RECT 291.620 121.655 291.790 121.825 ;
        RECT 291.620 121.295 291.790 121.465 ;
        RECT 291.620 116.905 291.790 117.075 ;
        RECT 291.620 116.545 291.790 116.715 ;
        RECT 291.620 116.185 291.790 116.355 ;
        RECT 291.620 115.825 291.790 115.995 ;
        RECT 291.620 111.435 291.790 111.605 ;
        RECT 291.620 111.075 291.790 111.245 ;
        RECT 291.620 110.715 291.790 110.885 ;
        RECT 291.620 110.355 291.790 110.525 ;
        RECT 270.460 105.605 270.630 105.775 ;
        RECT 270.460 105.245 270.630 105.415 ;
        RECT 275.750 105.605 275.920 105.775 ;
        RECT 270.460 104.885 270.630 105.055 ;
        RECT 275.750 105.245 275.920 105.415 ;
        RECT 281.040 105.605 281.210 105.775 ;
        RECT 275.750 104.885 275.920 105.055 ;
        RECT 281.040 105.245 281.210 105.415 ;
        RECT 291.620 105.965 291.790 106.135 ;
        RECT 296.910 127.485 297.080 127.655 ;
        RECT 296.910 127.125 297.080 127.295 ;
        RECT 296.910 126.765 297.080 126.935 ;
        RECT 310.560 127.565 310.730 127.735 ;
        RECT 310.560 127.205 310.730 127.375 ;
        RECT 315.850 127.565 316.020 127.735 ;
        RECT 321.140 127.565 321.310 127.735 ;
        RECT 326.430 127.565 326.600 127.735 ;
        RECT 331.720 127.565 331.890 127.735 ;
        RECT 310.560 126.845 310.730 127.015 ;
        RECT 310.560 126.485 310.730 126.655 ;
        RECT 315.850 127.205 316.020 127.375 ;
        RECT 315.850 126.845 316.020 127.015 ;
        RECT 315.850 126.485 316.020 126.655 ;
        RECT 296.910 122.375 297.080 122.545 ;
        RECT 296.910 122.015 297.080 122.185 ;
        RECT 296.910 121.655 297.080 121.825 ;
        RECT 296.910 121.295 297.080 121.465 ;
        RECT 296.910 116.905 297.080 117.075 ;
        RECT 296.910 116.545 297.080 116.715 ;
        RECT 296.910 116.185 297.080 116.355 ;
        RECT 296.910 115.825 297.080 115.995 ;
        RECT 298.070 113.500 299.320 121.230 ;
        RECT 310.560 122.095 310.730 122.265 ;
        RECT 310.560 121.735 310.730 121.905 ;
        RECT 310.560 121.375 310.730 121.545 ;
        RECT 310.560 121.015 310.730 121.185 ;
        RECT 315.850 122.095 316.020 122.265 ;
        RECT 315.850 121.735 316.020 121.905 ;
        RECT 315.850 121.375 316.020 121.545 ;
        RECT 315.850 121.015 316.020 121.185 ;
        RECT 307.550 119.975 307.720 120.145 ;
        RECT 307.550 119.615 307.720 119.785 ;
        RECT 307.550 119.255 307.720 119.425 ;
        RECT 307.550 118.895 307.720 119.065 ;
        RECT 307.550 118.535 307.720 118.705 ;
        RECT 307.550 118.175 307.720 118.345 ;
        RECT 307.550 117.815 307.720 117.985 ;
        RECT 307.550 117.455 307.720 117.625 ;
        RECT 307.550 117.095 307.720 117.265 ;
        RECT 307.550 116.735 307.720 116.905 ;
        RECT 307.550 116.375 307.720 116.545 ;
        RECT 307.550 116.015 307.720 116.185 ;
        RECT 307.550 115.655 307.720 115.825 ;
        RECT 307.550 115.295 307.720 115.465 ;
        RECT 307.550 114.935 307.720 115.105 ;
        RECT 307.550 114.575 307.720 114.745 ;
        RECT 307.550 114.215 307.720 114.385 ;
        RECT 310.560 116.625 310.730 116.795 ;
        RECT 310.560 116.265 310.730 116.435 ;
        RECT 310.560 115.905 310.730 116.075 ;
        RECT 310.560 115.545 310.730 115.715 ;
        RECT 315.850 116.625 316.020 116.795 ;
        RECT 315.850 116.265 316.020 116.435 ;
        RECT 315.850 115.905 316.020 116.075 ;
        RECT 315.850 115.545 316.020 115.715 ;
        RECT 296.910 111.435 297.080 111.605 ;
        RECT 296.910 111.075 297.080 111.245 ;
        RECT 296.910 110.715 297.080 110.885 ;
        RECT 296.910 110.355 297.080 110.525 ;
        RECT 286.330 105.605 286.500 105.775 ;
        RECT 286.330 105.245 286.500 105.415 ;
        RECT 296.910 105.965 297.080 106.135 ;
        RECT 310.560 111.155 310.730 111.325 ;
        RECT 310.560 110.795 310.730 110.965 ;
        RECT 310.560 110.435 310.730 110.605 ;
        RECT 310.560 110.075 310.730 110.245 ;
        RECT 315.850 111.155 316.020 111.325 ;
        RECT 315.850 110.795 316.020 110.965 ;
        RECT 315.850 110.435 316.020 110.605 ;
        RECT 315.850 110.075 316.020 110.245 ;
        RECT 291.620 105.605 291.790 105.775 ;
        RECT 291.620 105.245 291.790 105.415 ;
        RECT 296.910 105.605 297.080 105.775 ;
        RECT 310.560 105.685 310.730 105.855 ;
        RECT 281.040 104.885 281.210 105.055 ;
        RECT 286.330 104.885 286.500 105.055 ;
        RECT 291.620 104.885 291.790 105.055 ;
        RECT 296.910 105.245 297.080 105.415 ;
        RECT 315.850 105.685 316.020 105.855 ;
        RECT 321.140 127.205 321.310 127.375 ;
        RECT 321.140 126.845 321.310 127.015 ;
        RECT 321.140 126.485 321.310 126.655 ;
        RECT 321.140 122.095 321.310 122.265 ;
        RECT 321.140 121.735 321.310 121.905 ;
        RECT 321.140 121.375 321.310 121.545 ;
        RECT 321.140 121.015 321.310 121.185 ;
        RECT 321.140 116.625 321.310 116.795 ;
        RECT 321.140 116.265 321.310 116.435 ;
        RECT 321.140 115.905 321.310 116.075 ;
        RECT 321.140 115.545 321.310 115.715 ;
        RECT 321.140 111.155 321.310 111.325 ;
        RECT 321.140 110.795 321.310 110.965 ;
        RECT 321.140 110.435 321.310 110.605 ;
        RECT 321.140 110.075 321.310 110.245 ;
        RECT 321.140 105.685 321.310 105.855 ;
        RECT 337.010 127.565 337.180 127.735 ;
        RECT 342.870 127.555 343.040 127.725 ;
        RECT 326.430 127.205 326.600 127.375 ;
        RECT 326.430 126.845 326.600 127.015 ;
        RECT 326.430 126.485 326.600 126.655 ;
        RECT 326.430 122.095 326.600 122.265 ;
        RECT 326.430 121.735 326.600 121.905 ;
        RECT 326.430 121.375 326.600 121.545 ;
        RECT 326.430 121.015 326.600 121.185 ;
        RECT 326.430 116.625 326.600 116.795 ;
        RECT 326.430 116.265 326.600 116.435 ;
        RECT 326.430 115.905 326.600 116.075 ;
        RECT 326.430 115.545 326.600 115.715 ;
        RECT 326.430 111.155 326.600 111.325 ;
        RECT 326.430 110.795 326.600 110.965 ;
        RECT 326.430 110.435 326.600 110.605 ;
        RECT 326.430 110.075 326.600 110.245 ;
        RECT 326.430 105.685 326.600 105.855 ;
        RECT 331.720 127.205 331.890 127.375 ;
        RECT 331.720 126.845 331.890 127.015 ;
        RECT 331.720 126.485 331.890 126.655 ;
        RECT 331.720 122.095 331.890 122.265 ;
        RECT 331.720 121.735 331.890 121.905 ;
        RECT 331.720 121.375 331.890 121.545 ;
        RECT 331.720 121.015 331.890 121.185 ;
        RECT 331.720 116.625 331.890 116.795 ;
        RECT 331.720 116.265 331.890 116.435 ;
        RECT 331.720 115.905 331.890 116.075 ;
        RECT 331.720 115.545 331.890 115.715 ;
        RECT 331.720 111.155 331.890 111.325 ;
        RECT 331.720 110.795 331.890 110.965 ;
        RECT 331.720 110.435 331.890 110.605 ;
        RECT 331.720 110.075 331.890 110.245 ;
        RECT 310.560 105.325 310.730 105.495 ;
        RECT 296.910 104.885 297.080 105.055 ;
        RECT 310.560 104.965 310.730 105.135 ;
        RECT 315.850 105.325 316.020 105.495 ;
        RECT 310.560 104.605 310.730 104.775 ;
        RECT 315.850 104.965 316.020 105.135 ;
        RECT 321.140 105.325 321.310 105.495 ;
        RECT 315.850 104.605 316.020 104.775 ;
        RECT 321.140 104.965 321.310 105.135 ;
        RECT 331.720 105.685 331.890 105.855 ;
        RECT 337.010 127.205 337.180 127.375 ;
        RECT 337.010 126.845 337.180 127.015 ;
        RECT 342.870 127.195 343.040 127.365 ;
        RECT 348.160 127.555 348.330 127.725 ;
        RECT 353.450 127.555 353.620 127.725 ;
        RECT 358.740 127.555 358.910 127.725 ;
        RECT 364.030 127.555 364.200 127.725 ;
        RECT 342.870 126.835 343.040 127.005 ;
        RECT 337.010 126.485 337.180 126.655 ;
        RECT 337.010 122.095 337.180 122.265 ;
        RECT 337.010 121.735 337.180 121.905 ;
        RECT 337.010 121.375 337.180 121.545 ;
        RECT 337.010 121.015 337.180 121.185 ;
        RECT 337.010 116.625 337.180 116.795 ;
        RECT 337.010 116.265 337.180 116.435 ;
        RECT 337.010 115.905 337.180 116.075 ;
        RECT 337.010 115.545 337.180 115.715 ;
        RECT 337.010 111.155 337.180 111.325 ;
        RECT 337.010 110.795 337.180 110.965 ;
        RECT 337.010 110.435 337.180 110.605 ;
        RECT 337.010 110.075 337.180 110.245 ;
        RECT 326.430 105.325 326.600 105.495 ;
        RECT 326.430 104.965 326.600 105.135 ;
        RECT 337.010 105.685 337.180 105.855 ;
        RECT 339.860 119.965 340.030 120.135 ;
        RECT 339.860 119.605 340.030 119.775 ;
        RECT 339.860 119.245 340.030 119.415 ;
        RECT 339.860 118.885 340.030 119.055 ;
        RECT 339.860 118.525 340.030 118.695 ;
        RECT 339.860 118.165 340.030 118.335 ;
        RECT 339.860 117.805 340.030 117.975 ;
        RECT 339.860 117.445 340.030 117.615 ;
        RECT 339.860 117.085 340.030 117.255 ;
        RECT 339.860 116.725 340.030 116.895 ;
        RECT 339.860 116.365 340.030 116.535 ;
        RECT 339.860 116.005 340.030 116.175 ;
        RECT 339.860 115.645 340.030 115.815 ;
        RECT 339.860 115.285 340.030 115.455 ;
        RECT 339.860 114.925 340.030 115.095 ;
        RECT 339.860 114.565 340.030 114.735 ;
        RECT 339.860 114.205 340.030 114.375 ;
        RECT 331.720 105.325 331.890 105.495 ;
        RECT 331.720 104.965 331.890 105.135 ;
        RECT 337.010 105.325 337.180 105.495 ;
        RECT 321.140 104.605 321.310 104.775 ;
        RECT 326.430 104.605 326.600 104.775 ;
        RECT 331.720 104.605 331.890 104.775 ;
        RECT 337.010 104.965 337.180 105.135 ;
        RECT 337.010 104.605 337.180 104.775 ;
        RECT 270.460 98.525 270.630 98.695 ;
        RECT 275.750 98.525 275.920 98.695 ;
        RECT 267.450 90.935 267.620 91.105 ;
        RECT 267.450 90.575 267.620 90.745 ;
        RECT 267.450 90.215 267.620 90.385 ;
        RECT 267.450 89.855 267.620 90.025 ;
        RECT 267.450 89.495 267.620 89.665 ;
        RECT 267.450 89.135 267.620 89.305 ;
        RECT 267.450 88.775 267.620 88.945 ;
        RECT 267.450 88.415 267.620 88.585 ;
        RECT 267.450 88.055 267.620 88.225 ;
        RECT 267.450 87.695 267.620 87.865 ;
        RECT 267.450 87.335 267.620 87.505 ;
        RECT 267.450 86.975 267.620 87.145 ;
        RECT 267.450 86.615 267.620 86.785 ;
        RECT 267.450 86.255 267.620 86.425 ;
        RECT 267.450 85.895 267.620 86.065 ;
        RECT 267.450 85.535 267.620 85.705 ;
        RECT 267.450 85.175 267.620 85.345 ;
        RECT 264.340 76.215 264.510 76.385 ;
        RECT 264.340 75.855 264.510 76.025 ;
        RECT 264.340 75.495 264.510 75.665 ;
        RECT 234.930 61.585 235.100 61.755 ;
        RECT 234.930 61.225 235.100 61.395 ;
        RECT 234.930 60.865 235.100 61.035 ;
        RECT 234.930 60.505 235.100 60.675 ;
        RECT 234.930 60.145 235.100 60.315 ;
        RECT 234.930 59.785 235.100 59.955 ;
        RECT 234.930 59.425 235.100 59.595 ;
        RECT 234.930 59.065 235.100 59.235 ;
        RECT 234.930 58.705 235.100 58.875 ;
        RECT 234.930 58.345 235.100 58.515 ;
        RECT 234.930 57.985 235.100 58.155 ;
        RECT 234.930 57.625 235.100 57.795 ;
        RECT 234.930 57.265 235.100 57.435 ;
        RECT 234.930 56.905 235.100 57.075 ;
        RECT 234.930 56.545 235.100 56.715 ;
        RECT 234.930 56.185 235.100 56.355 ;
        RECT 234.930 55.825 235.100 55.995 ;
        RECT 226.160 46.825 226.330 46.995 ;
        RECT 226.160 46.465 226.330 46.635 ;
        RECT 231.450 46.825 231.620 46.995 ;
        RECT 215.580 46.105 215.750 46.275 ;
        RECT 220.870 46.105 221.040 46.275 ;
        RECT 226.160 46.105 226.330 46.275 ;
        RECT 231.450 46.465 231.620 46.635 ;
        RECT 231.450 46.105 231.620 46.275 ;
        RECT 202.080 31.935 202.250 32.105 ;
        RECT 202.080 31.575 202.250 31.745 ;
        RECT 202.080 31.215 202.250 31.385 ;
        RECT 202.080 30.855 202.250 31.025 ;
        RECT 202.080 30.495 202.250 30.665 ;
        RECT 202.080 30.135 202.250 30.305 ;
        RECT 202.080 29.775 202.250 29.945 ;
        RECT 202.080 29.415 202.250 29.585 ;
        RECT 202.080 29.055 202.250 29.225 ;
        RECT 202.080 28.695 202.250 28.865 ;
        RECT 202.080 28.335 202.250 28.505 ;
        RECT 202.080 27.975 202.250 28.145 ;
        RECT 205.090 39.525 205.260 39.695 ;
        RECT 205.090 39.165 205.260 39.335 ;
        RECT 210.380 39.525 210.550 39.695 ;
        RECT 215.670 39.525 215.840 39.695 ;
        RECT 220.960 39.525 221.130 39.695 ;
        RECT 226.250 39.525 226.420 39.695 ;
        RECT 205.090 38.805 205.260 38.975 ;
        RECT 205.090 38.445 205.260 38.615 ;
        RECT 210.380 39.165 210.550 39.335 ;
        RECT 210.380 38.805 210.550 38.975 ;
        RECT 210.380 38.445 210.550 38.615 ;
        RECT 205.090 34.055 205.260 34.225 ;
        RECT 205.090 33.695 205.260 33.865 ;
        RECT 205.090 33.335 205.260 33.505 ;
        RECT 205.090 32.975 205.260 33.145 ;
        RECT 210.380 34.055 210.550 34.225 ;
        RECT 210.380 33.695 210.550 33.865 ;
        RECT 210.380 33.335 210.550 33.505 ;
        RECT 210.380 32.975 210.550 33.145 ;
        RECT 205.090 28.585 205.260 28.755 ;
        RECT 205.090 28.225 205.260 28.395 ;
        RECT 169.630 27.615 169.800 27.785 ;
        RECT 169.630 27.255 169.800 27.425 ;
        RECT 169.630 26.895 169.800 27.065 ;
        RECT 169.630 26.535 169.800 26.705 ;
        RECT 169.630 26.175 169.800 26.345 ;
        RECT 202.080 27.615 202.250 27.785 ;
        RECT 202.080 27.255 202.250 27.425 ;
        RECT 202.080 26.895 202.250 27.065 ;
        RECT 202.080 26.535 202.250 26.705 ;
        RECT 202.080 26.175 202.250 26.345 ;
        RECT 96.190 17.255 96.360 17.425 ;
        RECT 96.190 16.895 96.360 17.065 ;
        RECT 101.480 17.255 101.650 17.425 ;
        RECT 85.610 16.535 85.780 16.705 ;
        RECT 90.900 16.535 91.070 16.705 ;
        RECT 96.190 16.535 96.360 16.705 ;
        RECT 101.480 16.895 101.650 17.065 ;
        RECT 101.480 16.535 101.650 16.705 ;
        RECT -96.485 11.700 -96.315 11.870 ;
        RECT -95.195 11.700 -95.025 11.870 ;
        RECT -93.905 11.700 -93.735 11.870 ;
        RECT -92.615 11.700 -92.445 11.870 ;
        RECT -91.325 11.700 -91.155 11.870 ;
        RECT -90.035 11.700 -89.865 11.870 ;
        RECT -88.745 11.700 -88.575 11.870 ;
        RECT -87.455 11.700 -87.285 11.870 ;
        RECT -86.165 11.700 -85.995 11.870 ;
        RECT -84.875 11.700 -84.705 11.870 ;
        RECT -83.585 11.700 -83.415 11.870 ;
        RECT -82.295 11.700 -82.125 11.870 ;
        RECT -81.005 11.700 -80.835 11.870 ;
        RECT -79.715 11.700 -79.545 11.870 ;
        RECT -78.425 11.700 -78.255 11.870 ;
        RECT -77.135 11.700 -76.965 11.870 ;
        RECT -75.845 11.700 -75.675 11.870 ;
        RECT -74.555 11.700 -74.385 11.870 ;
        RECT -73.265 11.700 -73.095 11.870 ;
        RECT -71.975 11.700 -71.805 11.870 ;
        RECT -90.700 8.825 -77.210 11.155 ;
        RECT 205.090 27.865 205.260 28.035 ;
        RECT 205.090 27.505 205.260 27.675 ;
        RECT 210.380 28.585 210.550 28.755 ;
        RECT 210.380 28.225 210.550 28.395 ;
        RECT 210.380 27.865 210.550 28.035 ;
        RECT 210.380 27.505 210.550 27.675 ;
        RECT 205.090 23.115 205.260 23.285 ;
        RECT 205.090 22.755 205.260 22.925 ;
        RECT 205.090 22.395 205.260 22.565 ;
        RECT 205.090 22.035 205.260 22.205 ;
        RECT 210.380 23.115 210.550 23.285 ;
        RECT 210.380 22.755 210.550 22.925 ;
        RECT 210.380 22.395 210.550 22.565 ;
        RECT 210.380 22.035 210.550 22.205 ;
        RECT 205.090 17.645 205.260 17.815 ;
        RECT 210.380 17.645 210.550 17.815 ;
        RECT 215.670 39.165 215.840 39.335 ;
        RECT 215.670 38.805 215.840 38.975 ;
        RECT 215.670 38.445 215.840 38.615 ;
        RECT 215.670 34.055 215.840 34.225 ;
        RECT 215.670 33.695 215.840 33.865 ;
        RECT 215.670 33.335 215.840 33.505 ;
        RECT 215.670 32.975 215.840 33.145 ;
        RECT 215.670 28.585 215.840 28.755 ;
        RECT 215.670 28.225 215.840 28.395 ;
        RECT 215.670 27.865 215.840 28.035 ;
        RECT 215.670 27.505 215.840 27.675 ;
        RECT 215.670 23.115 215.840 23.285 ;
        RECT 215.670 22.755 215.840 22.925 ;
        RECT 215.670 22.395 215.840 22.565 ;
        RECT 215.670 22.035 215.840 22.205 ;
        RECT 215.670 17.645 215.840 17.815 ;
        RECT 231.540 39.525 231.710 39.695 ;
        RECT 220.960 39.165 221.130 39.335 ;
        RECT 220.960 38.805 221.130 38.975 ;
        RECT 220.960 38.445 221.130 38.615 ;
        RECT 220.960 34.055 221.130 34.225 ;
        RECT 220.960 33.695 221.130 33.865 ;
        RECT 220.960 33.335 221.130 33.505 ;
        RECT 220.960 32.975 221.130 33.145 ;
        RECT 220.960 28.585 221.130 28.755 ;
        RECT 220.960 28.225 221.130 28.395 ;
        RECT 220.960 27.865 221.130 28.035 ;
        RECT 220.960 27.505 221.130 27.675 ;
        RECT 220.960 23.115 221.130 23.285 ;
        RECT 220.960 22.755 221.130 22.925 ;
        RECT 220.960 22.395 221.130 22.565 ;
        RECT 220.960 22.035 221.130 22.205 ;
        RECT 220.960 17.645 221.130 17.815 ;
        RECT 226.250 39.165 226.420 39.335 ;
        RECT 226.250 38.805 226.420 38.975 ;
        RECT 231.540 39.165 231.710 39.335 ;
        RECT 231.540 38.805 231.710 38.975 ;
        RECT 226.250 38.445 226.420 38.615 ;
        RECT 226.250 34.055 226.420 34.225 ;
        RECT 226.250 33.695 226.420 33.865 ;
        RECT 226.250 33.335 226.420 33.505 ;
        RECT 226.250 32.975 226.420 33.145 ;
        RECT 226.250 28.585 226.420 28.755 ;
        RECT 226.250 28.225 226.420 28.395 ;
        RECT 226.250 27.865 226.420 28.035 ;
        RECT 226.250 27.505 226.420 27.675 ;
        RECT 226.250 23.115 226.420 23.285 ;
        RECT 226.250 22.755 226.420 22.925 ;
        RECT 226.250 22.395 226.420 22.565 ;
        RECT 226.250 22.035 226.420 22.205 ;
        RECT 205.090 17.285 205.260 17.455 ;
        RECT 205.090 16.925 205.260 17.095 ;
        RECT 210.380 17.285 210.550 17.455 ;
        RECT 205.090 16.565 205.260 16.735 ;
        RECT 210.380 16.925 210.550 17.095 ;
        RECT 215.670 17.285 215.840 17.455 ;
        RECT 210.380 16.565 210.550 16.735 ;
        RECT 215.670 16.925 215.840 17.095 ;
        RECT 226.250 17.645 226.420 17.815 ;
        RECT 231.540 38.445 231.710 38.615 ;
        RECT 231.540 34.055 231.710 34.225 ;
        RECT 231.540 33.695 231.710 33.865 ;
        RECT 231.540 33.335 231.710 33.505 ;
        RECT 231.540 32.975 231.710 33.145 ;
        RECT 231.540 28.585 231.710 28.755 ;
        RECT 231.540 28.225 231.710 28.395 ;
        RECT 231.540 27.865 231.710 28.035 ;
        RECT 231.540 27.505 231.710 27.675 ;
        RECT 237.940 69.175 238.110 69.345 ;
        RECT 237.940 68.815 238.110 68.985 ;
        RECT 243.230 69.175 243.400 69.345 ;
        RECT 248.520 69.175 248.690 69.345 ;
        RECT 253.810 69.175 253.980 69.345 ;
        RECT 259.100 69.175 259.270 69.345 ;
        RECT 237.940 68.455 238.110 68.625 ;
        RECT 237.940 68.095 238.110 68.265 ;
        RECT 243.230 68.815 243.400 68.985 ;
        RECT 243.230 68.455 243.400 68.625 ;
        RECT 243.230 68.095 243.400 68.265 ;
        RECT 237.940 63.705 238.110 63.875 ;
        RECT 237.940 63.345 238.110 63.515 ;
        RECT 237.940 62.985 238.110 63.155 ;
        RECT 237.940 62.625 238.110 62.795 ;
        RECT 243.230 63.705 243.400 63.875 ;
        RECT 243.230 63.345 243.400 63.515 ;
        RECT 243.230 62.985 243.400 63.155 ;
        RECT 243.230 62.625 243.400 62.795 ;
        RECT 237.940 58.235 238.110 58.405 ;
        RECT 237.940 57.875 238.110 58.045 ;
        RECT 237.940 57.515 238.110 57.685 ;
        RECT 237.940 57.155 238.110 57.325 ;
        RECT 243.230 58.235 243.400 58.405 ;
        RECT 243.230 57.875 243.400 58.045 ;
        RECT 243.230 57.515 243.400 57.685 ;
        RECT 243.230 57.155 243.400 57.325 ;
        RECT 237.940 52.765 238.110 52.935 ;
        RECT 237.940 52.405 238.110 52.575 ;
        RECT 237.940 52.045 238.110 52.215 ;
        RECT 237.940 51.685 238.110 51.855 ;
        RECT 243.230 52.765 243.400 52.935 ;
        RECT 243.230 52.405 243.400 52.575 ;
        RECT 243.230 52.045 243.400 52.215 ;
        RECT 243.230 51.685 243.400 51.855 ;
        RECT 237.940 47.295 238.110 47.465 ;
        RECT 243.230 47.295 243.400 47.465 ;
        RECT 248.520 68.815 248.690 68.985 ;
        RECT 248.520 68.455 248.690 68.625 ;
        RECT 248.520 68.095 248.690 68.265 ;
        RECT 248.520 63.705 248.690 63.875 ;
        RECT 248.520 63.345 248.690 63.515 ;
        RECT 248.520 62.985 248.690 63.155 ;
        RECT 248.520 62.625 248.690 62.795 ;
        RECT 248.520 58.235 248.690 58.405 ;
        RECT 248.520 57.875 248.690 58.045 ;
        RECT 248.520 57.515 248.690 57.685 ;
        RECT 248.520 57.155 248.690 57.325 ;
        RECT 248.520 52.765 248.690 52.935 ;
        RECT 248.520 52.405 248.690 52.575 ;
        RECT 248.520 52.045 248.690 52.215 ;
        RECT 248.520 51.685 248.690 51.855 ;
        RECT 248.520 47.295 248.690 47.465 ;
        RECT 264.390 69.175 264.560 69.345 ;
        RECT 253.810 68.815 253.980 68.985 ;
        RECT 253.810 68.455 253.980 68.625 ;
        RECT 253.810 68.095 253.980 68.265 ;
        RECT 253.810 63.705 253.980 63.875 ;
        RECT 253.810 63.345 253.980 63.515 ;
        RECT 253.810 62.985 253.980 63.155 ;
        RECT 253.810 62.625 253.980 62.795 ;
        RECT 253.810 58.235 253.980 58.405 ;
        RECT 253.810 57.875 253.980 58.045 ;
        RECT 253.810 57.515 253.980 57.685 ;
        RECT 253.810 57.155 253.980 57.325 ;
        RECT 253.810 52.765 253.980 52.935 ;
        RECT 253.810 52.405 253.980 52.575 ;
        RECT 253.810 52.045 253.980 52.215 ;
        RECT 253.810 51.685 253.980 51.855 ;
        RECT 253.810 47.295 253.980 47.465 ;
        RECT 259.100 68.815 259.270 68.985 ;
        RECT 259.100 68.455 259.270 68.625 ;
        RECT 259.100 68.095 259.270 68.265 ;
        RECT 259.100 63.705 259.270 63.875 ;
        RECT 259.100 63.345 259.270 63.515 ;
        RECT 259.100 62.985 259.270 63.155 ;
        RECT 259.100 62.625 259.270 62.795 ;
        RECT 259.100 58.235 259.270 58.405 ;
        RECT 259.100 57.875 259.270 58.045 ;
        RECT 259.100 57.515 259.270 57.685 ;
        RECT 259.100 57.155 259.270 57.325 ;
        RECT 259.100 52.765 259.270 52.935 ;
        RECT 259.100 52.405 259.270 52.575 ;
        RECT 259.100 52.045 259.270 52.215 ;
        RECT 259.100 51.685 259.270 51.855 ;
        RECT 237.940 46.935 238.110 47.105 ;
        RECT 237.940 46.575 238.110 46.745 ;
        RECT 243.230 46.935 243.400 47.105 ;
        RECT 237.940 46.215 238.110 46.385 ;
        RECT 243.230 46.575 243.400 46.745 ;
        RECT 248.520 46.935 248.690 47.105 ;
        RECT 243.230 46.215 243.400 46.385 ;
        RECT 248.520 46.575 248.690 46.745 ;
        RECT 259.100 47.295 259.270 47.465 ;
        RECT 264.390 68.815 264.560 68.985 ;
        RECT 264.390 68.455 264.560 68.625 ;
        RECT 264.390 68.095 264.560 68.265 ;
        RECT 264.390 63.705 264.560 63.875 ;
        RECT 264.390 63.345 264.560 63.515 ;
        RECT 264.390 62.985 264.560 63.155 ;
        RECT 264.390 62.625 264.560 62.795 ;
        RECT 264.390 58.235 264.560 58.405 ;
        RECT 264.390 57.875 264.560 58.045 ;
        RECT 264.390 57.515 264.560 57.685 ;
        RECT 264.390 57.155 264.560 57.325 ;
        RECT 264.390 52.765 264.560 52.935 ;
        RECT 264.390 52.405 264.560 52.575 ;
        RECT 264.390 52.045 264.560 52.215 ;
        RECT 264.390 51.685 264.560 51.855 ;
        RECT 253.810 46.935 253.980 47.105 ;
        RECT 253.810 46.575 253.980 46.745 ;
        RECT 264.390 47.295 264.560 47.465 ;
        RECT 270.460 98.165 270.630 98.335 ;
        RECT 281.040 98.525 281.210 98.695 ;
        RECT 286.330 98.525 286.500 98.695 ;
        RECT 291.620 98.525 291.790 98.695 ;
        RECT 270.460 97.805 270.630 97.975 ;
        RECT 270.460 97.445 270.630 97.615 ;
        RECT 275.750 98.165 275.920 98.335 ;
        RECT 275.750 97.805 275.920 97.975 ;
        RECT 275.750 97.445 275.920 97.615 ;
        RECT 270.460 93.055 270.630 93.225 ;
        RECT 270.460 92.695 270.630 92.865 ;
        RECT 270.460 92.335 270.630 92.505 ;
        RECT 270.460 91.975 270.630 92.145 ;
        RECT 275.750 93.055 275.920 93.225 ;
        RECT 275.750 92.695 275.920 92.865 ;
        RECT 275.750 92.335 275.920 92.505 ;
        RECT 275.750 91.975 275.920 92.145 ;
        RECT 270.460 87.585 270.630 87.755 ;
        RECT 270.460 87.225 270.630 87.395 ;
        RECT 270.460 86.865 270.630 87.035 ;
        RECT 270.460 86.505 270.630 86.675 ;
        RECT 275.750 87.585 275.920 87.755 ;
        RECT 275.750 87.225 275.920 87.395 ;
        RECT 275.750 86.865 275.920 87.035 ;
        RECT 275.750 86.505 275.920 86.675 ;
        RECT 270.460 82.115 270.630 82.285 ;
        RECT 270.460 81.755 270.630 81.925 ;
        RECT 270.460 81.395 270.630 81.565 ;
        RECT 270.460 81.035 270.630 81.205 ;
        RECT 275.750 82.115 275.920 82.285 ;
        RECT 275.750 81.755 275.920 81.925 ;
        RECT 275.750 81.395 275.920 81.565 ;
        RECT 275.750 81.035 275.920 81.205 ;
        RECT 270.460 76.645 270.630 76.815 ;
        RECT 275.750 76.645 275.920 76.815 ;
        RECT 281.040 98.165 281.210 98.335 ;
        RECT 281.040 97.805 281.210 97.975 ;
        RECT 281.040 97.445 281.210 97.615 ;
        RECT 281.040 93.055 281.210 93.225 ;
        RECT 281.040 92.695 281.210 92.865 ;
        RECT 281.040 92.335 281.210 92.505 ;
        RECT 281.040 91.975 281.210 92.145 ;
        RECT 281.040 87.585 281.210 87.755 ;
        RECT 281.040 87.225 281.210 87.395 ;
        RECT 281.040 86.865 281.210 87.035 ;
        RECT 281.040 86.505 281.210 86.675 ;
        RECT 281.040 82.115 281.210 82.285 ;
        RECT 281.040 81.755 281.210 81.925 ;
        RECT 281.040 81.395 281.210 81.565 ;
        RECT 281.040 81.035 281.210 81.205 ;
        RECT 281.040 76.645 281.210 76.815 ;
        RECT 296.910 98.525 297.080 98.695 ;
        RECT 286.330 98.165 286.500 98.335 ;
        RECT 286.330 97.805 286.500 97.975 ;
        RECT 286.330 97.445 286.500 97.615 ;
        RECT 286.330 93.055 286.500 93.225 ;
        RECT 286.330 92.695 286.500 92.865 ;
        RECT 286.330 92.335 286.500 92.505 ;
        RECT 286.330 91.975 286.500 92.145 ;
        RECT 286.330 87.585 286.500 87.755 ;
        RECT 286.330 87.225 286.500 87.395 ;
        RECT 286.330 86.865 286.500 87.035 ;
        RECT 286.330 86.505 286.500 86.675 ;
        RECT 286.330 82.115 286.500 82.285 ;
        RECT 286.330 81.755 286.500 81.925 ;
        RECT 286.330 81.395 286.500 81.565 ;
        RECT 286.330 81.035 286.500 81.205 ;
        RECT 286.330 76.645 286.500 76.815 ;
        RECT 291.620 98.165 291.790 98.335 ;
        RECT 291.620 97.805 291.790 97.975 ;
        RECT 291.620 97.445 291.790 97.615 ;
        RECT 291.620 93.055 291.790 93.225 ;
        RECT 291.620 92.695 291.790 92.865 ;
        RECT 291.620 92.335 291.790 92.505 ;
        RECT 291.620 91.975 291.790 92.145 ;
        RECT 291.620 87.585 291.790 87.755 ;
        RECT 291.620 87.225 291.790 87.395 ;
        RECT 291.620 86.865 291.790 87.035 ;
        RECT 291.620 86.505 291.790 86.675 ;
        RECT 291.620 82.115 291.790 82.285 ;
        RECT 291.620 81.755 291.790 81.925 ;
        RECT 291.620 81.395 291.790 81.565 ;
        RECT 291.620 81.035 291.790 81.205 ;
        RECT 270.460 76.285 270.630 76.455 ;
        RECT 270.460 75.925 270.630 76.095 ;
        RECT 275.750 76.285 275.920 76.455 ;
        RECT 270.460 75.565 270.630 75.735 ;
        RECT 275.750 75.925 275.920 76.095 ;
        RECT 281.040 76.285 281.210 76.455 ;
        RECT 275.750 75.565 275.920 75.735 ;
        RECT 281.040 75.925 281.210 76.095 ;
        RECT 291.620 76.645 291.790 76.815 ;
        RECT 296.910 98.165 297.080 98.335 ;
        RECT 296.910 97.805 297.080 97.975 ;
        RECT 296.910 97.445 297.080 97.615 ;
        RECT 310.590 98.375 310.760 98.545 ;
        RECT 310.590 98.015 310.760 98.185 ;
        RECT 315.880 98.375 316.050 98.545 ;
        RECT 321.170 98.375 321.340 98.545 ;
        RECT 326.460 98.375 326.630 98.545 ;
        RECT 331.750 98.375 331.920 98.545 ;
        RECT 310.590 97.655 310.760 97.825 ;
        RECT 310.590 97.295 310.760 97.465 ;
        RECT 315.880 98.015 316.050 98.185 ;
        RECT 315.880 97.655 316.050 97.825 ;
        RECT 315.880 97.295 316.050 97.465 ;
        RECT 296.910 93.055 297.080 93.225 ;
        RECT 296.910 92.695 297.080 92.865 ;
        RECT 296.910 92.335 297.080 92.505 ;
        RECT 296.910 91.975 297.080 92.145 ;
        RECT 296.910 87.585 297.080 87.755 ;
        RECT 296.910 87.225 297.080 87.395 ;
        RECT 296.910 86.865 297.080 87.035 ;
        RECT 296.910 86.505 297.080 86.675 ;
        RECT 298.530 84.925 299.420 92.295 ;
        RECT 310.590 92.905 310.760 93.075 ;
        RECT 310.590 92.545 310.760 92.715 ;
        RECT 310.590 92.185 310.760 92.355 ;
        RECT 310.590 91.825 310.760 91.995 ;
        RECT 315.880 92.905 316.050 93.075 ;
        RECT 315.880 92.545 316.050 92.715 ;
        RECT 315.880 92.185 316.050 92.355 ;
        RECT 315.880 91.825 316.050 91.995 ;
        RECT 307.580 90.785 307.750 90.955 ;
        RECT 307.580 90.425 307.750 90.595 ;
        RECT 307.580 90.065 307.750 90.235 ;
        RECT 307.580 89.705 307.750 89.875 ;
        RECT 307.580 89.345 307.750 89.515 ;
        RECT 307.580 88.985 307.750 89.155 ;
        RECT 307.580 88.625 307.750 88.795 ;
        RECT 307.580 88.265 307.750 88.435 ;
        RECT 307.580 87.905 307.750 88.075 ;
        RECT 307.580 87.545 307.750 87.715 ;
        RECT 307.580 87.185 307.750 87.355 ;
        RECT 307.580 86.825 307.750 86.995 ;
        RECT 307.580 86.465 307.750 86.635 ;
        RECT 307.580 86.105 307.750 86.275 ;
        RECT 307.580 85.745 307.750 85.915 ;
        RECT 307.580 85.385 307.750 85.555 ;
        RECT 307.580 85.025 307.750 85.195 ;
        RECT 310.590 87.435 310.760 87.605 ;
        RECT 310.590 87.075 310.760 87.245 ;
        RECT 310.590 86.715 310.760 86.885 ;
        RECT 310.590 86.355 310.760 86.525 ;
        RECT 315.880 87.435 316.050 87.605 ;
        RECT 315.880 87.075 316.050 87.245 ;
        RECT 315.880 86.715 316.050 86.885 ;
        RECT 315.880 86.355 316.050 86.525 ;
        RECT 296.910 82.115 297.080 82.285 ;
        RECT 296.910 81.755 297.080 81.925 ;
        RECT 296.910 81.395 297.080 81.565 ;
        RECT 296.910 81.035 297.080 81.205 ;
        RECT 286.330 76.285 286.500 76.455 ;
        RECT 286.330 75.925 286.500 76.095 ;
        RECT 296.910 76.645 297.080 76.815 ;
        RECT 310.590 81.965 310.760 82.135 ;
        RECT 310.590 81.605 310.760 81.775 ;
        RECT 310.590 81.245 310.760 81.415 ;
        RECT 310.590 80.885 310.760 81.055 ;
        RECT 315.880 81.965 316.050 82.135 ;
        RECT 315.880 81.605 316.050 81.775 ;
        RECT 315.880 81.245 316.050 81.415 ;
        RECT 315.880 80.885 316.050 81.055 ;
        RECT 291.620 76.285 291.790 76.455 ;
        RECT 291.620 75.925 291.790 76.095 ;
        RECT 310.590 76.495 310.760 76.665 ;
        RECT 296.910 76.285 297.080 76.455 ;
        RECT 281.040 75.565 281.210 75.735 ;
        RECT 286.330 75.565 286.500 75.735 ;
        RECT 291.620 75.565 291.790 75.735 ;
        RECT 296.910 75.925 297.080 76.095 ;
        RECT 315.880 76.495 316.050 76.665 ;
        RECT 321.170 98.015 321.340 98.185 ;
        RECT 321.170 97.655 321.340 97.825 ;
        RECT 321.170 97.295 321.340 97.465 ;
        RECT 321.170 92.905 321.340 93.075 ;
        RECT 321.170 92.545 321.340 92.715 ;
        RECT 321.170 92.185 321.340 92.355 ;
        RECT 321.170 91.825 321.340 91.995 ;
        RECT 321.170 87.435 321.340 87.605 ;
        RECT 321.170 87.075 321.340 87.245 ;
        RECT 321.170 86.715 321.340 86.885 ;
        RECT 321.170 86.355 321.340 86.525 ;
        RECT 321.170 81.965 321.340 82.135 ;
        RECT 321.170 81.605 321.340 81.775 ;
        RECT 321.170 81.245 321.340 81.415 ;
        RECT 321.170 80.885 321.340 81.055 ;
        RECT 321.170 76.495 321.340 76.665 ;
        RECT 337.040 98.375 337.210 98.545 ;
        RECT 326.460 98.015 326.630 98.185 ;
        RECT 326.460 97.655 326.630 97.825 ;
        RECT 326.460 97.295 326.630 97.465 ;
        RECT 326.460 92.905 326.630 93.075 ;
        RECT 326.460 92.545 326.630 92.715 ;
        RECT 326.460 92.185 326.630 92.355 ;
        RECT 326.460 91.825 326.630 91.995 ;
        RECT 326.460 87.435 326.630 87.605 ;
        RECT 326.460 87.075 326.630 87.245 ;
        RECT 326.460 86.715 326.630 86.885 ;
        RECT 326.460 86.355 326.630 86.525 ;
        RECT 326.460 81.965 326.630 82.135 ;
        RECT 326.460 81.605 326.630 81.775 ;
        RECT 326.460 81.245 326.630 81.415 ;
        RECT 326.460 80.885 326.630 81.055 ;
        RECT 326.460 76.495 326.630 76.665 ;
        RECT 331.750 98.015 331.920 98.185 ;
        RECT 331.750 97.655 331.920 97.825 ;
        RECT 331.750 97.295 331.920 97.465 ;
        RECT 331.750 92.905 331.920 93.075 ;
        RECT 331.750 92.545 331.920 92.715 ;
        RECT 331.750 92.185 331.920 92.355 ;
        RECT 331.750 91.825 331.920 91.995 ;
        RECT 331.750 87.435 331.920 87.605 ;
        RECT 331.750 87.075 331.920 87.245 ;
        RECT 331.750 86.715 331.920 86.885 ;
        RECT 331.750 86.355 331.920 86.525 ;
        RECT 331.750 81.965 331.920 82.135 ;
        RECT 331.750 81.605 331.920 81.775 ;
        RECT 331.750 81.245 331.920 81.415 ;
        RECT 331.750 80.885 331.920 81.055 ;
        RECT 310.590 76.135 310.760 76.305 ;
        RECT 296.910 75.565 297.080 75.735 ;
        RECT 310.590 75.775 310.760 75.945 ;
        RECT 315.880 76.135 316.050 76.305 ;
        RECT 310.590 75.415 310.760 75.585 ;
        RECT 315.880 75.775 316.050 75.945 ;
        RECT 321.170 76.135 321.340 76.305 ;
        RECT 315.880 75.415 316.050 75.585 ;
        RECT 321.170 75.775 321.340 75.945 ;
        RECT 331.750 76.495 331.920 76.665 ;
        RECT 337.040 98.015 337.210 98.185 ;
        RECT 337.040 97.655 337.210 97.825 ;
        RECT 337.040 97.295 337.210 97.465 ;
        RECT 337.040 92.905 337.210 93.075 ;
        RECT 337.040 92.545 337.210 92.715 ;
        RECT 337.040 92.185 337.210 92.355 ;
        RECT 337.040 91.825 337.210 91.995 ;
        RECT 337.040 87.435 337.210 87.605 ;
        RECT 337.040 87.075 337.210 87.245 ;
        RECT 337.040 86.715 337.210 86.885 ;
        RECT 337.040 86.355 337.210 86.525 ;
        RECT 337.040 81.965 337.210 82.135 ;
        RECT 337.040 81.605 337.210 81.775 ;
        RECT 337.040 81.245 337.210 81.415 ;
        RECT 337.040 80.885 337.210 81.055 ;
        RECT 326.460 76.135 326.630 76.305 ;
        RECT 326.460 75.775 326.630 75.945 ;
        RECT 337.040 76.495 337.210 76.665 ;
        RECT 342.870 126.475 343.040 126.645 ;
        RECT 348.160 127.195 348.330 127.365 ;
        RECT 348.160 126.835 348.330 127.005 ;
        RECT 348.160 126.475 348.330 126.645 ;
        RECT 342.870 122.085 343.040 122.255 ;
        RECT 342.870 121.725 343.040 121.895 ;
        RECT 342.870 121.365 343.040 121.535 ;
        RECT 342.870 121.005 343.040 121.175 ;
        RECT 348.160 122.085 348.330 122.255 ;
        RECT 348.160 121.725 348.330 121.895 ;
        RECT 348.160 121.365 348.330 121.535 ;
        RECT 348.160 121.005 348.330 121.175 ;
        RECT 342.870 116.615 343.040 116.785 ;
        RECT 342.870 116.255 343.040 116.425 ;
        RECT 342.870 115.895 343.040 116.065 ;
        RECT 342.870 115.535 343.040 115.705 ;
        RECT 348.160 116.615 348.330 116.785 ;
        RECT 348.160 116.255 348.330 116.425 ;
        RECT 348.160 115.895 348.330 116.065 ;
        RECT 348.160 115.535 348.330 115.705 ;
        RECT 342.870 111.145 343.040 111.315 ;
        RECT 342.870 110.785 343.040 110.955 ;
        RECT 342.870 110.425 343.040 110.595 ;
        RECT 342.870 110.065 343.040 110.235 ;
        RECT 348.160 111.145 348.330 111.315 ;
        RECT 348.160 110.785 348.330 110.955 ;
        RECT 348.160 110.425 348.330 110.595 ;
        RECT 348.160 110.065 348.330 110.235 ;
        RECT 342.870 105.675 343.040 105.845 ;
        RECT 348.160 105.675 348.330 105.845 ;
        RECT 353.450 127.195 353.620 127.365 ;
        RECT 353.450 126.835 353.620 127.005 ;
        RECT 353.450 126.475 353.620 126.645 ;
        RECT 353.450 122.085 353.620 122.255 ;
        RECT 353.450 121.725 353.620 121.895 ;
        RECT 353.450 121.365 353.620 121.535 ;
        RECT 353.450 121.005 353.620 121.175 ;
        RECT 353.450 116.615 353.620 116.785 ;
        RECT 353.450 116.255 353.620 116.425 ;
        RECT 353.450 115.895 353.620 116.065 ;
        RECT 353.450 115.535 353.620 115.705 ;
        RECT 353.450 111.145 353.620 111.315 ;
        RECT 353.450 110.785 353.620 110.955 ;
        RECT 353.450 110.425 353.620 110.595 ;
        RECT 353.450 110.065 353.620 110.235 ;
        RECT 353.450 105.675 353.620 105.845 ;
        RECT 369.320 127.555 369.490 127.725 ;
        RECT 358.740 127.195 358.910 127.365 ;
        RECT 358.740 126.835 358.910 127.005 ;
        RECT 358.740 126.475 358.910 126.645 ;
        RECT 358.740 122.085 358.910 122.255 ;
        RECT 358.740 121.725 358.910 121.895 ;
        RECT 358.740 121.365 358.910 121.535 ;
        RECT 358.740 121.005 358.910 121.175 ;
        RECT 358.740 116.615 358.910 116.785 ;
        RECT 358.740 116.255 358.910 116.425 ;
        RECT 358.740 115.895 358.910 116.065 ;
        RECT 358.740 115.535 358.910 115.705 ;
        RECT 358.740 111.145 358.910 111.315 ;
        RECT 358.740 110.785 358.910 110.955 ;
        RECT 358.740 110.425 358.910 110.595 ;
        RECT 358.740 110.065 358.910 110.235 ;
        RECT 358.740 105.675 358.910 105.845 ;
        RECT 364.030 127.195 364.200 127.365 ;
        RECT 364.030 126.835 364.200 127.005 ;
        RECT 364.030 126.475 364.200 126.645 ;
        RECT 364.030 122.085 364.200 122.255 ;
        RECT 364.030 121.725 364.200 121.895 ;
        RECT 364.030 121.365 364.200 121.535 ;
        RECT 364.030 121.005 364.200 121.175 ;
        RECT 364.030 116.615 364.200 116.785 ;
        RECT 364.030 116.255 364.200 116.425 ;
        RECT 364.030 115.895 364.200 116.065 ;
        RECT 364.030 115.535 364.200 115.705 ;
        RECT 364.030 111.145 364.200 111.315 ;
        RECT 364.030 110.785 364.200 110.955 ;
        RECT 364.030 110.425 364.200 110.595 ;
        RECT 364.030 110.065 364.200 110.235 ;
        RECT 342.870 105.315 343.040 105.485 ;
        RECT 342.870 104.955 343.040 105.125 ;
        RECT 348.160 105.315 348.330 105.485 ;
        RECT 342.870 104.595 343.040 104.765 ;
        RECT 348.160 104.955 348.330 105.125 ;
        RECT 353.450 105.315 353.620 105.485 ;
        RECT 348.160 104.595 348.330 104.765 ;
        RECT 353.450 104.955 353.620 105.125 ;
        RECT 364.030 105.675 364.200 105.845 ;
        RECT 369.320 127.195 369.490 127.365 ;
        RECT 381.630 127.425 381.800 127.595 ;
        RECT 369.320 126.835 369.490 127.005 ;
        RECT 369.320 126.475 369.490 126.645 ;
        RECT 381.630 127.065 381.800 127.235 ;
        RECT 392.210 127.425 392.380 127.595 ;
        RECT 402.790 127.425 402.960 127.595 ;
        RECT 413.940 127.415 414.110 127.585 ;
        RECT 381.630 126.705 381.800 126.875 ;
        RECT 381.630 126.345 381.800 126.515 ;
        RECT 369.320 122.085 369.490 122.255 ;
        RECT 369.320 121.725 369.490 121.895 ;
        RECT 369.320 121.365 369.490 121.535 ;
        RECT 369.320 121.005 369.490 121.175 ;
        RECT 369.320 116.615 369.490 116.785 ;
        RECT 369.320 116.255 369.490 116.425 ;
        RECT 369.320 115.895 369.490 116.065 ;
        RECT 369.320 115.535 369.490 115.705 ;
        RECT 369.320 111.145 369.490 111.315 ;
        RECT 369.320 110.785 369.490 110.955 ;
        RECT 369.320 110.425 369.490 110.595 ;
        RECT 369.320 110.065 369.490 110.235 ;
        RECT 358.740 105.315 358.910 105.485 ;
        RECT 358.740 104.955 358.910 105.125 ;
        RECT 369.320 105.675 369.490 105.845 ;
        RECT 373.330 119.835 373.500 120.005 ;
        RECT 373.330 119.475 373.500 119.645 ;
        RECT 373.330 119.115 373.500 119.285 ;
        RECT 373.330 118.755 373.500 118.925 ;
        RECT 373.330 118.395 373.500 118.565 ;
        RECT 373.330 118.035 373.500 118.205 ;
        RECT 373.330 117.675 373.500 117.845 ;
        RECT 373.330 117.315 373.500 117.485 ;
        RECT 373.330 116.955 373.500 117.125 ;
        RECT 373.330 116.595 373.500 116.765 ;
        RECT 373.330 116.235 373.500 116.405 ;
        RECT 373.330 115.875 373.500 116.045 ;
        RECT 373.330 115.515 373.500 115.685 ;
        RECT 373.330 115.155 373.500 115.325 ;
        RECT 373.330 114.795 373.500 114.965 ;
        RECT 373.330 114.435 373.500 114.605 ;
        RECT 373.330 114.075 373.500 114.245 ;
        RECT 364.030 105.315 364.200 105.485 ;
        RECT 364.030 104.955 364.200 105.125 ;
        RECT 369.320 105.315 369.490 105.485 ;
        RECT 353.450 104.595 353.620 104.765 ;
        RECT 358.740 104.595 358.910 104.765 ;
        RECT 364.030 104.595 364.200 104.765 ;
        RECT 369.320 104.955 369.490 105.125 ;
        RECT 369.320 104.595 369.490 104.765 ;
        RECT 339.900 90.845 340.070 91.015 ;
        RECT 339.900 90.485 340.070 90.655 ;
        RECT 339.900 90.125 340.070 90.295 ;
        RECT 339.900 89.765 340.070 89.935 ;
        RECT 339.900 89.405 340.070 89.575 ;
        RECT 339.900 89.045 340.070 89.215 ;
        RECT 339.900 88.685 340.070 88.855 ;
        RECT 339.900 88.325 340.070 88.495 ;
        RECT 339.900 87.965 340.070 88.135 ;
        RECT 339.900 87.605 340.070 87.775 ;
        RECT 339.900 87.245 340.070 87.415 ;
        RECT 339.900 86.885 340.070 87.055 ;
        RECT 339.900 86.525 340.070 86.695 ;
        RECT 339.900 86.165 340.070 86.335 ;
        RECT 339.900 85.805 340.070 85.975 ;
        RECT 339.900 85.445 340.070 85.615 ;
        RECT 339.900 85.085 340.070 85.255 ;
        RECT 331.750 76.135 331.920 76.305 ;
        RECT 331.750 75.775 331.920 75.945 ;
        RECT 337.040 76.135 337.210 76.305 ;
        RECT 321.170 75.415 321.340 75.585 ;
        RECT 326.460 75.415 326.630 75.585 ;
        RECT 331.750 75.415 331.920 75.585 ;
        RECT 337.040 75.775 337.210 75.945 ;
        RECT 337.040 75.415 337.210 75.585 ;
        RECT 267.500 61.655 267.670 61.825 ;
        RECT 267.500 61.295 267.670 61.465 ;
        RECT 267.500 60.935 267.670 61.105 ;
        RECT 267.500 60.575 267.670 60.745 ;
        RECT 267.500 60.215 267.670 60.385 ;
        RECT 267.500 59.855 267.670 60.025 ;
        RECT 267.500 59.495 267.670 59.665 ;
        RECT 267.500 59.135 267.670 59.305 ;
        RECT 267.500 58.775 267.670 58.945 ;
        RECT 267.500 58.415 267.670 58.585 ;
        RECT 267.500 58.055 267.670 58.225 ;
        RECT 267.500 57.695 267.670 57.865 ;
        RECT 267.500 57.335 267.670 57.505 ;
        RECT 267.500 56.975 267.670 57.145 ;
        RECT 267.500 56.615 267.670 56.785 ;
        RECT 267.500 56.255 267.670 56.425 ;
        RECT 267.500 55.895 267.670 56.065 ;
        RECT 259.100 46.935 259.270 47.105 ;
        RECT 259.100 46.575 259.270 46.745 ;
        RECT 264.390 46.935 264.560 47.105 ;
        RECT 248.520 46.215 248.690 46.385 ;
        RECT 253.810 46.215 253.980 46.385 ;
        RECT 259.100 46.215 259.270 46.385 ;
        RECT 264.390 46.575 264.560 46.745 ;
        RECT 264.390 46.215 264.560 46.385 ;
        RECT 235.020 32.045 235.190 32.215 ;
        RECT 235.020 31.685 235.190 31.855 ;
        RECT 235.020 31.325 235.190 31.495 ;
        RECT 235.020 30.965 235.190 31.135 ;
        RECT 235.020 30.605 235.190 30.775 ;
        RECT 235.020 30.245 235.190 30.415 ;
        RECT 235.020 29.885 235.190 30.055 ;
        RECT 235.020 29.525 235.190 29.695 ;
        RECT 235.020 29.165 235.190 29.335 ;
        RECT 235.020 28.805 235.190 28.975 ;
        RECT 235.020 28.445 235.190 28.615 ;
        RECT 235.020 28.085 235.190 28.255 ;
        RECT 235.020 27.725 235.190 27.895 ;
        RECT 235.020 27.365 235.190 27.535 ;
        RECT 235.020 27.005 235.190 27.175 ;
        RECT 238.030 39.635 238.200 39.805 ;
        RECT 238.030 39.275 238.200 39.445 ;
        RECT 243.320 39.635 243.490 39.805 ;
        RECT 248.610 39.635 248.780 39.805 ;
        RECT 253.900 39.635 254.070 39.805 ;
        RECT 259.190 39.635 259.360 39.805 ;
        RECT 238.030 38.915 238.200 39.085 ;
        RECT 238.030 38.555 238.200 38.725 ;
        RECT 243.320 39.275 243.490 39.445 ;
        RECT 243.320 38.915 243.490 39.085 ;
        RECT 243.320 38.555 243.490 38.725 ;
        RECT 238.030 34.165 238.200 34.335 ;
        RECT 238.030 33.805 238.200 33.975 ;
        RECT 238.030 33.445 238.200 33.615 ;
        RECT 238.030 33.085 238.200 33.255 ;
        RECT 243.320 34.165 243.490 34.335 ;
        RECT 243.320 33.805 243.490 33.975 ;
        RECT 243.320 33.445 243.490 33.615 ;
        RECT 243.320 33.085 243.490 33.255 ;
        RECT 238.030 28.695 238.200 28.865 ;
        RECT 238.030 28.335 238.200 28.505 ;
        RECT 238.030 27.975 238.200 28.145 ;
        RECT 238.030 27.615 238.200 27.785 ;
        RECT 243.320 28.695 243.490 28.865 ;
        RECT 243.320 28.335 243.490 28.505 ;
        RECT 243.320 27.975 243.490 28.145 ;
        RECT 243.320 27.615 243.490 27.785 ;
        RECT 235.020 26.645 235.190 26.815 ;
        RECT 235.020 26.285 235.190 26.455 ;
        RECT 231.540 23.115 231.710 23.285 ;
        RECT 231.540 22.755 231.710 22.925 ;
        RECT 231.540 22.395 231.710 22.565 ;
        RECT 231.540 22.035 231.710 22.205 ;
        RECT 220.960 17.285 221.130 17.455 ;
        RECT 220.960 16.925 221.130 17.095 ;
        RECT 231.540 17.645 231.710 17.815 ;
        RECT 238.030 23.225 238.200 23.395 ;
        RECT 238.030 22.865 238.200 23.035 ;
        RECT 238.030 22.505 238.200 22.675 ;
        RECT 238.030 22.145 238.200 22.315 ;
        RECT 243.320 23.225 243.490 23.395 ;
        RECT 243.320 22.865 243.490 23.035 ;
        RECT 243.320 22.505 243.490 22.675 ;
        RECT 243.320 22.145 243.490 22.315 ;
        RECT 238.030 17.755 238.200 17.925 ;
        RECT 226.250 17.285 226.420 17.455 ;
        RECT 226.250 16.925 226.420 17.095 ;
        RECT 231.540 17.285 231.710 17.455 ;
        RECT 215.670 16.565 215.840 16.735 ;
        RECT 220.960 16.565 221.130 16.735 ;
        RECT 226.250 16.565 226.420 16.735 ;
        RECT 231.540 16.925 231.710 17.095 ;
        RECT 243.320 17.755 243.490 17.925 ;
        RECT 248.610 39.275 248.780 39.445 ;
        RECT 248.610 38.915 248.780 39.085 ;
        RECT 248.610 38.555 248.780 38.725 ;
        RECT 248.610 34.165 248.780 34.335 ;
        RECT 248.610 33.805 248.780 33.975 ;
        RECT 248.610 33.445 248.780 33.615 ;
        RECT 248.610 33.085 248.780 33.255 ;
        RECT 248.610 28.695 248.780 28.865 ;
        RECT 248.610 28.335 248.780 28.505 ;
        RECT 248.610 27.975 248.780 28.145 ;
        RECT 248.610 27.615 248.780 27.785 ;
        RECT 248.610 23.225 248.780 23.395 ;
        RECT 248.610 22.865 248.780 23.035 ;
        RECT 248.610 22.505 248.780 22.675 ;
        RECT 248.610 22.145 248.780 22.315 ;
        RECT 248.610 17.755 248.780 17.925 ;
        RECT 264.480 39.635 264.650 39.805 ;
        RECT 253.900 39.275 254.070 39.445 ;
        RECT 253.900 38.915 254.070 39.085 ;
        RECT 253.900 38.555 254.070 38.725 ;
        RECT 253.900 34.165 254.070 34.335 ;
        RECT 253.900 33.805 254.070 33.975 ;
        RECT 253.900 33.445 254.070 33.615 ;
        RECT 253.900 33.085 254.070 33.255 ;
        RECT 253.900 28.695 254.070 28.865 ;
        RECT 253.900 28.335 254.070 28.505 ;
        RECT 253.900 27.975 254.070 28.145 ;
        RECT 253.900 27.615 254.070 27.785 ;
        RECT 253.900 23.225 254.070 23.395 ;
        RECT 253.900 22.865 254.070 23.035 ;
        RECT 253.900 22.505 254.070 22.675 ;
        RECT 253.900 22.145 254.070 22.315 ;
        RECT 253.900 17.755 254.070 17.925 ;
        RECT 259.190 39.275 259.360 39.445 ;
        RECT 259.190 38.915 259.360 39.085 ;
        RECT 264.480 39.275 264.650 39.445 ;
        RECT 259.190 38.555 259.360 38.725 ;
        RECT 259.190 34.165 259.360 34.335 ;
        RECT 259.190 33.805 259.360 33.975 ;
        RECT 259.190 33.445 259.360 33.615 ;
        RECT 259.190 33.085 259.360 33.255 ;
        RECT 259.190 28.695 259.360 28.865 ;
        RECT 259.190 28.335 259.360 28.505 ;
        RECT 259.190 27.975 259.360 28.145 ;
        RECT 259.190 27.615 259.360 27.785 ;
        RECT 259.190 23.225 259.360 23.395 ;
        RECT 259.190 22.865 259.360 23.035 ;
        RECT 259.190 22.505 259.360 22.675 ;
        RECT 259.190 22.145 259.360 22.315 ;
        RECT 238.030 17.395 238.200 17.565 ;
        RECT 238.030 17.035 238.200 17.205 ;
        RECT 243.320 17.395 243.490 17.565 ;
        RECT 231.540 16.565 231.710 16.735 ;
        RECT 238.030 16.675 238.200 16.845 ;
        RECT 243.320 17.035 243.490 17.205 ;
        RECT 248.610 17.395 248.780 17.565 ;
        RECT 243.320 16.675 243.490 16.845 ;
        RECT 248.610 17.035 248.780 17.205 ;
        RECT 259.190 17.755 259.360 17.925 ;
        RECT 264.480 38.915 264.650 39.085 ;
        RECT 264.480 38.555 264.650 38.725 ;
        RECT 264.480 34.165 264.650 34.335 ;
        RECT 264.480 33.805 264.650 33.975 ;
        RECT 264.480 33.445 264.650 33.615 ;
        RECT 264.480 33.085 264.650 33.255 ;
        RECT 264.480 28.695 264.650 28.865 ;
        RECT 264.480 28.335 264.650 28.505 ;
        RECT 264.480 27.975 264.650 28.145 ;
        RECT 264.480 27.615 264.650 27.785 ;
        RECT 270.510 69.245 270.680 69.415 ;
        RECT 270.510 68.885 270.680 69.055 ;
        RECT 275.800 69.245 275.970 69.415 ;
        RECT 281.090 69.245 281.260 69.415 ;
        RECT 286.380 69.245 286.550 69.415 ;
        RECT 291.670 69.245 291.840 69.415 ;
        RECT 270.510 68.525 270.680 68.695 ;
        RECT 270.510 68.165 270.680 68.335 ;
        RECT 275.800 68.885 275.970 69.055 ;
        RECT 275.800 68.525 275.970 68.695 ;
        RECT 275.800 68.165 275.970 68.335 ;
        RECT 270.510 63.775 270.680 63.945 ;
        RECT 270.510 63.415 270.680 63.585 ;
        RECT 270.510 63.055 270.680 63.225 ;
        RECT 270.510 62.695 270.680 62.865 ;
        RECT 275.800 63.775 275.970 63.945 ;
        RECT 275.800 63.415 275.970 63.585 ;
        RECT 275.800 63.055 275.970 63.225 ;
        RECT 275.800 62.695 275.970 62.865 ;
        RECT 270.510 58.305 270.680 58.475 ;
        RECT 270.510 57.945 270.680 58.115 ;
        RECT 270.510 57.585 270.680 57.755 ;
        RECT 270.510 57.225 270.680 57.395 ;
        RECT 275.800 58.305 275.970 58.475 ;
        RECT 275.800 57.945 275.970 58.115 ;
        RECT 275.800 57.585 275.970 57.755 ;
        RECT 275.800 57.225 275.970 57.395 ;
        RECT 270.510 52.835 270.680 53.005 ;
        RECT 270.510 52.475 270.680 52.645 ;
        RECT 270.510 52.115 270.680 52.285 ;
        RECT 270.510 51.755 270.680 51.925 ;
        RECT 275.800 52.835 275.970 53.005 ;
        RECT 275.800 52.475 275.970 52.645 ;
        RECT 275.800 52.115 275.970 52.285 ;
        RECT 275.800 51.755 275.970 51.925 ;
        RECT 270.510 47.365 270.680 47.535 ;
        RECT 275.800 47.365 275.970 47.535 ;
        RECT 281.090 68.885 281.260 69.055 ;
        RECT 281.090 68.525 281.260 68.695 ;
        RECT 281.090 68.165 281.260 68.335 ;
        RECT 281.090 63.775 281.260 63.945 ;
        RECT 281.090 63.415 281.260 63.585 ;
        RECT 281.090 63.055 281.260 63.225 ;
        RECT 281.090 62.695 281.260 62.865 ;
        RECT 281.090 58.305 281.260 58.475 ;
        RECT 281.090 57.945 281.260 58.115 ;
        RECT 281.090 57.585 281.260 57.755 ;
        RECT 281.090 57.225 281.260 57.395 ;
        RECT 281.090 52.835 281.260 53.005 ;
        RECT 281.090 52.475 281.260 52.645 ;
        RECT 281.090 52.115 281.260 52.285 ;
        RECT 281.090 51.755 281.260 51.925 ;
        RECT 281.090 47.365 281.260 47.535 ;
        RECT 296.960 69.245 297.130 69.415 ;
        RECT 286.380 68.885 286.550 69.055 ;
        RECT 286.380 68.525 286.550 68.695 ;
        RECT 286.380 68.165 286.550 68.335 ;
        RECT 286.380 63.775 286.550 63.945 ;
        RECT 286.380 63.415 286.550 63.585 ;
        RECT 286.380 63.055 286.550 63.225 ;
        RECT 286.380 62.695 286.550 62.865 ;
        RECT 286.380 58.305 286.550 58.475 ;
        RECT 286.380 57.945 286.550 58.115 ;
        RECT 286.380 57.585 286.550 57.755 ;
        RECT 286.380 57.225 286.550 57.395 ;
        RECT 286.380 52.835 286.550 53.005 ;
        RECT 286.380 52.475 286.550 52.645 ;
        RECT 286.380 52.115 286.550 52.285 ;
        RECT 286.380 51.755 286.550 51.925 ;
        RECT 286.380 47.365 286.550 47.535 ;
        RECT 291.670 68.885 291.840 69.055 ;
        RECT 291.670 68.525 291.840 68.695 ;
        RECT 291.670 68.165 291.840 68.335 ;
        RECT 291.670 63.775 291.840 63.945 ;
        RECT 291.670 63.415 291.840 63.585 ;
        RECT 291.670 63.055 291.840 63.225 ;
        RECT 291.670 62.695 291.840 62.865 ;
        RECT 291.670 58.305 291.840 58.475 ;
        RECT 291.670 57.945 291.840 58.115 ;
        RECT 291.670 57.585 291.840 57.755 ;
        RECT 291.670 57.225 291.840 57.395 ;
        RECT 291.670 52.835 291.840 53.005 ;
        RECT 291.670 52.475 291.840 52.645 ;
        RECT 291.670 52.115 291.840 52.285 ;
        RECT 291.670 51.755 291.840 51.925 ;
        RECT 270.510 47.005 270.680 47.175 ;
        RECT 270.510 46.645 270.680 46.815 ;
        RECT 275.800 47.005 275.970 47.175 ;
        RECT 270.510 46.285 270.680 46.455 ;
        RECT 275.800 46.645 275.970 46.815 ;
        RECT 281.090 47.005 281.260 47.175 ;
        RECT 275.800 46.285 275.970 46.455 ;
        RECT 281.090 46.645 281.260 46.815 ;
        RECT 291.670 47.365 291.840 47.535 ;
        RECT 296.960 68.885 297.130 69.055 ;
        RECT 310.590 69.085 310.760 69.255 ;
        RECT 296.960 68.525 297.130 68.695 ;
        RECT 296.960 68.165 297.130 68.335 ;
        RECT 296.960 63.775 297.130 63.945 ;
        RECT 296.960 63.415 297.130 63.585 ;
        RECT 310.590 68.725 310.760 68.895 ;
        RECT 315.880 69.085 316.050 69.255 ;
        RECT 321.170 69.085 321.340 69.255 ;
        RECT 326.460 69.085 326.630 69.255 ;
        RECT 331.750 69.085 331.920 69.255 ;
        RECT 310.590 68.365 310.760 68.535 ;
        RECT 310.590 68.005 310.760 68.175 ;
        RECT 315.880 68.725 316.050 68.895 ;
        RECT 315.880 68.365 316.050 68.535 ;
        RECT 315.880 68.005 316.050 68.175 ;
        RECT 310.590 63.615 310.760 63.785 ;
        RECT 296.960 63.055 297.130 63.225 ;
        RECT 296.960 62.695 297.130 62.865 ;
        RECT 296.960 58.305 297.130 58.475 ;
        RECT 296.960 57.945 297.130 58.115 ;
        RECT 296.960 57.585 297.130 57.755 ;
        RECT 296.960 57.225 297.130 57.395 ;
        RECT 298.635 55.950 299.525 62.600 ;
        RECT 310.590 63.255 310.760 63.425 ;
        RECT 310.590 62.895 310.760 63.065 ;
        RECT 310.590 62.535 310.760 62.705 ;
        RECT 315.880 63.615 316.050 63.785 ;
        RECT 315.880 63.255 316.050 63.425 ;
        RECT 315.880 62.895 316.050 63.065 ;
        RECT 315.880 62.535 316.050 62.705 ;
        RECT 307.580 61.495 307.750 61.665 ;
        RECT 307.580 61.135 307.750 61.305 ;
        RECT 307.580 60.775 307.750 60.945 ;
        RECT 307.580 60.415 307.750 60.585 ;
        RECT 307.580 60.055 307.750 60.225 ;
        RECT 307.580 59.695 307.750 59.865 ;
        RECT 307.580 59.335 307.750 59.505 ;
        RECT 307.580 58.975 307.750 59.145 ;
        RECT 307.580 58.615 307.750 58.785 ;
        RECT 307.580 58.255 307.750 58.425 ;
        RECT 307.580 57.895 307.750 58.065 ;
        RECT 307.580 57.535 307.750 57.705 ;
        RECT 307.580 57.175 307.750 57.345 ;
        RECT 307.580 56.815 307.750 56.985 ;
        RECT 307.580 56.455 307.750 56.625 ;
        RECT 307.580 56.095 307.750 56.265 ;
        RECT 307.580 55.735 307.750 55.905 ;
        RECT 310.590 58.145 310.760 58.315 ;
        RECT 310.590 57.785 310.760 57.955 ;
        RECT 310.590 57.425 310.760 57.595 ;
        RECT 310.590 57.065 310.760 57.235 ;
        RECT 315.880 58.145 316.050 58.315 ;
        RECT 315.880 57.785 316.050 57.955 ;
        RECT 315.880 57.425 316.050 57.595 ;
        RECT 315.880 57.065 316.050 57.235 ;
        RECT 296.960 52.835 297.130 53.005 ;
        RECT 296.960 52.475 297.130 52.645 ;
        RECT 296.960 52.115 297.130 52.285 ;
        RECT 296.960 51.755 297.130 51.925 ;
        RECT 286.380 47.005 286.550 47.175 ;
        RECT 286.380 46.645 286.550 46.815 ;
        RECT 296.960 47.365 297.130 47.535 ;
        RECT 310.590 52.675 310.760 52.845 ;
        RECT 310.590 52.315 310.760 52.485 ;
        RECT 310.590 51.955 310.760 52.125 ;
        RECT 310.590 51.595 310.760 51.765 ;
        RECT 315.880 52.675 316.050 52.845 ;
        RECT 315.880 52.315 316.050 52.485 ;
        RECT 315.880 51.955 316.050 52.125 ;
        RECT 315.880 51.595 316.050 51.765 ;
        RECT 291.670 47.005 291.840 47.175 ;
        RECT 291.670 46.645 291.840 46.815 ;
        RECT 310.590 47.205 310.760 47.375 ;
        RECT 296.960 47.005 297.130 47.175 ;
        RECT 281.090 46.285 281.260 46.455 ;
        RECT 286.380 46.285 286.550 46.455 ;
        RECT 291.670 46.285 291.840 46.455 ;
        RECT 296.960 46.645 297.130 46.815 ;
        RECT 315.880 47.205 316.050 47.375 ;
        RECT 321.170 68.725 321.340 68.895 ;
        RECT 321.170 68.365 321.340 68.535 ;
        RECT 321.170 68.005 321.340 68.175 ;
        RECT 321.170 63.615 321.340 63.785 ;
        RECT 321.170 63.255 321.340 63.425 ;
        RECT 321.170 62.895 321.340 63.065 ;
        RECT 321.170 62.535 321.340 62.705 ;
        RECT 321.170 58.145 321.340 58.315 ;
        RECT 321.170 57.785 321.340 57.955 ;
        RECT 321.170 57.425 321.340 57.595 ;
        RECT 321.170 57.065 321.340 57.235 ;
        RECT 321.170 52.675 321.340 52.845 ;
        RECT 321.170 52.315 321.340 52.485 ;
        RECT 321.170 51.955 321.340 52.125 ;
        RECT 321.170 51.595 321.340 51.765 ;
        RECT 321.170 47.205 321.340 47.375 ;
        RECT 337.040 69.085 337.210 69.255 ;
        RECT 326.460 68.725 326.630 68.895 ;
        RECT 326.460 68.365 326.630 68.535 ;
        RECT 326.460 68.005 326.630 68.175 ;
        RECT 326.460 63.615 326.630 63.785 ;
        RECT 326.460 63.255 326.630 63.425 ;
        RECT 326.460 62.895 326.630 63.065 ;
        RECT 326.460 62.535 326.630 62.705 ;
        RECT 326.460 58.145 326.630 58.315 ;
        RECT 326.460 57.785 326.630 57.955 ;
        RECT 326.460 57.425 326.630 57.595 ;
        RECT 326.460 57.065 326.630 57.235 ;
        RECT 326.460 52.675 326.630 52.845 ;
        RECT 326.460 52.315 326.630 52.485 ;
        RECT 326.460 51.955 326.630 52.125 ;
        RECT 326.460 51.595 326.630 51.765 ;
        RECT 326.460 47.205 326.630 47.375 ;
        RECT 331.750 68.725 331.920 68.895 ;
        RECT 331.750 68.365 331.920 68.535 ;
        RECT 331.750 68.005 331.920 68.175 ;
        RECT 331.750 63.615 331.920 63.785 ;
        RECT 331.750 63.255 331.920 63.425 ;
        RECT 331.750 62.895 331.920 63.065 ;
        RECT 331.750 62.535 331.920 62.705 ;
        RECT 331.750 58.145 331.920 58.315 ;
        RECT 331.750 57.785 331.920 57.955 ;
        RECT 331.750 57.425 331.920 57.595 ;
        RECT 331.750 57.065 331.920 57.235 ;
        RECT 331.750 52.675 331.920 52.845 ;
        RECT 331.750 52.315 331.920 52.485 ;
        RECT 331.750 51.955 331.920 52.125 ;
        RECT 331.750 51.595 331.920 51.765 ;
        RECT 310.590 46.845 310.760 47.015 ;
        RECT 296.960 46.285 297.130 46.455 ;
        RECT 310.590 46.485 310.760 46.655 ;
        RECT 315.880 46.845 316.050 47.015 ;
        RECT 310.590 46.125 310.760 46.295 ;
        RECT 315.880 46.485 316.050 46.655 ;
        RECT 321.170 46.845 321.340 47.015 ;
        RECT 315.880 46.125 316.050 46.295 ;
        RECT 321.170 46.485 321.340 46.655 ;
        RECT 331.750 47.205 331.920 47.375 ;
        RECT 337.040 68.725 337.210 68.895 ;
        RECT 337.040 68.365 337.210 68.535 ;
        RECT 337.040 68.005 337.210 68.175 ;
        RECT 337.040 63.615 337.210 63.785 ;
        RECT 337.040 63.255 337.210 63.425 ;
        RECT 337.040 62.895 337.210 63.065 ;
        RECT 337.040 62.535 337.210 62.705 ;
        RECT 337.040 58.145 337.210 58.315 ;
        RECT 337.040 57.785 337.210 57.955 ;
        RECT 337.040 57.425 337.210 57.595 ;
        RECT 337.040 57.065 337.210 57.235 ;
        RECT 337.040 52.675 337.210 52.845 ;
        RECT 337.040 52.315 337.210 52.485 ;
        RECT 337.040 51.955 337.210 52.125 ;
        RECT 337.040 51.595 337.210 51.765 ;
        RECT 326.460 46.845 326.630 47.015 ;
        RECT 326.460 46.485 326.630 46.655 ;
        RECT 337.040 47.205 337.210 47.375 ;
        RECT 342.910 98.435 343.080 98.605 ;
        RECT 342.910 98.075 343.080 98.245 ;
        RECT 348.200 98.435 348.370 98.605 ;
        RECT 353.490 98.435 353.660 98.605 ;
        RECT 358.780 98.435 358.950 98.605 ;
        RECT 364.070 98.435 364.240 98.605 ;
        RECT 342.910 97.715 343.080 97.885 ;
        RECT 342.910 97.355 343.080 97.525 ;
        RECT 348.200 98.075 348.370 98.245 ;
        RECT 348.200 97.715 348.370 97.885 ;
        RECT 348.200 97.355 348.370 97.525 ;
        RECT 342.910 92.965 343.080 93.135 ;
        RECT 342.910 92.605 343.080 92.775 ;
        RECT 342.910 92.245 343.080 92.415 ;
        RECT 342.910 91.885 343.080 92.055 ;
        RECT 348.200 92.965 348.370 93.135 ;
        RECT 348.200 92.605 348.370 92.775 ;
        RECT 348.200 92.245 348.370 92.415 ;
        RECT 348.200 91.885 348.370 92.055 ;
        RECT 342.910 87.495 343.080 87.665 ;
        RECT 342.910 87.135 343.080 87.305 ;
        RECT 342.910 86.775 343.080 86.945 ;
        RECT 342.910 86.415 343.080 86.585 ;
        RECT 348.200 87.495 348.370 87.665 ;
        RECT 348.200 87.135 348.370 87.305 ;
        RECT 348.200 86.775 348.370 86.945 ;
        RECT 348.200 86.415 348.370 86.585 ;
        RECT 342.910 82.025 343.080 82.195 ;
        RECT 342.910 81.665 343.080 81.835 ;
        RECT 342.910 81.305 343.080 81.475 ;
        RECT 342.910 80.945 343.080 81.115 ;
        RECT 348.200 82.025 348.370 82.195 ;
        RECT 348.200 81.665 348.370 81.835 ;
        RECT 348.200 81.305 348.370 81.475 ;
        RECT 348.200 80.945 348.370 81.115 ;
        RECT 342.910 76.555 343.080 76.725 ;
        RECT 348.200 76.555 348.370 76.725 ;
        RECT 353.490 98.075 353.660 98.245 ;
        RECT 353.490 97.715 353.660 97.885 ;
        RECT 353.490 97.355 353.660 97.525 ;
        RECT 353.490 92.965 353.660 93.135 ;
        RECT 353.490 92.605 353.660 92.775 ;
        RECT 353.490 92.245 353.660 92.415 ;
        RECT 353.490 91.885 353.660 92.055 ;
        RECT 353.490 87.495 353.660 87.665 ;
        RECT 353.490 87.135 353.660 87.305 ;
        RECT 353.490 86.775 353.660 86.945 ;
        RECT 353.490 86.415 353.660 86.585 ;
        RECT 353.490 82.025 353.660 82.195 ;
        RECT 353.490 81.665 353.660 81.835 ;
        RECT 353.490 81.305 353.660 81.475 ;
        RECT 353.490 80.945 353.660 81.115 ;
        RECT 353.490 76.555 353.660 76.725 ;
        RECT 369.360 98.435 369.530 98.605 ;
        RECT 358.780 98.075 358.950 98.245 ;
        RECT 358.780 97.715 358.950 97.885 ;
        RECT 358.780 97.355 358.950 97.525 ;
        RECT 358.780 92.965 358.950 93.135 ;
        RECT 358.780 92.605 358.950 92.775 ;
        RECT 358.780 92.245 358.950 92.415 ;
        RECT 358.780 91.885 358.950 92.055 ;
        RECT 358.780 87.495 358.950 87.665 ;
        RECT 358.780 87.135 358.950 87.305 ;
        RECT 358.780 86.775 358.950 86.945 ;
        RECT 358.780 86.415 358.950 86.585 ;
        RECT 358.780 82.025 358.950 82.195 ;
        RECT 358.780 81.665 358.950 81.835 ;
        RECT 358.780 81.305 358.950 81.475 ;
        RECT 358.780 80.945 358.950 81.115 ;
        RECT 358.780 76.555 358.950 76.725 ;
        RECT 364.070 98.075 364.240 98.245 ;
        RECT 364.070 97.715 364.240 97.885 ;
        RECT 364.070 97.355 364.240 97.525 ;
        RECT 364.070 92.965 364.240 93.135 ;
        RECT 364.070 92.605 364.240 92.775 ;
        RECT 364.070 92.245 364.240 92.415 ;
        RECT 364.070 91.885 364.240 92.055 ;
        RECT 364.070 87.495 364.240 87.665 ;
        RECT 364.070 87.135 364.240 87.305 ;
        RECT 364.070 86.775 364.240 86.945 ;
        RECT 364.070 86.415 364.240 86.585 ;
        RECT 364.070 82.025 364.240 82.195 ;
        RECT 364.070 81.665 364.240 81.835 ;
        RECT 364.070 81.305 364.240 81.475 ;
        RECT 364.070 80.945 364.240 81.115 ;
        RECT 342.910 76.195 343.080 76.365 ;
        RECT 342.910 75.835 343.080 76.005 ;
        RECT 348.200 76.195 348.370 76.365 ;
        RECT 342.910 75.475 343.080 75.645 ;
        RECT 348.200 75.835 348.370 76.005 ;
        RECT 353.490 76.195 353.660 76.365 ;
        RECT 348.200 75.475 348.370 75.645 ;
        RECT 353.490 75.835 353.660 76.005 ;
        RECT 364.070 76.555 364.240 76.725 ;
        RECT 369.360 98.075 369.530 98.245 ;
        RECT 369.360 97.715 369.530 97.885 ;
        RECT 369.360 97.355 369.530 97.525 ;
        RECT 369.360 92.965 369.530 93.135 ;
        RECT 369.360 92.605 369.530 92.775 ;
        RECT 369.360 92.245 369.530 92.415 ;
        RECT 369.360 91.885 369.530 92.055 ;
        RECT 369.360 87.495 369.530 87.665 ;
        RECT 369.360 87.135 369.530 87.305 ;
        RECT 369.360 86.775 369.530 86.945 ;
        RECT 369.360 86.415 369.530 86.585 ;
        RECT 369.360 82.025 369.530 82.195 ;
        RECT 369.360 81.665 369.530 81.835 ;
        RECT 369.360 81.305 369.530 81.475 ;
        RECT 369.360 80.945 369.530 81.115 ;
        RECT 358.780 76.195 358.950 76.365 ;
        RECT 358.780 75.835 358.950 76.005 ;
        RECT 369.360 76.555 369.530 76.725 ;
        RECT 381.630 121.955 381.800 122.125 ;
        RECT 381.630 121.595 381.800 121.765 ;
        RECT 381.630 121.235 381.800 121.405 ;
        RECT 381.630 120.875 381.800 121.045 ;
        RECT 381.630 116.485 381.800 116.655 ;
        RECT 381.630 116.125 381.800 116.295 ;
        RECT 381.630 115.765 381.800 115.935 ;
        RECT 381.630 115.405 381.800 115.575 ;
        RECT 381.630 111.015 381.800 111.185 ;
        RECT 381.630 110.655 381.800 110.825 ;
        RECT 381.630 110.295 381.800 110.465 ;
        RECT 381.630 109.935 381.800 110.105 ;
        RECT 381.630 105.545 381.800 105.715 ;
        RECT 392.210 127.065 392.380 127.235 ;
        RECT 392.210 126.705 392.380 126.875 ;
        RECT 392.210 126.345 392.380 126.515 ;
        RECT 392.210 121.955 392.380 122.125 ;
        RECT 392.210 121.595 392.380 121.765 ;
        RECT 392.210 121.235 392.380 121.405 ;
        RECT 392.210 120.875 392.380 121.045 ;
        RECT 392.210 116.485 392.380 116.655 ;
        RECT 392.210 116.125 392.380 116.295 ;
        RECT 392.210 115.765 392.380 115.935 ;
        RECT 392.210 115.405 392.380 115.575 ;
        RECT 392.210 111.015 392.380 111.185 ;
        RECT 392.210 110.655 392.380 110.825 ;
        RECT 392.210 110.295 392.380 110.465 ;
        RECT 392.210 109.935 392.380 110.105 ;
        RECT 392.210 105.545 392.380 105.715 ;
        RECT 402.790 127.065 402.960 127.235 ;
        RECT 402.790 126.705 402.960 126.875 ;
        RECT 402.790 126.345 402.960 126.515 ;
        RECT 413.940 127.055 414.110 127.225 ;
        RECT 424.520 127.415 424.690 127.585 ;
        RECT 435.100 127.415 435.270 127.585 ;
        RECT 442.510 127.385 442.680 127.555 ;
        RECT 413.940 126.695 414.110 126.865 ;
        RECT 413.940 126.335 414.110 126.505 ;
        RECT 402.790 121.955 402.960 122.125 ;
        RECT 402.790 121.595 402.960 121.765 ;
        RECT 402.790 121.235 402.960 121.405 ;
        RECT 402.790 120.875 402.960 121.045 ;
        RECT 402.790 116.485 402.960 116.655 ;
        RECT 402.790 116.125 402.960 116.295 ;
        RECT 402.790 115.765 402.960 115.935 ;
        RECT 402.790 115.405 402.960 115.575 ;
        RECT 402.790 111.015 402.960 111.185 ;
        RECT 402.790 110.655 402.960 110.825 ;
        RECT 402.790 110.295 402.960 110.465 ;
        RECT 402.790 109.935 402.960 110.105 ;
        RECT 402.790 105.545 402.960 105.715 ;
        RECT 405.640 119.825 405.810 119.995 ;
        RECT 405.640 119.465 405.810 119.635 ;
        RECT 405.640 119.105 405.810 119.275 ;
        RECT 405.640 118.745 405.810 118.915 ;
        RECT 405.640 118.385 405.810 118.555 ;
        RECT 405.640 118.025 405.810 118.195 ;
        RECT 405.640 117.665 405.810 117.835 ;
        RECT 405.640 117.305 405.810 117.475 ;
        RECT 405.640 116.945 405.810 117.115 ;
        RECT 405.640 116.585 405.810 116.755 ;
        RECT 405.640 116.225 405.810 116.395 ;
        RECT 405.640 115.865 405.810 116.035 ;
        RECT 405.640 115.505 405.810 115.675 ;
        RECT 405.640 115.145 405.810 115.315 ;
        RECT 405.640 114.785 405.810 114.955 ;
        RECT 405.640 114.425 405.810 114.595 ;
        RECT 405.640 114.065 405.810 114.235 ;
        RECT 381.630 105.185 381.800 105.355 ;
        RECT 381.630 104.825 381.800 104.995 ;
        RECT 392.210 105.185 392.380 105.355 ;
        RECT 392.210 104.825 392.380 104.995 ;
        RECT 402.790 105.185 402.960 105.355 ;
        RECT 402.790 104.825 402.960 104.995 ;
        RECT 381.630 104.465 381.800 104.635 ;
        RECT 392.210 104.465 392.380 104.635 ;
        RECT 402.790 104.465 402.960 104.635 ;
        RECT 413.940 121.945 414.110 122.115 ;
        RECT 413.940 121.585 414.110 121.755 ;
        RECT 413.940 121.225 414.110 121.395 ;
        RECT 413.940 120.865 414.110 121.035 ;
        RECT 413.940 116.475 414.110 116.645 ;
        RECT 413.940 116.115 414.110 116.285 ;
        RECT 413.940 115.755 414.110 115.925 ;
        RECT 413.940 115.395 414.110 115.565 ;
        RECT 413.940 111.005 414.110 111.175 ;
        RECT 413.940 110.645 414.110 110.815 ;
        RECT 413.940 110.285 414.110 110.455 ;
        RECT 413.940 109.925 414.110 110.095 ;
        RECT 413.940 105.535 414.110 105.705 ;
        RECT 424.520 127.055 424.690 127.225 ;
        RECT 424.520 126.695 424.690 126.865 ;
        RECT 424.520 126.335 424.690 126.505 ;
        RECT 424.520 121.945 424.690 122.115 ;
        RECT 424.520 121.585 424.690 121.755 ;
        RECT 424.520 121.225 424.690 121.395 ;
        RECT 424.520 120.865 424.690 121.035 ;
        RECT 424.520 116.475 424.690 116.645 ;
        RECT 424.520 116.115 424.690 116.285 ;
        RECT 424.520 115.755 424.690 115.925 ;
        RECT 424.520 115.395 424.690 115.565 ;
        RECT 424.520 111.005 424.690 111.175 ;
        RECT 424.520 110.645 424.690 110.815 ;
        RECT 424.520 110.285 424.690 110.455 ;
        RECT 424.520 109.925 424.690 110.095 ;
        RECT 424.520 105.535 424.690 105.705 ;
        RECT 435.100 127.055 435.270 127.225 ;
        RECT 435.100 126.695 435.270 126.865 ;
        RECT 435.100 126.335 435.270 126.505 ;
        RECT 442.510 127.025 442.680 127.195 ;
        RECT 447.800 127.385 447.970 127.555 ;
        RECT 453.090 127.385 453.260 127.555 ;
        RECT 458.380 127.385 458.550 127.555 ;
        RECT 463.670 127.385 463.840 127.555 ;
        RECT 442.510 126.665 442.680 126.835 ;
        RECT 442.510 126.305 442.680 126.475 ;
        RECT 447.800 127.025 447.970 127.195 ;
        RECT 447.800 126.665 447.970 126.835 ;
        RECT 447.800 126.305 447.970 126.475 ;
        RECT 435.100 121.945 435.270 122.115 ;
        RECT 435.100 121.585 435.270 121.755 ;
        RECT 435.100 121.225 435.270 121.395 ;
        RECT 435.100 120.865 435.270 121.035 ;
        RECT 435.100 116.475 435.270 116.645 ;
        RECT 435.100 116.115 435.270 116.285 ;
        RECT 435.100 115.755 435.270 115.925 ;
        RECT 435.100 115.395 435.270 115.565 ;
        RECT 435.100 111.005 435.270 111.175 ;
        RECT 435.100 110.645 435.270 110.815 ;
        RECT 435.100 110.285 435.270 110.455 ;
        RECT 435.100 109.925 435.270 110.095 ;
        RECT 435.100 105.535 435.270 105.705 ;
        RECT 439.500 119.795 439.670 119.965 ;
        RECT 439.500 119.435 439.670 119.605 ;
        RECT 439.500 119.075 439.670 119.245 ;
        RECT 439.500 118.715 439.670 118.885 ;
        RECT 439.500 118.355 439.670 118.525 ;
        RECT 439.500 117.995 439.670 118.165 ;
        RECT 439.500 117.635 439.670 117.805 ;
        RECT 439.500 117.275 439.670 117.445 ;
        RECT 439.500 116.915 439.670 117.085 ;
        RECT 439.500 116.555 439.670 116.725 ;
        RECT 439.500 116.195 439.670 116.365 ;
        RECT 439.500 115.835 439.670 116.005 ;
        RECT 439.500 115.475 439.670 115.645 ;
        RECT 439.500 115.115 439.670 115.285 ;
        RECT 439.500 114.755 439.670 114.925 ;
        RECT 439.500 114.395 439.670 114.565 ;
        RECT 439.500 114.035 439.670 114.205 ;
        RECT 413.940 105.175 414.110 105.345 ;
        RECT 413.940 104.815 414.110 104.985 ;
        RECT 424.520 105.175 424.690 105.345 ;
        RECT 424.520 104.815 424.690 104.985 ;
        RECT 435.100 105.175 435.270 105.345 ;
        RECT 435.100 104.815 435.270 104.985 ;
        RECT 413.940 104.455 414.110 104.625 ;
        RECT 424.520 104.455 424.690 104.625 ;
        RECT 435.100 104.455 435.270 104.625 ;
        RECT 381.660 98.235 381.830 98.405 ;
        RECT 373.360 90.645 373.530 90.815 ;
        RECT 373.360 90.285 373.530 90.455 ;
        RECT 373.360 89.925 373.530 90.095 ;
        RECT 373.360 89.565 373.530 89.735 ;
        RECT 373.360 89.205 373.530 89.375 ;
        RECT 373.360 88.845 373.530 89.015 ;
        RECT 373.360 88.485 373.530 88.655 ;
        RECT 373.360 88.125 373.530 88.295 ;
        RECT 373.360 87.765 373.530 87.935 ;
        RECT 373.360 87.405 373.530 87.575 ;
        RECT 373.360 87.045 373.530 87.215 ;
        RECT 373.360 86.685 373.530 86.855 ;
        RECT 373.360 86.325 373.530 86.495 ;
        RECT 373.360 85.965 373.530 86.135 ;
        RECT 373.360 85.605 373.530 85.775 ;
        RECT 373.360 85.245 373.530 85.415 ;
        RECT 373.360 84.885 373.530 85.055 ;
        RECT 364.070 76.195 364.240 76.365 ;
        RECT 364.070 75.835 364.240 76.005 ;
        RECT 369.360 76.195 369.530 76.365 ;
        RECT 353.490 75.475 353.660 75.645 ;
        RECT 358.780 75.475 358.950 75.645 ;
        RECT 364.070 75.475 364.240 75.645 ;
        RECT 369.360 75.835 369.530 76.005 ;
        RECT 369.360 75.475 369.530 75.645 ;
        RECT 339.920 61.485 340.090 61.655 ;
        RECT 339.920 61.125 340.090 61.295 ;
        RECT 339.920 60.765 340.090 60.935 ;
        RECT 339.920 60.405 340.090 60.575 ;
        RECT 339.920 60.045 340.090 60.215 ;
        RECT 339.920 59.685 340.090 59.855 ;
        RECT 339.920 59.325 340.090 59.495 ;
        RECT 339.920 58.965 340.090 59.135 ;
        RECT 339.920 58.605 340.090 58.775 ;
        RECT 339.920 58.245 340.090 58.415 ;
        RECT 339.920 57.885 340.090 58.055 ;
        RECT 339.920 57.525 340.090 57.695 ;
        RECT 339.920 57.165 340.090 57.335 ;
        RECT 339.920 56.805 340.090 56.975 ;
        RECT 339.920 56.445 340.090 56.615 ;
        RECT 339.920 56.085 340.090 56.255 ;
        RECT 339.920 55.725 340.090 55.895 ;
        RECT 331.750 46.845 331.920 47.015 ;
        RECT 331.750 46.485 331.920 46.655 ;
        RECT 337.040 46.845 337.210 47.015 ;
        RECT 321.170 46.125 321.340 46.295 ;
        RECT 326.460 46.125 326.630 46.295 ;
        RECT 331.750 46.125 331.920 46.295 ;
        RECT 337.040 46.485 337.210 46.655 ;
        RECT 337.040 46.125 337.210 46.295 ;
        RECT 267.590 32.115 267.760 32.285 ;
        RECT 267.590 31.755 267.760 31.925 ;
        RECT 267.590 31.395 267.760 31.565 ;
        RECT 267.590 31.035 267.760 31.205 ;
        RECT 267.590 30.675 267.760 30.845 ;
        RECT 267.590 30.315 267.760 30.485 ;
        RECT 267.590 29.955 267.760 30.125 ;
        RECT 267.590 29.595 267.760 29.765 ;
        RECT 267.590 29.235 267.760 29.405 ;
        RECT 267.590 28.875 267.760 29.045 ;
        RECT 267.590 28.515 267.760 28.685 ;
        RECT 267.590 28.155 267.760 28.325 ;
        RECT 267.590 27.795 267.760 27.965 ;
        RECT 267.590 27.435 267.760 27.605 ;
        RECT 267.590 27.075 267.760 27.245 ;
        RECT 267.590 26.715 267.760 26.885 ;
        RECT 270.600 39.705 270.770 39.875 ;
        RECT 270.600 39.345 270.770 39.515 ;
        RECT 275.890 39.705 276.060 39.875 ;
        RECT 281.180 39.705 281.350 39.875 ;
        RECT 286.470 39.705 286.640 39.875 ;
        RECT 291.760 39.705 291.930 39.875 ;
        RECT 270.600 38.985 270.770 39.155 ;
        RECT 270.600 38.625 270.770 38.795 ;
        RECT 275.890 39.345 276.060 39.515 ;
        RECT 275.890 38.985 276.060 39.155 ;
        RECT 275.890 38.625 276.060 38.795 ;
        RECT 270.600 34.235 270.770 34.405 ;
        RECT 270.600 33.875 270.770 34.045 ;
        RECT 270.600 33.515 270.770 33.685 ;
        RECT 270.600 33.155 270.770 33.325 ;
        RECT 275.890 34.235 276.060 34.405 ;
        RECT 275.890 33.875 276.060 34.045 ;
        RECT 275.890 33.515 276.060 33.685 ;
        RECT 275.890 33.155 276.060 33.325 ;
        RECT 270.600 28.765 270.770 28.935 ;
        RECT 270.600 28.405 270.770 28.575 ;
        RECT 270.600 28.045 270.770 28.215 ;
        RECT 270.600 27.685 270.770 27.855 ;
        RECT 275.890 28.765 276.060 28.935 ;
        RECT 275.890 28.405 276.060 28.575 ;
        RECT 275.890 28.045 276.060 28.215 ;
        RECT 275.890 27.685 276.060 27.855 ;
        RECT 267.590 26.355 267.760 26.525 ;
        RECT 264.480 23.225 264.650 23.395 ;
        RECT 264.480 22.865 264.650 23.035 ;
        RECT 264.480 22.505 264.650 22.675 ;
        RECT 264.480 22.145 264.650 22.315 ;
        RECT 253.900 17.395 254.070 17.565 ;
        RECT 253.900 17.035 254.070 17.205 ;
        RECT 264.480 17.755 264.650 17.925 ;
        RECT 270.600 23.295 270.770 23.465 ;
        RECT 270.600 22.935 270.770 23.105 ;
        RECT 270.600 22.575 270.770 22.745 ;
        RECT 270.600 22.215 270.770 22.385 ;
        RECT 275.890 23.295 276.060 23.465 ;
        RECT 275.890 22.935 276.060 23.105 ;
        RECT 275.890 22.575 276.060 22.745 ;
        RECT 275.890 22.215 276.060 22.385 ;
        RECT 270.600 17.825 270.770 17.995 ;
        RECT 259.190 17.395 259.360 17.565 ;
        RECT 259.190 17.035 259.360 17.205 ;
        RECT 264.480 17.395 264.650 17.565 ;
        RECT 248.610 16.675 248.780 16.845 ;
        RECT 253.900 16.675 254.070 16.845 ;
        RECT 259.190 16.675 259.360 16.845 ;
        RECT 264.480 17.035 264.650 17.205 ;
        RECT 275.890 17.825 276.060 17.995 ;
        RECT 281.180 39.345 281.350 39.515 ;
        RECT 281.180 38.985 281.350 39.155 ;
        RECT 281.180 38.625 281.350 38.795 ;
        RECT 281.180 34.235 281.350 34.405 ;
        RECT 281.180 33.875 281.350 34.045 ;
        RECT 281.180 33.515 281.350 33.685 ;
        RECT 281.180 33.155 281.350 33.325 ;
        RECT 281.180 28.765 281.350 28.935 ;
        RECT 281.180 28.405 281.350 28.575 ;
        RECT 281.180 28.045 281.350 28.215 ;
        RECT 281.180 27.685 281.350 27.855 ;
        RECT 281.180 23.295 281.350 23.465 ;
        RECT 281.180 22.935 281.350 23.105 ;
        RECT 281.180 22.575 281.350 22.745 ;
        RECT 281.180 22.215 281.350 22.385 ;
        RECT 281.180 17.825 281.350 17.995 ;
        RECT 297.050 39.705 297.220 39.875 ;
        RECT 286.470 39.345 286.640 39.515 ;
        RECT 286.470 38.985 286.640 39.155 ;
        RECT 286.470 38.625 286.640 38.795 ;
        RECT 286.470 34.235 286.640 34.405 ;
        RECT 286.470 33.875 286.640 34.045 ;
        RECT 286.470 33.515 286.640 33.685 ;
        RECT 286.470 33.155 286.640 33.325 ;
        RECT 286.470 28.765 286.640 28.935 ;
        RECT 286.470 28.405 286.640 28.575 ;
        RECT 286.470 28.045 286.640 28.215 ;
        RECT 286.470 27.685 286.640 27.855 ;
        RECT 286.470 23.295 286.640 23.465 ;
        RECT 286.470 22.935 286.640 23.105 ;
        RECT 286.470 22.575 286.640 22.745 ;
        RECT 286.470 22.215 286.640 22.385 ;
        RECT 286.470 17.825 286.640 17.995 ;
        RECT 291.760 39.345 291.930 39.515 ;
        RECT 297.050 39.345 297.220 39.515 ;
        RECT 310.590 39.795 310.760 39.965 ;
        RECT 310.590 39.435 310.760 39.605 ;
        RECT 315.880 39.795 316.050 39.965 ;
        RECT 321.170 39.795 321.340 39.965 ;
        RECT 326.460 39.795 326.630 39.965 ;
        RECT 331.750 39.795 331.920 39.965 ;
        RECT 291.760 38.985 291.930 39.155 ;
        RECT 291.760 38.625 291.930 38.795 ;
        RECT 291.760 34.235 291.930 34.405 ;
        RECT 291.760 33.875 291.930 34.045 ;
        RECT 291.760 33.515 291.930 33.685 ;
        RECT 291.760 33.155 291.930 33.325 ;
        RECT 291.760 28.765 291.930 28.935 ;
        RECT 291.760 28.405 291.930 28.575 ;
        RECT 291.760 28.045 291.930 28.215 ;
        RECT 291.760 27.685 291.930 27.855 ;
        RECT 291.760 23.295 291.930 23.465 ;
        RECT 291.760 22.935 291.930 23.105 ;
        RECT 291.760 22.575 291.930 22.745 ;
        RECT 291.760 22.215 291.930 22.385 ;
        RECT 270.600 17.465 270.770 17.635 ;
        RECT 270.600 17.105 270.770 17.275 ;
        RECT 275.890 17.465 276.060 17.635 ;
        RECT 264.480 16.675 264.650 16.845 ;
        RECT 270.600 16.745 270.770 16.915 ;
        RECT 275.890 17.105 276.060 17.275 ;
        RECT 281.180 17.465 281.350 17.635 ;
        RECT 275.890 16.745 276.060 16.915 ;
        RECT 281.180 17.105 281.350 17.275 ;
        RECT 291.760 17.825 291.930 17.995 ;
        RECT 297.050 38.985 297.220 39.155 ;
        RECT 297.050 38.625 297.220 38.795 ;
        RECT 297.050 34.235 297.220 34.405 ;
        RECT 310.590 39.075 310.760 39.245 ;
        RECT 310.590 38.715 310.760 38.885 ;
        RECT 315.880 39.435 316.050 39.605 ;
        RECT 315.880 39.075 316.050 39.245 ;
        RECT 315.880 38.715 316.050 38.885 ;
        RECT 310.590 34.325 310.760 34.495 ;
        RECT 297.050 33.875 297.220 34.045 ;
        RECT 297.050 33.515 297.220 33.685 ;
        RECT 297.050 33.155 297.220 33.325 ;
        RECT 297.050 28.765 297.220 28.935 ;
        RECT 297.050 28.405 297.220 28.575 ;
        RECT 297.050 28.045 297.220 28.215 ;
        RECT 297.050 27.685 297.220 27.855 ;
        RECT 298.570 26.810 299.100 33.460 ;
        RECT 310.590 33.965 310.760 34.135 ;
        RECT 310.590 33.605 310.760 33.775 ;
        RECT 310.590 33.245 310.760 33.415 ;
        RECT 315.880 34.325 316.050 34.495 ;
        RECT 315.880 33.965 316.050 34.135 ;
        RECT 315.880 33.605 316.050 33.775 ;
        RECT 315.880 33.245 316.050 33.415 ;
        RECT 307.580 32.205 307.750 32.375 ;
        RECT 307.580 31.845 307.750 32.015 ;
        RECT 307.580 31.485 307.750 31.655 ;
        RECT 307.580 31.125 307.750 31.295 ;
        RECT 307.580 30.765 307.750 30.935 ;
        RECT 307.580 30.405 307.750 30.575 ;
        RECT 307.580 30.045 307.750 30.215 ;
        RECT 307.580 29.685 307.750 29.855 ;
        RECT 297.050 23.295 297.220 23.465 ;
        RECT 297.050 22.935 297.220 23.105 ;
        RECT 297.050 22.575 297.220 22.745 ;
        RECT 297.050 22.215 297.220 22.385 ;
        RECT 286.470 17.465 286.640 17.635 ;
        RECT 286.470 17.105 286.640 17.275 ;
        RECT 297.050 17.825 297.220 17.995 ;
        RECT 291.760 17.465 291.930 17.635 ;
        RECT 291.760 17.105 291.930 17.275 ;
        RECT 297.050 17.465 297.220 17.635 ;
        RECT 281.180 16.745 281.350 16.915 ;
        RECT 286.470 16.745 286.640 16.915 ;
        RECT 291.760 16.745 291.930 16.915 ;
        RECT 297.050 17.105 297.220 17.275 ;
        RECT 297.050 16.745 297.220 16.915 ;
        RECT 307.580 29.325 307.750 29.495 ;
        RECT 307.580 28.965 307.750 29.135 ;
        RECT 307.580 28.605 307.750 28.775 ;
        RECT 307.580 28.245 307.750 28.415 ;
        RECT 307.580 27.885 307.750 28.055 ;
        RECT 307.580 27.525 307.750 27.695 ;
        RECT 307.580 27.165 307.750 27.335 ;
        RECT 307.580 26.805 307.750 26.975 ;
        RECT 307.580 26.445 307.750 26.615 ;
        RECT 310.590 28.855 310.760 29.025 ;
        RECT 310.590 28.495 310.760 28.665 ;
        RECT 310.590 28.135 310.760 28.305 ;
        RECT 310.590 27.775 310.760 27.945 ;
        RECT 315.880 28.855 316.050 29.025 ;
        RECT 315.880 28.495 316.050 28.665 ;
        RECT 315.880 28.135 316.050 28.305 ;
        RECT 315.880 27.775 316.050 27.945 ;
        RECT 310.590 23.385 310.760 23.555 ;
        RECT 310.590 23.025 310.760 23.195 ;
        RECT 310.590 22.665 310.760 22.835 ;
        RECT 310.590 22.305 310.760 22.475 ;
        RECT 315.880 23.385 316.050 23.555 ;
        RECT 315.880 23.025 316.050 23.195 ;
        RECT 315.880 22.665 316.050 22.835 ;
        RECT 315.880 22.305 316.050 22.475 ;
        RECT 310.590 17.915 310.760 18.085 ;
        RECT 315.880 17.915 316.050 18.085 ;
        RECT 321.170 39.435 321.340 39.605 ;
        RECT 321.170 39.075 321.340 39.245 ;
        RECT 321.170 38.715 321.340 38.885 ;
        RECT 321.170 34.325 321.340 34.495 ;
        RECT 321.170 33.965 321.340 34.135 ;
        RECT 321.170 33.605 321.340 33.775 ;
        RECT 321.170 33.245 321.340 33.415 ;
        RECT 321.170 28.855 321.340 29.025 ;
        RECT 321.170 28.495 321.340 28.665 ;
        RECT 321.170 28.135 321.340 28.305 ;
        RECT 321.170 27.775 321.340 27.945 ;
        RECT 321.170 23.385 321.340 23.555 ;
        RECT 321.170 23.025 321.340 23.195 ;
        RECT 321.170 22.665 321.340 22.835 ;
        RECT 321.170 22.305 321.340 22.475 ;
        RECT 321.170 17.915 321.340 18.085 ;
        RECT 337.040 39.795 337.210 39.965 ;
        RECT 326.460 39.435 326.630 39.605 ;
        RECT 326.460 39.075 326.630 39.245 ;
        RECT 326.460 38.715 326.630 38.885 ;
        RECT 326.460 34.325 326.630 34.495 ;
        RECT 326.460 33.965 326.630 34.135 ;
        RECT 326.460 33.605 326.630 33.775 ;
        RECT 326.460 33.245 326.630 33.415 ;
        RECT 326.460 28.855 326.630 29.025 ;
        RECT 326.460 28.495 326.630 28.665 ;
        RECT 326.460 28.135 326.630 28.305 ;
        RECT 326.460 27.775 326.630 27.945 ;
        RECT 326.460 23.385 326.630 23.555 ;
        RECT 326.460 23.025 326.630 23.195 ;
        RECT 326.460 22.665 326.630 22.835 ;
        RECT 326.460 22.305 326.630 22.475 ;
        RECT 326.460 17.915 326.630 18.085 ;
        RECT 331.750 39.435 331.920 39.605 ;
        RECT 331.750 39.075 331.920 39.245 ;
        RECT 331.750 38.715 331.920 38.885 ;
        RECT 331.750 34.325 331.920 34.495 ;
        RECT 331.750 33.965 331.920 34.135 ;
        RECT 331.750 33.605 331.920 33.775 ;
        RECT 331.750 33.245 331.920 33.415 ;
        RECT 331.750 28.855 331.920 29.025 ;
        RECT 331.750 28.495 331.920 28.665 ;
        RECT 331.750 28.135 331.920 28.305 ;
        RECT 331.750 27.775 331.920 27.945 ;
        RECT 331.750 23.385 331.920 23.555 ;
        RECT 331.750 23.025 331.920 23.195 ;
        RECT 331.750 22.665 331.920 22.835 ;
        RECT 331.750 22.305 331.920 22.475 ;
        RECT 310.590 17.555 310.760 17.725 ;
        RECT 310.590 17.195 310.760 17.365 ;
        RECT 315.880 17.555 316.050 17.725 ;
        RECT 310.590 16.835 310.760 17.005 ;
        RECT 315.880 17.195 316.050 17.365 ;
        RECT 321.170 17.555 321.340 17.725 ;
        RECT 315.880 16.835 316.050 17.005 ;
        RECT 321.170 17.195 321.340 17.365 ;
        RECT 331.750 17.915 331.920 18.085 ;
        RECT 337.040 39.435 337.210 39.605 ;
        RECT 337.040 39.075 337.210 39.245 ;
        RECT 337.040 38.715 337.210 38.885 ;
        RECT 337.040 34.325 337.210 34.495 ;
        RECT 337.040 33.965 337.210 34.135 ;
        RECT 337.040 33.605 337.210 33.775 ;
        RECT 337.040 33.245 337.210 33.415 ;
        RECT 337.040 28.855 337.210 29.025 ;
        RECT 337.040 28.495 337.210 28.665 ;
        RECT 337.040 28.135 337.210 28.305 ;
        RECT 337.040 27.775 337.210 27.945 ;
        RECT 342.930 69.075 343.100 69.245 ;
        RECT 342.930 68.715 343.100 68.885 ;
        RECT 348.220 69.075 348.390 69.245 ;
        RECT 353.510 69.075 353.680 69.245 ;
        RECT 358.800 69.075 358.970 69.245 ;
        RECT 364.090 69.075 364.260 69.245 ;
        RECT 342.930 68.355 343.100 68.525 ;
        RECT 342.930 67.995 343.100 68.165 ;
        RECT 348.220 68.715 348.390 68.885 ;
        RECT 348.220 68.355 348.390 68.525 ;
        RECT 348.220 67.995 348.390 68.165 ;
        RECT 342.930 63.605 343.100 63.775 ;
        RECT 342.930 63.245 343.100 63.415 ;
        RECT 342.930 62.885 343.100 63.055 ;
        RECT 342.930 62.525 343.100 62.695 ;
        RECT 348.220 63.605 348.390 63.775 ;
        RECT 348.220 63.245 348.390 63.415 ;
        RECT 348.220 62.885 348.390 63.055 ;
        RECT 348.220 62.525 348.390 62.695 ;
        RECT 342.930 58.135 343.100 58.305 ;
        RECT 342.930 57.775 343.100 57.945 ;
        RECT 342.930 57.415 343.100 57.585 ;
        RECT 342.930 57.055 343.100 57.225 ;
        RECT 348.220 58.135 348.390 58.305 ;
        RECT 348.220 57.775 348.390 57.945 ;
        RECT 348.220 57.415 348.390 57.585 ;
        RECT 348.220 57.055 348.390 57.225 ;
        RECT 342.930 52.665 343.100 52.835 ;
        RECT 342.930 52.305 343.100 52.475 ;
        RECT 342.930 51.945 343.100 52.115 ;
        RECT 342.930 51.585 343.100 51.755 ;
        RECT 348.220 52.665 348.390 52.835 ;
        RECT 348.220 52.305 348.390 52.475 ;
        RECT 348.220 51.945 348.390 52.115 ;
        RECT 348.220 51.585 348.390 51.755 ;
        RECT 342.930 47.195 343.100 47.365 ;
        RECT 348.220 47.195 348.390 47.365 ;
        RECT 353.510 68.715 353.680 68.885 ;
        RECT 353.510 68.355 353.680 68.525 ;
        RECT 353.510 67.995 353.680 68.165 ;
        RECT 353.510 63.605 353.680 63.775 ;
        RECT 353.510 63.245 353.680 63.415 ;
        RECT 353.510 62.885 353.680 63.055 ;
        RECT 353.510 62.525 353.680 62.695 ;
        RECT 353.510 58.135 353.680 58.305 ;
        RECT 353.510 57.775 353.680 57.945 ;
        RECT 353.510 57.415 353.680 57.585 ;
        RECT 353.510 57.055 353.680 57.225 ;
        RECT 353.510 52.665 353.680 52.835 ;
        RECT 353.510 52.305 353.680 52.475 ;
        RECT 353.510 51.945 353.680 52.115 ;
        RECT 353.510 51.585 353.680 51.755 ;
        RECT 353.510 47.195 353.680 47.365 ;
        RECT 369.380 69.075 369.550 69.245 ;
        RECT 358.800 68.715 358.970 68.885 ;
        RECT 358.800 68.355 358.970 68.525 ;
        RECT 358.800 67.995 358.970 68.165 ;
        RECT 358.800 63.605 358.970 63.775 ;
        RECT 358.800 63.245 358.970 63.415 ;
        RECT 358.800 62.885 358.970 63.055 ;
        RECT 358.800 62.525 358.970 62.695 ;
        RECT 358.800 58.135 358.970 58.305 ;
        RECT 358.800 57.775 358.970 57.945 ;
        RECT 358.800 57.415 358.970 57.585 ;
        RECT 358.800 57.055 358.970 57.225 ;
        RECT 358.800 52.665 358.970 52.835 ;
        RECT 358.800 52.305 358.970 52.475 ;
        RECT 358.800 51.945 358.970 52.115 ;
        RECT 358.800 51.585 358.970 51.755 ;
        RECT 358.800 47.195 358.970 47.365 ;
        RECT 364.090 68.715 364.260 68.885 ;
        RECT 364.090 68.355 364.260 68.525 ;
        RECT 364.090 67.995 364.260 68.165 ;
        RECT 364.090 63.605 364.260 63.775 ;
        RECT 364.090 63.245 364.260 63.415 ;
        RECT 364.090 62.885 364.260 63.055 ;
        RECT 364.090 62.525 364.260 62.695 ;
        RECT 364.090 58.135 364.260 58.305 ;
        RECT 364.090 57.775 364.260 57.945 ;
        RECT 364.090 57.415 364.260 57.585 ;
        RECT 364.090 57.055 364.260 57.225 ;
        RECT 364.090 52.665 364.260 52.835 ;
        RECT 364.090 52.305 364.260 52.475 ;
        RECT 364.090 51.945 364.260 52.115 ;
        RECT 364.090 51.585 364.260 51.755 ;
        RECT 342.930 46.835 343.100 47.005 ;
        RECT 342.930 46.475 343.100 46.645 ;
        RECT 348.220 46.835 348.390 47.005 ;
        RECT 342.930 46.115 343.100 46.285 ;
        RECT 348.220 46.475 348.390 46.645 ;
        RECT 353.510 46.835 353.680 47.005 ;
        RECT 348.220 46.115 348.390 46.285 ;
        RECT 353.510 46.475 353.680 46.645 ;
        RECT 364.090 47.195 364.260 47.365 ;
        RECT 369.380 68.715 369.550 68.885 ;
        RECT 369.380 68.355 369.550 68.525 ;
        RECT 369.380 67.995 369.550 68.165 ;
        RECT 369.380 63.605 369.550 63.775 ;
        RECT 369.380 63.245 369.550 63.415 ;
        RECT 369.380 62.885 369.550 63.055 ;
        RECT 369.380 62.525 369.550 62.695 ;
        RECT 369.380 58.135 369.550 58.305 ;
        RECT 369.380 57.775 369.550 57.945 ;
        RECT 369.380 57.415 369.550 57.585 ;
        RECT 369.380 57.055 369.550 57.225 ;
        RECT 369.380 52.665 369.550 52.835 ;
        RECT 369.380 52.305 369.550 52.475 ;
        RECT 369.380 51.945 369.550 52.115 ;
        RECT 369.380 51.585 369.550 51.755 ;
        RECT 358.800 46.835 358.970 47.005 ;
        RECT 358.800 46.475 358.970 46.645 ;
        RECT 369.380 47.195 369.550 47.365 ;
        RECT 381.660 97.875 381.830 98.045 ;
        RECT 392.240 98.235 392.410 98.405 ;
        RECT 402.820 98.235 402.990 98.405 ;
        RECT 381.660 97.515 381.830 97.685 ;
        RECT 381.660 97.155 381.830 97.325 ;
        RECT 381.660 92.765 381.830 92.935 ;
        RECT 381.660 92.405 381.830 92.575 ;
        RECT 381.660 92.045 381.830 92.215 ;
        RECT 381.660 91.685 381.830 91.855 ;
        RECT 381.660 87.295 381.830 87.465 ;
        RECT 381.660 86.935 381.830 87.105 ;
        RECT 381.660 86.575 381.830 86.745 ;
        RECT 381.660 86.215 381.830 86.385 ;
        RECT 381.660 81.825 381.830 81.995 ;
        RECT 381.660 81.465 381.830 81.635 ;
        RECT 381.660 81.105 381.830 81.275 ;
        RECT 381.660 80.745 381.830 80.915 ;
        RECT 381.660 76.355 381.830 76.525 ;
        RECT 392.240 97.875 392.410 98.045 ;
        RECT 392.240 97.515 392.410 97.685 ;
        RECT 392.240 97.155 392.410 97.325 ;
        RECT 392.240 92.765 392.410 92.935 ;
        RECT 392.240 92.405 392.410 92.575 ;
        RECT 392.240 92.045 392.410 92.215 ;
        RECT 392.240 91.685 392.410 91.855 ;
        RECT 392.240 87.295 392.410 87.465 ;
        RECT 392.240 86.935 392.410 87.105 ;
        RECT 392.240 86.575 392.410 86.745 ;
        RECT 392.240 86.215 392.410 86.385 ;
        RECT 392.240 81.825 392.410 81.995 ;
        RECT 392.240 81.465 392.410 81.635 ;
        RECT 392.240 81.105 392.410 81.275 ;
        RECT 392.240 80.745 392.410 80.915 ;
        RECT 392.240 76.355 392.410 76.525 ;
        RECT 402.820 97.875 402.990 98.045 ;
        RECT 402.820 97.515 402.990 97.685 ;
        RECT 402.820 97.155 402.990 97.325 ;
        RECT 402.820 92.765 402.990 92.935 ;
        RECT 402.820 92.405 402.990 92.575 ;
        RECT 402.820 92.045 402.990 92.215 ;
        RECT 402.820 91.685 402.990 91.855 ;
        RECT 402.820 87.295 402.990 87.465 ;
        RECT 402.820 86.935 402.990 87.105 ;
        RECT 402.820 86.575 402.990 86.745 ;
        RECT 402.820 86.215 402.990 86.385 ;
        RECT 402.820 81.825 402.990 81.995 ;
        RECT 402.820 81.465 402.990 81.635 ;
        RECT 402.820 81.105 402.990 81.275 ;
        RECT 402.820 80.745 402.990 80.915 ;
        RECT 402.820 76.355 402.990 76.525 ;
        RECT 413.980 98.295 414.150 98.465 ;
        RECT 405.680 90.705 405.850 90.875 ;
        RECT 405.680 90.345 405.850 90.515 ;
        RECT 405.680 89.985 405.850 90.155 ;
        RECT 405.680 89.625 405.850 89.795 ;
        RECT 405.680 89.265 405.850 89.435 ;
        RECT 405.680 88.905 405.850 89.075 ;
        RECT 405.680 88.545 405.850 88.715 ;
        RECT 405.680 88.185 405.850 88.355 ;
        RECT 405.680 87.825 405.850 87.995 ;
        RECT 405.680 87.465 405.850 87.635 ;
        RECT 405.680 87.105 405.850 87.275 ;
        RECT 405.680 86.745 405.850 86.915 ;
        RECT 405.680 86.385 405.850 86.555 ;
        RECT 405.680 86.025 405.850 86.195 ;
        RECT 405.680 85.665 405.850 85.835 ;
        RECT 405.680 85.305 405.850 85.475 ;
        RECT 405.680 84.945 405.850 85.115 ;
        RECT 381.660 75.995 381.830 76.165 ;
        RECT 381.660 75.635 381.830 75.805 ;
        RECT 392.240 75.995 392.410 76.165 ;
        RECT 392.240 75.635 392.410 75.805 ;
        RECT 402.820 75.995 402.990 76.165 ;
        RECT 402.820 75.635 402.990 75.805 ;
        RECT 381.660 75.275 381.830 75.445 ;
        RECT 392.240 75.275 392.410 75.445 ;
        RECT 402.820 75.275 402.990 75.445 ;
        RECT 413.980 97.935 414.150 98.105 ;
        RECT 424.560 98.295 424.730 98.465 ;
        RECT 435.140 98.295 435.310 98.465 ;
        RECT 413.980 97.575 414.150 97.745 ;
        RECT 413.980 97.215 414.150 97.385 ;
        RECT 413.980 92.825 414.150 92.995 ;
        RECT 413.980 92.465 414.150 92.635 ;
        RECT 413.980 92.105 414.150 92.275 ;
        RECT 413.980 91.745 414.150 91.915 ;
        RECT 413.980 87.355 414.150 87.525 ;
        RECT 413.980 86.995 414.150 87.165 ;
        RECT 413.980 86.635 414.150 86.805 ;
        RECT 413.980 86.275 414.150 86.445 ;
        RECT 413.980 81.885 414.150 82.055 ;
        RECT 413.980 81.525 414.150 81.695 ;
        RECT 413.980 81.165 414.150 81.335 ;
        RECT 413.980 80.805 414.150 80.975 ;
        RECT 413.980 76.415 414.150 76.585 ;
        RECT 424.560 97.935 424.730 98.105 ;
        RECT 424.560 97.575 424.730 97.745 ;
        RECT 424.560 97.215 424.730 97.385 ;
        RECT 424.560 92.825 424.730 92.995 ;
        RECT 424.560 92.465 424.730 92.635 ;
        RECT 424.560 92.105 424.730 92.275 ;
        RECT 424.560 91.745 424.730 91.915 ;
        RECT 424.560 87.355 424.730 87.525 ;
        RECT 424.560 86.995 424.730 87.165 ;
        RECT 424.560 86.635 424.730 86.805 ;
        RECT 424.560 86.275 424.730 86.445 ;
        RECT 424.560 81.885 424.730 82.055 ;
        RECT 424.560 81.525 424.730 81.695 ;
        RECT 424.560 81.165 424.730 81.335 ;
        RECT 424.560 80.805 424.730 80.975 ;
        RECT 424.560 76.415 424.730 76.585 ;
        RECT 435.140 97.935 435.310 98.105 ;
        RECT 435.140 97.575 435.310 97.745 ;
        RECT 435.140 97.215 435.310 97.385 ;
        RECT 435.140 92.825 435.310 92.995 ;
        RECT 435.140 92.465 435.310 92.635 ;
        RECT 435.140 92.105 435.310 92.275 ;
        RECT 435.140 91.745 435.310 91.915 ;
        RECT 435.140 87.355 435.310 87.525 ;
        RECT 435.140 86.995 435.310 87.165 ;
        RECT 435.140 86.635 435.310 86.805 ;
        RECT 435.140 86.275 435.310 86.445 ;
        RECT 435.140 81.885 435.310 82.055 ;
        RECT 435.140 81.525 435.310 81.695 ;
        RECT 435.140 81.165 435.310 81.335 ;
        RECT 435.140 80.805 435.310 80.975 ;
        RECT 435.140 76.415 435.310 76.585 ;
        RECT 442.510 121.915 442.680 122.085 ;
        RECT 442.510 121.555 442.680 121.725 ;
        RECT 442.510 121.195 442.680 121.365 ;
        RECT 442.510 120.835 442.680 121.005 ;
        RECT 447.800 121.915 447.970 122.085 ;
        RECT 447.800 121.555 447.970 121.725 ;
        RECT 447.800 121.195 447.970 121.365 ;
        RECT 447.800 120.835 447.970 121.005 ;
        RECT 442.510 116.445 442.680 116.615 ;
        RECT 442.510 116.085 442.680 116.255 ;
        RECT 442.510 115.725 442.680 115.895 ;
        RECT 442.510 115.365 442.680 115.535 ;
        RECT 447.800 116.445 447.970 116.615 ;
        RECT 447.800 116.085 447.970 116.255 ;
        RECT 447.800 115.725 447.970 115.895 ;
        RECT 447.800 115.365 447.970 115.535 ;
        RECT 442.510 110.975 442.680 111.145 ;
        RECT 442.510 110.615 442.680 110.785 ;
        RECT 442.510 110.255 442.680 110.425 ;
        RECT 442.510 109.895 442.680 110.065 ;
        RECT 447.800 110.975 447.970 111.145 ;
        RECT 447.800 110.615 447.970 110.785 ;
        RECT 447.800 110.255 447.970 110.425 ;
        RECT 447.800 109.895 447.970 110.065 ;
        RECT 442.510 105.505 442.680 105.675 ;
        RECT 447.800 105.505 447.970 105.675 ;
        RECT 453.090 127.025 453.260 127.195 ;
        RECT 453.090 126.665 453.260 126.835 ;
        RECT 453.090 126.305 453.260 126.475 ;
        RECT 453.090 121.915 453.260 122.085 ;
        RECT 453.090 121.555 453.260 121.725 ;
        RECT 453.090 121.195 453.260 121.365 ;
        RECT 453.090 120.835 453.260 121.005 ;
        RECT 453.090 116.445 453.260 116.615 ;
        RECT 453.090 116.085 453.260 116.255 ;
        RECT 453.090 115.725 453.260 115.895 ;
        RECT 453.090 115.365 453.260 115.535 ;
        RECT 453.090 110.975 453.260 111.145 ;
        RECT 453.090 110.615 453.260 110.785 ;
        RECT 453.090 110.255 453.260 110.425 ;
        RECT 453.090 109.895 453.260 110.065 ;
        RECT 453.090 105.505 453.260 105.675 ;
        RECT 468.960 127.385 469.130 127.555 ;
        RECT 474.820 127.375 474.990 127.545 ;
        RECT 458.380 127.025 458.550 127.195 ;
        RECT 458.380 126.665 458.550 126.835 ;
        RECT 458.380 126.305 458.550 126.475 ;
        RECT 458.380 121.915 458.550 122.085 ;
        RECT 458.380 121.555 458.550 121.725 ;
        RECT 458.380 121.195 458.550 121.365 ;
        RECT 458.380 120.835 458.550 121.005 ;
        RECT 458.380 116.445 458.550 116.615 ;
        RECT 458.380 116.085 458.550 116.255 ;
        RECT 458.380 115.725 458.550 115.895 ;
        RECT 458.380 115.365 458.550 115.535 ;
        RECT 458.380 110.975 458.550 111.145 ;
        RECT 458.380 110.615 458.550 110.785 ;
        RECT 458.380 110.255 458.550 110.425 ;
        RECT 458.380 109.895 458.550 110.065 ;
        RECT 458.380 105.505 458.550 105.675 ;
        RECT 463.670 127.025 463.840 127.195 ;
        RECT 463.670 126.665 463.840 126.835 ;
        RECT 463.670 126.305 463.840 126.475 ;
        RECT 463.670 121.915 463.840 122.085 ;
        RECT 463.670 121.555 463.840 121.725 ;
        RECT 463.670 121.195 463.840 121.365 ;
        RECT 463.670 120.835 463.840 121.005 ;
        RECT 463.670 116.445 463.840 116.615 ;
        RECT 463.670 116.085 463.840 116.255 ;
        RECT 463.670 115.725 463.840 115.895 ;
        RECT 463.670 115.365 463.840 115.535 ;
        RECT 463.670 110.975 463.840 111.145 ;
        RECT 463.670 110.615 463.840 110.785 ;
        RECT 463.670 110.255 463.840 110.425 ;
        RECT 463.670 109.895 463.840 110.065 ;
        RECT 442.510 105.145 442.680 105.315 ;
        RECT 442.510 104.785 442.680 104.955 ;
        RECT 447.800 105.145 447.970 105.315 ;
        RECT 442.510 104.425 442.680 104.595 ;
        RECT 447.800 104.785 447.970 104.955 ;
        RECT 453.090 105.145 453.260 105.315 ;
        RECT 447.800 104.425 447.970 104.595 ;
        RECT 453.090 104.785 453.260 104.955 ;
        RECT 463.670 105.505 463.840 105.675 ;
        RECT 468.960 127.025 469.130 127.195 ;
        RECT 468.960 126.665 469.130 126.835 ;
        RECT 468.960 126.305 469.130 126.475 ;
        RECT 474.820 127.015 474.990 127.185 ;
        RECT 480.110 127.375 480.280 127.545 ;
        RECT 485.400 127.375 485.570 127.545 ;
        RECT 490.690 127.375 490.860 127.545 ;
        RECT 495.980 127.375 496.150 127.545 ;
        RECT 474.820 126.655 474.990 126.825 ;
        RECT 474.820 126.295 474.990 126.465 ;
        RECT 480.110 127.015 480.280 127.185 ;
        RECT 480.110 126.655 480.280 126.825 ;
        RECT 480.110 126.295 480.280 126.465 ;
        RECT 468.960 121.915 469.130 122.085 ;
        RECT 468.960 121.555 469.130 121.725 ;
        RECT 468.960 121.195 469.130 121.365 ;
        RECT 468.960 120.835 469.130 121.005 ;
        RECT 468.960 116.445 469.130 116.615 ;
        RECT 468.960 116.085 469.130 116.255 ;
        RECT 468.960 115.725 469.130 115.895 ;
        RECT 468.960 115.365 469.130 115.535 ;
        RECT 468.960 110.975 469.130 111.145 ;
        RECT 468.960 110.615 469.130 110.785 ;
        RECT 468.960 110.255 469.130 110.425 ;
        RECT 468.960 109.895 469.130 110.065 ;
        RECT 458.380 105.145 458.550 105.315 ;
        RECT 458.380 104.785 458.550 104.955 ;
        RECT 468.960 105.505 469.130 105.675 ;
        RECT 471.810 119.785 471.980 119.955 ;
        RECT 471.810 119.425 471.980 119.595 ;
        RECT 471.810 119.065 471.980 119.235 ;
        RECT 471.810 118.705 471.980 118.875 ;
        RECT 471.810 118.345 471.980 118.515 ;
        RECT 471.810 117.985 471.980 118.155 ;
        RECT 471.810 117.625 471.980 117.795 ;
        RECT 471.810 117.265 471.980 117.435 ;
        RECT 471.810 116.905 471.980 117.075 ;
        RECT 471.810 116.545 471.980 116.715 ;
        RECT 471.810 116.185 471.980 116.355 ;
        RECT 471.810 115.825 471.980 115.995 ;
        RECT 471.810 115.465 471.980 115.635 ;
        RECT 471.810 115.105 471.980 115.275 ;
        RECT 471.810 114.745 471.980 114.915 ;
        RECT 471.810 114.385 471.980 114.555 ;
        RECT 471.810 114.025 471.980 114.195 ;
        RECT 463.670 105.145 463.840 105.315 ;
        RECT 463.670 104.785 463.840 104.955 ;
        RECT 468.960 105.145 469.130 105.315 ;
        RECT 453.090 104.425 453.260 104.595 ;
        RECT 458.380 104.425 458.550 104.595 ;
        RECT 463.670 104.425 463.840 104.595 ;
        RECT 468.960 104.785 469.130 104.955 ;
        RECT 468.960 104.425 469.130 104.595 ;
        RECT 439.530 90.605 439.700 90.775 ;
        RECT 439.530 90.245 439.700 90.415 ;
        RECT 439.530 89.885 439.700 90.055 ;
        RECT 439.530 89.525 439.700 89.695 ;
        RECT 439.530 89.165 439.700 89.335 ;
        RECT 439.530 88.805 439.700 88.975 ;
        RECT 439.530 88.445 439.700 88.615 ;
        RECT 439.530 88.085 439.700 88.255 ;
        RECT 439.530 87.725 439.700 87.895 ;
        RECT 439.530 87.365 439.700 87.535 ;
        RECT 439.530 87.005 439.700 87.175 ;
        RECT 439.530 86.645 439.700 86.815 ;
        RECT 439.530 86.285 439.700 86.455 ;
        RECT 439.530 85.925 439.700 86.095 ;
        RECT 439.530 85.565 439.700 85.735 ;
        RECT 439.530 85.205 439.700 85.375 ;
        RECT 439.530 84.845 439.700 85.015 ;
        RECT 413.980 76.055 414.150 76.225 ;
        RECT 413.980 75.695 414.150 75.865 ;
        RECT 424.560 76.055 424.730 76.225 ;
        RECT 424.560 75.695 424.730 75.865 ;
        RECT 435.140 76.055 435.310 76.225 ;
        RECT 435.140 75.695 435.310 75.865 ;
        RECT 413.980 75.335 414.150 75.505 ;
        RECT 424.560 75.335 424.730 75.505 ;
        RECT 435.140 75.335 435.310 75.505 ;
        RECT 381.660 68.945 381.830 69.115 ;
        RECT 373.360 61.355 373.530 61.525 ;
        RECT 373.360 60.995 373.530 61.165 ;
        RECT 373.360 60.635 373.530 60.805 ;
        RECT 373.360 60.275 373.530 60.445 ;
        RECT 373.360 59.915 373.530 60.085 ;
        RECT 373.360 59.555 373.530 59.725 ;
        RECT 373.360 59.195 373.530 59.365 ;
        RECT 373.360 58.835 373.530 59.005 ;
        RECT 373.360 58.475 373.530 58.645 ;
        RECT 373.360 58.115 373.530 58.285 ;
        RECT 373.360 57.755 373.530 57.925 ;
        RECT 373.360 57.395 373.530 57.565 ;
        RECT 373.360 57.035 373.530 57.205 ;
        RECT 373.360 56.675 373.530 56.845 ;
        RECT 373.360 56.315 373.530 56.485 ;
        RECT 373.360 55.955 373.530 56.125 ;
        RECT 373.360 55.595 373.530 55.765 ;
        RECT 364.090 46.835 364.260 47.005 ;
        RECT 364.090 46.475 364.260 46.645 ;
        RECT 369.380 46.835 369.550 47.005 ;
        RECT 353.510 46.115 353.680 46.285 ;
        RECT 358.800 46.115 358.970 46.285 ;
        RECT 364.090 46.115 364.260 46.285 ;
        RECT 369.380 46.475 369.550 46.645 ;
        RECT 369.380 46.115 369.550 46.285 ;
        RECT 339.940 32.195 340.110 32.365 ;
        RECT 339.940 31.835 340.110 32.005 ;
        RECT 339.940 31.475 340.110 31.645 ;
        RECT 339.940 31.115 340.110 31.285 ;
        RECT 339.940 30.755 340.110 30.925 ;
        RECT 339.940 30.395 340.110 30.565 ;
        RECT 339.940 30.035 340.110 30.205 ;
        RECT 339.940 29.675 340.110 29.845 ;
        RECT 339.940 29.315 340.110 29.485 ;
        RECT 339.940 28.955 340.110 29.125 ;
        RECT 339.940 28.595 340.110 28.765 ;
        RECT 339.940 28.235 340.110 28.405 ;
        RECT 339.940 27.875 340.110 28.045 ;
        RECT 339.940 27.515 340.110 27.685 ;
        RECT 339.940 27.155 340.110 27.325 ;
        RECT 339.940 26.795 340.110 26.965 ;
        RECT 339.940 26.435 340.110 26.605 ;
        RECT 342.950 39.785 343.120 39.955 ;
        RECT 342.950 39.425 343.120 39.595 ;
        RECT 348.240 39.785 348.410 39.955 ;
        RECT 353.530 39.785 353.700 39.955 ;
        RECT 358.820 39.785 358.990 39.955 ;
        RECT 364.110 39.785 364.280 39.955 ;
        RECT 342.950 39.065 343.120 39.235 ;
        RECT 342.950 38.705 343.120 38.875 ;
        RECT 348.240 39.425 348.410 39.595 ;
        RECT 348.240 39.065 348.410 39.235 ;
        RECT 348.240 38.705 348.410 38.875 ;
        RECT 342.950 34.315 343.120 34.485 ;
        RECT 342.950 33.955 343.120 34.125 ;
        RECT 342.950 33.595 343.120 33.765 ;
        RECT 342.950 33.235 343.120 33.405 ;
        RECT 348.240 34.315 348.410 34.485 ;
        RECT 348.240 33.955 348.410 34.125 ;
        RECT 348.240 33.595 348.410 33.765 ;
        RECT 348.240 33.235 348.410 33.405 ;
        RECT 342.950 28.845 343.120 29.015 ;
        RECT 342.950 28.485 343.120 28.655 ;
        RECT 342.950 28.125 343.120 28.295 ;
        RECT 342.950 27.765 343.120 27.935 ;
        RECT 348.240 28.845 348.410 29.015 ;
        RECT 348.240 28.485 348.410 28.655 ;
        RECT 348.240 28.125 348.410 28.295 ;
        RECT 348.240 27.765 348.410 27.935 ;
        RECT 337.040 23.385 337.210 23.555 ;
        RECT 337.040 23.025 337.210 23.195 ;
        RECT 337.040 22.665 337.210 22.835 ;
        RECT 337.040 22.305 337.210 22.475 ;
        RECT 326.460 17.555 326.630 17.725 ;
        RECT 326.460 17.195 326.630 17.365 ;
        RECT 337.040 17.915 337.210 18.085 ;
        RECT 331.750 17.555 331.920 17.725 ;
        RECT 331.750 17.195 331.920 17.365 ;
        RECT 337.040 17.555 337.210 17.725 ;
        RECT 321.170 16.835 321.340 17.005 ;
        RECT 326.460 16.835 326.630 17.005 ;
        RECT 331.750 16.835 331.920 17.005 ;
        RECT 337.040 17.195 337.210 17.365 ;
        RECT 337.040 16.835 337.210 17.005 ;
        RECT 342.950 23.375 343.120 23.545 ;
        RECT 342.950 23.015 343.120 23.185 ;
        RECT 342.950 22.655 343.120 22.825 ;
        RECT 342.950 22.295 343.120 22.465 ;
        RECT 348.240 23.375 348.410 23.545 ;
        RECT 348.240 23.015 348.410 23.185 ;
        RECT 348.240 22.655 348.410 22.825 ;
        RECT 348.240 22.295 348.410 22.465 ;
        RECT 342.950 17.905 343.120 18.075 ;
        RECT 348.240 17.905 348.410 18.075 ;
        RECT 353.530 39.425 353.700 39.595 ;
        RECT 353.530 39.065 353.700 39.235 ;
        RECT 353.530 38.705 353.700 38.875 ;
        RECT 353.530 34.315 353.700 34.485 ;
        RECT 353.530 33.955 353.700 34.125 ;
        RECT 353.530 33.595 353.700 33.765 ;
        RECT 353.530 33.235 353.700 33.405 ;
        RECT 353.530 28.845 353.700 29.015 ;
        RECT 353.530 28.485 353.700 28.655 ;
        RECT 353.530 28.125 353.700 28.295 ;
        RECT 353.530 27.765 353.700 27.935 ;
        RECT 353.530 23.375 353.700 23.545 ;
        RECT 353.530 23.015 353.700 23.185 ;
        RECT 353.530 22.655 353.700 22.825 ;
        RECT 353.530 22.295 353.700 22.465 ;
        RECT 353.530 17.905 353.700 18.075 ;
        RECT 369.400 39.785 369.570 39.955 ;
        RECT 358.820 39.425 358.990 39.595 ;
        RECT 358.820 39.065 358.990 39.235 ;
        RECT 358.820 38.705 358.990 38.875 ;
        RECT 358.820 34.315 358.990 34.485 ;
        RECT 358.820 33.955 358.990 34.125 ;
        RECT 358.820 33.595 358.990 33.765 ;
        RECT 358.820 33.235 358.990 33.405 ;
        RECT 358.820 28.845 358.990 29.015 ;
        RECT 358.820 28.485 358.990 28.655 ;
        RECT 358.820 28.125 358.990 28.295 ;
        RECT 358.820 27.765 358.990 27.935 ;
        RECT 358.820 23.375 358.990 23.545 ;
        RECT 358.820 23.015 358.990 23.185 ;
        RECT 358.820 22.655 358.990 22.825 ;
        RECT 358.820 22.295 358.990 22.465 ;
        RECT 358.820 17.905 358.990 18.075 ;
        RECT 364.110 39.425 364.280 39.595 ;
        RECT 364.110 39.065 364.280 39.235 ;
        RECT 364.110 38.705 364.280 38.875 ;
        RECT 364.110 34.315 364.280 34.485 ;
        RECT 364.110 33.955 364.280 34.125 ;
        RECT 364.110 33.595 364.280 33.765 ;
        RECT 364.110 33.235 364.280 33.405 ;
        RECT 364.110 28.845 364.280 29.015 ;
        RECT 364.110 28.485 364.280 28.655 ;
        RECT 364.110 28.125 364.280 28.295 ;
        RECT 364.110 27.765 364.280 27.935 ;
        RECT 364.110 23.375 364.280 23.545 ;
        RECT 364.110 23.015 364.280 23.185 ;
        RECT 364.110 22.655 364.280 22.825 ;
        RECT 364.110 22.295 364.280 22.465 ;
        RECT 342.950 17.545 343.120 17.715 ;
        RECT 342.950 17.185 343.120 17.355 ;
        RECT 348.240 17.545 348.410 17.715 ;
        RECT 342.950 16.825 343.120 16.995 ;
        RECT 348.240 17.185 348.410 17.355 ;
        RECT 353.530 17.545 353.700 17.715 ;
        RECT 348.240 16.825 348.410 16.995 ;
        RECT 353.530 17.185 353.700 17.355 ;
        RECT 364.110 17.905 364.280 18.075 ;
        RECT 369.400 39.425 369.570 39.595 ;
        RECT 369.400 39.065 369.570 39.235 ;
        RECT 369.400 38.705 369.570 38.875 ;
        RECT 369.400 34.315 369.570 34.485 ;
        RECT 369.400 33.955 369.570 34.125 ;
        RECT 369.400 33.595 369.570 33.765 ;
        RECT 369.400 33.235 369.570 33.405 ;
        RECT 369.400 28.845 369.570 29.015 ;
        RECT 369.400 28.485 369.570 28.655 ;
        RECT 369.400 28.125 369.570 28.295 ;
        RECT 369.400 27.765 369.570 27.935 ;
        RECT 369.400 23.375 369.570 23.545 ;
        RECT 369.400 23.015 369.570 23.185 ;
        RECT 369.400 22.655 369.570 22.825 ;
        RECT 369.400 22.295 369.570 22.465 ;
        RECT 358.820 17.545 358.990 17.715 ;
        RECT 358.820 17.185 358.990 17.355 ;
        RECT 369.400 17.905 369.570 18.075 ;
        RECT 381.660 68.585 381.830 68.755 ;
        RECT 392.240 68.945 392.410 69.115 ;
        RECT 402.820 68.945 402.990 69.115 ;
        RECT 381.660 68.225 381.830 68.395 ;
        RECT 381.660 67.865 381.830 68.035 ;
        RECT 381.660 63.475 381.830 63.645 ;
        RECT 381.660 63.115 381.830 63.285 ;
        RECT 381.660 62.755 381.830 62.925 ;
        RECT 381.660 62.395 381.830 62.565 ;
        RECT 381.660 58.005 381.830 58.175 ;
        RECT 381.660 57.645 381.830 57.815 ;
        RECT 381.660 57.285 381.830 57.455 ;
        RECT 381.660 56.925 381.830 57.095 ;
        RECT 381.660 52.535 381.830 52.705 ;
        RECT 381.660 52.175 381.830 52.345 ;
        RECT 381.660 51.815 381.830 51.985 ;
        RECT 381.660 51.455 381.830 51.625 ;
        RECT 381.660 47.065 381.830 47.235 ;
        RECT 392.240 68.585 392.410 68.755 ;
        RECT 392.240 68.225 392.410 68.395 ;
        RECT 392.240 67.865 392.410 68.035 ;
        RECT 392.240 63.475 392.410 63.645 ;
        RECT 392.240 63.115 392.410 63.285 ;
        RECT 392.240 62.755 392.410 62.925 ;
        RECT 392.240 62.395 392.410 62.565 ;
        RECT 392.240 58.005 392.410 58.175 ;
        RECT 392.240 57.645 392.410 57.815 ;
        RECT 392.240 57.285 392.410 57.455 ;
        RECT 392.240 56.925 392.410 57.095 ;
        RECT 392.240 52.535 392.410 52.705 ;
        RECT 392.240 52.175 392.410 52.345 ;
        RECT 392.240 51.815 392.410 51.985 ;
        RECT 392.240 51.455 392.410 51.625 ;
        RECT 392.240 47.065 392.410 47.235 ;
        RECT 402.820 68.585 402.990 68.755 ;
        RECT 402.820 68.225 402.990 68.395 ;
        RECT 402.820 67.865 402.990 68.035 ;
        RECT 402.820 63.475 402.990 63.645 ;
        RECT 402.820 63.115 402.990 63.285 ;
        RECT 402.820 62.755 402.990 62.925 ;
        RECT 402.820 62.395 402.990 62.565 ;
        RECT 402.820 58.005 402.990 58.175 ;
        RECT 402.820 57.645 402.990 57.815 ;
        RECT 402.820 57.285 402.990 57.455 ;
        RECT 402.820 56.925 402.990 57.095 ;
        RECT 402.820 52.535 402.990 52.705 ;
        RECT 402.820 52.175 402.990 52.345 ;
        RECT 402.820 51.815 402.990 51.985 ;
        RECT 402.820 51.455 402.990 51.625 ;
        RECT 402.820 47.065 402.990 47.235 ;
        RECT 414.000 68.935 414.170 69.105 ;
        RECT 405.700 61.345 405.870 61.515 ;
        RECT 405.700 60.985 405.870 61.155 ;
        RECT 405.700 60.625 405.870 60.795 ;
        RECT 405.700 60.265 405.870 60.435 ;
        RECT 405.700 59.905 405.870 60.075 ;
        RECT 405.700 59.545 405.870 59.715 ;
        RECT 405.700 59.185 405.870 59.355 ;
        RECT 405.700 58.825 405.870 58.995 ;
        RECT 405.700 58.465 405.870 58.635 ;
        RECT 405.700 58.105 405.870 58.275 ;
        RECT 405.700 57.745 405.870 57.915 ;
        RECT 405.700 57.385 405.870 57.555 ;
        RECT 405.700 57.025 405.870 57.195 ;
        RECT 405.700 56.665 405.870 56.835 ;
        RECT 405.700 56.305 405.870 56.475 ;
        RECT 405.700 55.945 405.870 56.115 ;
        RECT 405.700 55.585 405.870 55.755 ;
        RECT 381.660 46.705 381.830 46.875 ;
        RECT 381.660 46.345 381.830 46.515 ;
        RECT 392.240 46.705 392.410 46.875 ;
        RECT 392.240 46.345 392.410 46.515 ;
        RECT 402.820 46.705 402.990 46.875 ;
        RECT 402.820 46.345 402.990 46.515 ;
        RECT 381.660 45.985 381.830 46.155 ;
        RECT 392.240 45.985 392.410 46.155 ;
        RECT 402.820 45.985 402.990 46.155 ;
        RECT 414.000 68.575 414.170 68.745 ;
        RECT 424.580 68.935 424.750 69.105 ;
        RECT 435.160 68.935 435.330 69.105 ;
        RECT 414.000 68.215 414.170 68.385 ;
        RECT 414.000 67.855 414.170 68.025 ;
        RECT 414.000 63.465 414.170 63.635 ;
        RECT 414.000 63.105 414.170 63.275 ;
        RECT 414.000 62.745 414.170 62.915 ;
        RECT 414.000 62.385 414.170 62.555 ;
        RECT 414.000 57.995 414.170 58.165 ;
        RECT 414.000 57.635 414.170 57.805 ;
        RECT 414.000 57.275 414.170 57.445 ;
        RECT 414.000 56.915 414.170 57.085 ;
        RECT 414.000 52.525 414.170 52.695 ;
        RECT 414.000 52.165 414.170 52.335 ;
        RECT 414.000 51.805 414.170 51.975 ;
        RECT 414.000 51.445 414.170 51.615 ;
        RECT 414.000 47.055 414.170 47.225 ;
        RECT 424.580 68.575 424.750 68.745 ;
        RECT 424.580 68.215 424.750 68.385 ;
        RECT 424.580 67.855 424.750 68.025 ;
        RECT 424.580 63.465 424.750 63.635 ;
        RECT 424.580 63.105 424.750 63.275 ;
        RECT 424.580 62.745 424.750 62.915 ;
        RECT 424.580 62.385 424.750 62.555 ;
        RECT 424.580 57.995 424.750 58.165 ;
        RECT 424.580 57.635 424.750 57.805 ;
        RECT 424.580 57.275 424.750 57.445 ;
        RECT 424.580 56.915 424.750 57.085 ;
        RECT 424.580 52.525 424.750 52.695 ;
        RECT 424.580 52.165 424.750 52.335 ;
        RECT 424.580 51.805 424.750 51.975 ;
        RECT 424.580 51.445 424.750 51.615 ;
        RECT 424.580 47.055 424.750 47.225 ;
        RECT 435.160 68.575 435.330 68.745 ;
        RECT 435.160 68.215 435.330 68.385 ;
        RECT 435.160 67.855 435.330 68.025 ;
        RECT 435.160 63.465 435.330 63.635 ;
        RECT 435.160 63.105 435.330 63.275 ;
        RECT 435.160 62.745 435.330 62.915 ;
        RECT 435.160 62.385 435.330 62.555 ;
        RECT 435.160 57.995 435.330 58.165 ;
        RECT 435.160 57.635 435.330 57.805 ;
        RECT 435.160 57.275 435.330 57.445 ;
        RECT 435.160 56.915 435.330 57.085 ;
        RECT 435.160 52.525 435.330 52.695 ;
        RECT 435.160 52.165 435.330 52.335 ;
        RECT 435.160 51.805 435.330 51.975 ;
        RECT 435.160 51.445 435.330 51.615 ;
        RECT 435.160 47.055 435.330 47.225 ;
        RECT 442.540 98.195 442.710 98.365 ;
        RECT 442.540 97.835 442.710 98.005 ;
        RECT 447.830 98.195 448.000 98.365 ;
        RECT 453.120 98.195 453.290 98.365 ;
        RECT 458.410 98.195 458.580 98.365 ;
        RECT 463.700 98.195 463.870 98.365 ;
        RECT 442.540 97.475 442.710 97.645 ;
        RECT 442.540 97.115 442.710 97.285 ;
        RECT 447.830 97.835 448.000 98.005 ;
        RECT 447.830 97.475 448.000 97.645 ;
        RECT 447.830 97.115 448.000 97.285 ;
        RECT 442.540 92.725 442.710 92.895 ;
        RECT 442.540 92.365 442.710 92.535 ;
        RECT 442.540 92.005 442.710 92.175 ;
        RECT 442.540 91.645 442.710 91.815 ;
        RECT 447.830 92.725 448.000 92.895 ;
        RECT 447.830 92.365 448.000 92.535 ;
        RECT 447.830 92.005 448.000 92.175 ;
        RECT 447.830 91.645 448.000 91.815 ;
        RECT 442.540 87.255 442.710 87.425 ;
        RECT 442.540 86.895 442.710 87.065 ;
        RECT 442.540 86.535 442.710 86.705 ;
        RECT 442.540 86.175 442.710 86.345 ;
        RECT 447.830 87.255 448.000 87.425 ;
        RECT 447.830 86.895 448.000 87.065 ;
        RECT 447.830 86.535 448.000 86.705 ;
        RECT 447.830 86.175 448.000 86.345 ;
        RECT 442.540 81.785 442.710 81.955 ;
        RECT 442.540 81.425 442.710 81.595 ;
        RECT 442.540 81.065 442.710 81.235 ;
        RECT 442.540 80.705 442.710 80.875 ;
        RECT 447.830 81.785 448.000 81.955 ;
        RECT 447.830 81.425 448.000 81.595 ;
        RECT 447.830 81.065 448.000 81.235 ;
        RECT 447.830 80.705 448.000 80.875 ;
        RECT 442.540 76.315 442.710 76.485 ;
        RECT 447.830 76.315 448.000 76.485 ;
        RECT 453.120 97.835 453.290 98.005 ;
        RECT 453.120 97.475 453.290 97.645 ;
        RECT 453.120 97.115 453.290 97.285 ;
        RECT 453.120 92.725 453.290 92.895 ;
        RECT 453.120 92.365 453.290 92.535 ;
        RECT 453.120 92.005 453.290 92.175 ;
        RECT 453.120 91.645 453.290 91.815 ;
        RECT 453.120 87.255 453.290 87.425 ;
        RECT 453.120 86.895 453.290 87.065 ;
        RECT 453.120 86.535 453.290 86.705 ;
        RECT 453.120 86.175 453.290 86.345 ;
        RECT 453.120 81.785 453.290 81.955 ;
        RECT 453.120 81.425 453.290 81.595 ;
        RECT 453.120 81.065 453.290 81.235 ;
        RECT 453.120 80.705 453.290 80.875 ;
        RECT 453.120 76.315 453.290 76.485 ;
        RECT 468.990 98.195 469.160 98.365 ;
        RECT 458.410 97.835 458.580 98.005 ;
        RECT 458.410 97.475 458.580 97.645 ;
        RECT 458.410 97.115 458.580 97.285 ;
        RECT 458.410 92.725 458.580 92.895 ;
        RECT 458.410 92.365 458.580 92.535 ;
        RECT 458.410 92.005 458.580 92.175 ;
        RECT 458.410 91.645 458.580 91.815 ;
        RECT 458.410 87.255 458.580 87.425 ;
        RECT 458.410 86.895 458.580 87.065 ;
        RECT 458.410 86.535 458.580 86.705 ;
        RECT 458.410 86.175 458.580 86.345 ;
        RECT 458.410 81.785 458.580 81.955 ;
        RECT 458.410 81.425 458.580 81.595 ;
        RECT 458.410 81.065 458.580 81.235 ;
        RECT 458.410 80.705 458.580 80.875 ;
        RECT 458.410 76.315 458.580 76.485 ;
        RECT 463.700 97.835 463.870 98.005 ;
        RECT 463.700 97.475 463.870 97.645 ;
        RECT 463.700 97.115 463.870 97.285 ;
        RECT 463.700 92.725 463.870 92.895 ;
        RECT 463.700 92.365 463.870 92.535 ;
        RECT 463.700 92.005 463.870 92.175 ;
        RECT 463.700 91.645 463.870 91.815 ;
        RECT 463.700 87.255 463.870 87.425 ;
        RECT 463.700 86.895 463.870 87.065 ;
        RECT 463.700 86.535 463.870 86.705 ;
        RECT 463.700 86.175 463.870 86.345 ;
        RECT 463.700 81.785 463.870 81.955 ;
        RECT 463.700 81.425 463.870 81.595 ;
        RECT 463.700 81.065 463.870 81.235 ;
        RECT 463.700 80.705 463.870 80.875 ;
        RECT 442.540 75.955 442.710 76.125 ;
        RECT 442.540 75.595 442.710 75.765 ;
        RECT 447.830 75.955 448.000 76.125 ;
        RECT 442.540 75.235 442.710 75.405 ;
        RECT 447.830 75.595 448.000 75.765 ;
        RECT 453.120 75.955 453.290 76.125 ;
        RECT 447.830 75.235 448.000 75.405 ;
        RECT 453.120 75.595 453.290 75.765 ;
        RECT 463.700 76.315 463.870 76.485 ;
        RECT 468.990 97.835 469.160 98.005 ;
        RECT 468.990 97.475 469.160 97.645 ;
        RECT 468.990 97.115 469.160 97.285 ;
        RECT 468.990 92.725 469.160 92.895 ;
        RECT 468.990 92.365 469.160 92.535 ;
        RECT 468.990 92.005 469.160 92.175 ;
        RECT 468.990 91.645 469.160 91.815 ;
        RECT 468.990 87.255 469.160 87.425 ;
        RECT 468.990 86.895 469.160 87.065 ;
        RECT 468.990 86.535 469.160 86.705 ;
        RECT 468.990 86.175 469.160 86.345 ;
        RECT 468.990 81.785 469.160 81.955 ;
        RECT 468.990 81.425 469.160 81.595 ;
        RECT 468.990 81.065 469.160 81.235 ;
        RECT 468.990 80.705 469.160 80.875 ;
        RECT 458.410 75.955 458.580 76.125 ;
        RECT 458.410 75.595 458.580 75.765 ;
        RECT 468.990 76.315 469.160 76.485 ;
        RECT 474.820 121.905 474.990 122.075 ;
        RECT 474.820 121.545 474.990 121.715 ;
        RECT 474.820 121.185 474.990 121.355 ;
        RECT 474.820 120.825 474.990 120.995 ;
        RECT 480.110 121.905 480.280 122.075 ;
        RECT 480.110 121.545 480.280 121.715 ;
        RECT 480.110 121.185 480.280 121.355 ;
        RECT 480.110 120.825 480.280 120.995 ;
        RECT 474.820 116.435 474.990 116.605 ;
        RECT 474.820 116.075 474.990 116.245 ;
        RECT 474.820 115.715 474.990 115.885 ;
        RECT 474.820 115.355 474.990 115.525 ;
        RECT 480.110 116.435 480.280 116.605 ;
        RECT 480.110 116.075 480.280 116.245 ;
        RECT 480.110 115.715 480.280 115.885 ;
        RECT 480.110 115.355 480.280 115.525 ;
        RECT 474.820 110.965 474.990 111.135 ;
        RECT 474.820 110.605 474.990 110.775 ;
        RECT 474.820 110.245 474.990 110.415 ;
        RECT 474.820 109.885 474.990 110.055 ;
        RECT 480.110 110.965 480.280 111.135 ;
        RECT 480.110 110.605 480.280 110.775 ;
        RECT 480.110 110.245 480.280 110.415 ;
        RECT 480.110 109.885 480.280 110.055 ;
        RECT 474.820 105.495 474.990 105.665 ;
        RECT 480.110 105.495 480.280 105.665 ;
        RECT 485.400 127.015 485.570 127.185 ;
        RECT 485.400 126.655 485.570 126.825 ;
        RECT 485.400 126.295 485.570 126.465 ;
        RECT 485.400 121.905 485.570 122.075 ;
        RECT 485.400 121.545 485.570 121.715 ;
        RECT 485.400 121.185 485.570 121.355 ;
        RECT 485.400 120.825 485.570 120.995 ;
        RECT 485.400 116.435 485.570 116.605 ;
        RECT 485.400 116.075 485.570 116.245 ;
        RECT 485.400 115.715 485.570 115.885 ;
        RECT 485.400 115.355 485.570 115.525 ;
        RECT 485.400 110.965 485.570 111.135 ;
        RECT 485.400 110.605 485.570 110.775 ;
        RECT 485.400 110.245 485.570 110.415 ;
        RECT 485.400 109.885 485.570 110.055 ;
        RECT 485.400 105.495 485.570 105.665 ;
        RECT 501.270 127.375 501.440 127.545 ;
        RECT 490.690 127.015 490.860 127.185 ;
        RECT 490.690 126.655 490.860 126.825 ;
        RECT 490.690 126.295 490.860 126.465 ;
        RECT 490.690 121.905 490.860 122.075 ;
        RECT 490.690 121.545 490.860 121.715 ;
        RECT 490.690 121.185 490.860 121.355 ;
        RECT 490.690 120.825 490.860 120.995 ;
        RECT 490.690 116.435 490.860 116.605 ;
        RECT 490.690 116.075 490.860 116.245 ;
        RECT 490.690 115.715 490.860 115.885 ;
        RECT 490.690 115.355 490.860 115.525 ;
        RECT 490.690 110.965 490.860 111.135 ;
        RECT 490.690 110.605 490.860 110.775 ;
        RECT 490.690 110.245 490.860 110.415 ;
        RECT 490.690 109.885 490.860 110.055 ;
        RECT 490.690 105.495 490.860 105.665 ;
        RECT 495.980 127.015 496.150 127.185 ;
        RECT 501.270 127.015 501.440 127.185 ;
        RECT 495.980 126.655 496.150 126.825 ;
        RECT 495.980 126.295 496.150 126.465 ;
        RECT 495.980 121.905 496.150 122.075 ;
        RECT 495.980 121.545 496.150 121.715 ;
        RECT 495.980 121.185 496.150 121.355 ;
        RECT 495.980 120.825 496.150 120.995 ;
        RECT 495.980 116.435 496.150 116.605 ;
        RECT 495.980 116.075 496.150 116.245 ;
        RECT 495.980 115.715 496.150 115.885 ;
        RECT 495.980 115.355 496.150 115.525 ;
        RECT 495.980 110.965 496.150 111.135 ;
        RECT 495.980 110.605 496.150 110.775 ;
        RECT 495.980 110.245 496.150 110.415 ;
        RECT 495.980 109.885 496.150 110.055 ;
        RECT 474.820 105.135 474.990 105.305 ;
        RECT 474.820 104.775 474.990 104.945 ;
        RECT 480.110 105.135 480.280 105.305 ;
        RECT 474.820 104.415 474.990 104.585 ;
        RECT 480.110 104.775 480.280 104.945 ;
        RECT 485.400 105.135 485.570 105.305 ;
        RECT 480.110 104.415 480.280 104.585 ;
        RECT 485.400 104.775 485.570 104.945 ;
        RECT 495.980 105.495 496.150 105.665 ;
        RECT 501.270 126.655 501.440 126.825 ;
        RECT 501.270 126.295 501.440 126.465 ;
        RECT 501.270 121.905 501.440 122.075 ;
        RECT 501.270 121.545 501.440 121.715 ;
        RECT 501.270 121.185 501.440 121.355 ;
        RECT 501.270 120.825 501.440 120.995 ;
        RECT 501.270 116.435 501.440 116.605 ;
        RECT 501.270 116.075 501.440 116.245 ;
        RECT 501.270 115.715 501.440 115.885 ;
        RECT 501.270 115.355 501.440 115.525 ;
        RECT 501.270 110.965 501.440 111.135 ;
        RECT 501.270 110.605 501.440 110.775 ;
        RECT 501.270 110.245 501.440 110.415 ;
        RECT 501.270 109.885 501.440 110.055 ;
        RECT 490.690 105.135 490.860 105.305 ;
        RECT 490.690 104.775 490.860 104.945 ;
        RECT 501.270 105.495 501.440 105.665 ;
        RECT 503.990 108.975 506.320 124.985 ;
        RECT 495.980 105.135 496.150 105.305 ;
        RECT 495.980 104.775 496.150 104.945 ;
        RECT 501.270 105.135 501.440 105.305 ;
        RECT 485.400 104.415 485.570 104.585 ;
        RECT 490.690 104.415 490.860 104.585 ;
        RECT 495.980 104.415 496.150 104.585 ;
        RECT 501.270 104.775 501.440 104.945 ;
        RECT 501.270 104.415 501.440 104.585 ;
        RECT 471.850 90.665 472.020 90.835 ;
        RECT 471.850 90.305 472.020 90.475 ;
        RECT 471.850 89.945 472.020 90.115 ;
        RECT 471.850 89.585 472.020 89.755 ;
        RECT 471.850 89.225 472.020 89.395 ;
        RECT 471.850 88.865 472.020 89.035 ;
        RECT 471.850 88.505 472.020 88.675 ;
        RECT 471.850 88.145 472.020 88.315 ;
        RECT 471.850 87.785 472.020 87.955 ;
        RECT 471.850 87.425 472.020 87.595 ;
        RECT 471.850 87.065 472.020 87.235 ;
        RECT 471.850 86.705 472.020 86.875 ;
        RECT 471.850 86.345 472.020 86.515 ;
        RECT 471.850 85.985 472.020 86.155 ;
        RECT 471.850 85.625 472.020 85.795 ;
        RECT 471.850 85.265 472.020 85.435 ;
        RECT 471.850 84.905 472.020 85.075 ;
        RECT 463.700 75.955 463.870 76.125 ;
        RECT 463.700 75.595 463.870 75.765 ;
        RECT 468.990 75.955 469.160 76.125 ;
        RECT 453.120 75.235 453.290 75.405 ;
        RECT 458.410 75.235 458.580 75.405 ;
        RECT 463.700 75.235 463.870 75.405 ;
        RECT 468.990 75.595 469.160 75.765 ;
        RECT 468.990 75.235 469.160 75.405 ;
        RECT 439.530 61.315 439.700 61.485 ;
        RECT 439.530 60.955 439.700 61.125 ;
        RECT 439.530 60.595 439.700 60.765 ;
        RECT 439.530 60.235 439.700 60.405 ;
        RECT 439.530 59.875 439.700 60.045 ;
        RECT 439.530 59.515 439.700 59.685 ;
        RECT 439.530 59.155 439.700 59.325 ;
        RECT 439.530 58.795 439.700 58.965 ;
        RECT 439.530 58.435 439.700 58.605 ;
        RECT 439.530 58.075 439.700 58.245 ;
        RECT 439.530 57.715 439.700 57.885 ;
        RECT 439.530 57.355 439.700 57.525 ;
        RECT 439.530 56.995 439.700 57.165 ;
        RECT 439.530 56.635 439.700 56.805 ;
        RECT 439.530 56.275 439.700 56.445 ;
        RECT 439.530 55.915 439.700 56.085 ;
        RECT 439.530 55.555 439.700 55.725 ;
        RECT 414.000 46.695 414.170 46.865 ;
        RECT 414.000 46.335 414.170 46.505 ;
        RECT 424.580 46.695 424.750 46.865 ;
        RECT 424.580 46.335 424.750 46.505 ;
        RECT 435.160 46.695 435.330 46.865 ;
        RECT 435.160 46.335 435.330 46.505 ;
        RECT 414.000 45.975 414.170 46.145 ;
        RECT 424.580 45.975 424.750 46.145 ;
        RECT 435.160 45.975 435.330 46.145 ;
        RECT 381.660 39.655 381.830 39.825 ;
        RECT 373.360 32.065 373.530 32.235 ;
        RECT 373.360 31.705 373.530 31.875 ;
        RECT 373.360 31.345 373.530 31.515 ;
        RECT 373.360 30.985 373.530 31.155 ;
        RECT 373.360 30.625 373.530 30.795 ;
        RECT 373.360 30.265 373.530 30.435 ;
        RECT 373.360 29.905 373.530 30.075 ;
        RECT 373.360 29.545 373.530 29.715 ;
        RECT 373.360 29.185 373.530 29.355 ;
        RECT 373.360 28.825 373.530 28.995 ;
        RECT 373.360 28.465 373.530 28.635 ;
        RECT 373.360 28.105 373.530 28.275 ;
        RECT 373.360 27.745 373.530 27.915 ;
        RECT 373.360 27.385 373.530 27.555 ;
        RECT 373.360 27.025 373.530 27.195 ;
        RECT 373.360 26.665 373.530 26.835 ;
        RECT 373.360 26.305 373.530 26.475 ;
        RECT 364.110 17.545 364.280 17.715 ;
        RECT 364.110 17.185 364.280 17.355 ;
        RECT 369.400 17.545 369.570 17.715 ;
        RECT 353.530 16.825 353.700 16.995 ;
        RECT 358.820 16.825 358.990 16.995 ;
        RECT 364.110 16.825 364.280 16.995 ;
        RECT 369.400 17.185 369.570 17.355 ;
        RECT 381.660 39.295 381.830 39.465 ;
        RECT 392.240 39.655 392.410 39.825 ;
        RECT 402.820 39.655 402.990 39.825 ;
        RECT 381.660 38.935 381.830 39.105 ;
        RECT 381.660 38.575 381.830 38.745 ;
        RECT 381.660 34.185 381.830 34.355 ;
        RECT 381.660 33.825 381.830 33.995 ;
        RECT 381.660 33.465 381.830 33.635 ;
        RECT 381.660 33.105 381.830 33.275 ;
        RECT 381.660 28.715 381.830 28.885 ;
        RECT 381.660 28.355 381.830 28.525 ;
        RECT 381.660 27.995 381.830 28.165 ;
        RECT 381.660 27.635 381.830 27.805 ;
        RECT 381.660 23.245 381.830 23.415 ;
        RECT 381.660 22.885 381.830 23.055 ;
        RECT 381.660 22.525 381.830 22.695 ;
        RECT 381.660 22.165 381.830 22.335 ;
        RECT 381.660 17.775 381.830 17.945 ;
        RECT 392.240 39.295 392.410 39.465 ;
        RECT 392.240 38.935 392.410 39.105 ;
        RECT 392.240 38.575 392.410 38.745 ;
        RECT 392.240 34.185 392.410 34.355 ;
        RECT 392.240 33.825 392.410 33.995 ;
        RECT 392.240 33.465 392.410 33.635 ;
        RECT 392.240 33.105 392.410 33.275 ;
        RECT 392.240 28.715 392.410 28.885 ;
        RECT 392.240 28.355 392.410 28.525 ;
        RECT 392.240 27.995 392.410 28.165 ;
        RECT 392.240 27.635 392.410 27.805 ;
        RECT 392.240 23.245 392.410 23.415 ;
        RECT 392.240 22.885 392.410 23.055 ;
        RECT 392.240 22.525 392.410 22.695 ;
        RECT 392.240 22.165 392.410 22.335 ;
        RECT 392.240 17.775 392.410 17.945 ;
        RECT 402.820 39.295 402.990 39.465 ;
        RECT 402.820 38.935 402.990 39.105 ;
        RECT 402.820 38.575 402.990 38.745 ;
        RECT 402.820 34.185 402.990 34.355 ;
        RECT 402.820 33.825 402.990 33.995 ;
        RECT 402.820 33.465 402.990 33.635 ;
        RECT 402.820 33.105 402.990 33.275 ;
        RECT 402.820 28.715 402.990 28.885 ;
        RECT 402.820 28.355 402.990 28.525 ;
        RECT 402.820 27.995 402.990 28.165 ;
        RECT 402.820 27.635 402.990 27.805 ;
        RECT 402.820 23.245 402.990 23.415 ;
        RECT 402.820 22.885 402.990 23.055 ;
        RECT 402.820 22.525 402.990 22.695 ;
        RECT 402.820 22.165 402.990 22.335 ;
        RECT 402.820 17.775 402.990 17.945 ;
        RECT 414.020 39.645 414.190 39.815 ;
        RECT 405.720 32.055 405.890 32.225 ;
        RECT 405.720 31.695 405.890 31.865 ;
        RECT 405.720 31.335 405.890 31.505 ;
        RECT 405.720 30.975 405.890 31.145 ;
        RECT 405.720 30.615 405.890 30.785 ;
        RECT 405.720 30.255 405.890 30.425 ;
        RECT 405.720 29.895 405.890 30.065 ;
        RECT 405.720 29.535 405.890 29.705 ;
        RECT 405.720 29.175 405.890 29.345 ;
        RECT 405.720 28.815 405.890 28.985 ;
        RECT 405.720 28.455 405.890 28.625 ;
        RECT 405.720 28.095 405.890 28.265 ;
        RECT 405.720 27.735 405.890 27.905 ;
        RECT 405.720 27.375 405.890 27.545 ;
        RECT 405.720 27.015 405.890 27.185 ;
        RECT 405.720 26.655 405.890 26.825 ;
        RECT 405.720 26.295 405.890 26.465 ;
        RECT 381.660 17.415 381.830 17.585 ;
        RECT 369.400 16.825 369.570 16.995 ;
        RECT 335.530 -0.805 346.140 4.045 ;
        RECT 381.660 17.055 381.830 17.225 ;
        RECT 392.240 17.415 392.410 17.585 ;
        RECT 392.240 17.055 392.410 17.225 ;
        RECT 402.820 17.415 402.990 17.585 ;
        RECT 414.020 39.285 414.190 39.455 ;
        RECT 424.600 39.645 424.770 39.815 ;
        RECT 435.180 39.645 435.350 39.815 ;
        RECT 414.020 38.925 414.190 39.095 ;
        RECT 414.020 38.565 414.190 38.735 ;
        RECT 414.020 34.175 414.190 34.345 ;
        RECT 414.020 33.815 414.190 33.985 ;
        RECT 414.020 33.455 414.190 33.625 ;
        RECT 414.020 33.095 414.190 33.265 ;
        RECT 414.020 28.705 414.190 28.875 ;
        RECT 414.020 28.345 414.190 28.515 ;
        RECT 414.020 27.985 414.190 28.155 ;
        RECT 414.020 27.625 414.190 27.795 ;
        RECT 414.020 23.235 414.190 23.405 ;
        RECT 414.020 22.875 414.190 23.045 ;
        RECT 414.020 22.515 414.190 22.685 ;
        RECT 414.020 22.155 414.190 22.325 ;
        RECT 414.020 17.765 414.190 17.935 ;
        RECT 424.600 39.285 424.770 39.455 ;
        RECT 424.600 38.925 424.770 39.095 ;
        RECT 424.600 38.565 424.770 38.735 ;
        RECT 424.600 34.175 424.770 34.345 ;
        RECT 424.600 33.815 424.770 33.985 ;
        RECT 424.600 33.455 424.770 33.625 ;
        RECT 424.600 33.095 424.770 33.265 ;
        RECT 424.600 28.705 424.770 28.875 ;
        RECT 424.600 28.345 424.770 28.515 ;
        RECT 424.600 27.985 424.770 28.155 ;
        RECT 424.600 27.625 424.770 27.795 ;
        RECT 424.600 23.235 424.770 23.405 ;
        RECT 424.600 22.875 424.770 23.045 ;
        RECT 424.600 22.515 424.770 22.685 ;
        RECT 424.600 22.155 424.770 22.325 ;
        RECT 424.600 17.765 424.770 17.935 ;
        RECT 435.180 39.285 435.350 39.455 ;
        RECT 435.180 38.925 435.350 39.095 ;
        RECT 435.180 38.565 435.350 38.735 ;
        RECT 435.180 34.175 435.350 34.345 ;
        RECT 435.180 33.815 435.350 33.985 ;
        RECT 435.180 33.455 435.350 33.625 ;
        RECT 435.180 33.095 435.350 33.265 ;
        RECT 435.180 28.705 435.350 28.875 ;
        RECT 435.180 28.345 435.350 28.515 ;
        RECT 435.180 27.985 435.350 28.155 ;
        RECT 435.180 27.625 435.350 27.795 ;
        RECT 435.180 23.235 435.350 23.405 ;
        RECT 435.180 22.875 435.350 23.045 ;
        RECT 435.180 22.515 435.350 22.685 ;
        RECT 435.180 22.155 435.350 22.325 ;
        RECT 435.180 17.765 435.350 17.935 ;
        RECT 442.540 68.905 442.710 69.075 ;
        RECT 442.540 68.545 442.710 68.715 ;
        RECT 447.830 68.905 448.000 69.075 ;
        RECT 453.120 68.905 453.290 69.075 ;
        RECT 458.410 68.905 458.580 69.075 ;
        RECT 463.700 68.905 463.870 69.075 ;
        RECT 442.540 68.185 442.710 68.355 ;
        RECT 442.540 67.825 442.710 67.995 ;
        RECT 447.830 68.545 448.000 68.715 ;
        RECT 447.830 68.185 448.000 68.355 ;
        RECT 447.830 67.825 448.000 67.995 ;
        RECT 442.540 63.435 442.710 63.605 ;
        RECT 442.540 63.075 442.710 63.245 ;
        RECT 442.540 62.715 442.710 62.885 ;
        RECT 442.540 62.355 442.710 62.525 ;
        RECT 447.830 63.435 448.000 63.605 ;
        RECT 447.830 63.075 448.000 63.245 ;
        RECT 447.830 62.715 448.000 62.885 ;
        RECT 447.830 62.355 448.000 62.525 ;
        RECT 442.540 57.965 442.710 58.135 ;
        RECT 442.540 57.605 442.710 57.775 ;
        RECT 442.540 57.245 442.710 57.415 ;
        RECT 442.540 56.885 442.710 57.055 ;
        RECT 447.830 57.965 448.000 58.135 ;
        RECT 447.830 57.605 448.000 57.775 ;
        RECT 447.830 57.245 448.000 57.415 ;
        RECT 447.830 56.885 448.000 57.055 ;
        RECT 442.540 52.495 442.710 52.665 ;
        RECT 442.540 52.135 442.710 52.305 ;
        RECT 442.540 51.775 442.710 51.945 ;
        RECT 442.540 51.415 442.710 51.585 ;
        RECT 447.830 52.495 448.000 52.665 ;
        RECT 447.830 52.135 448.000 52.305 ;
        RECT 447.830 51.775 448.000 51.945 ;
        RECT 447.830 51.415 448.000 51.585 ;
        RECT 442.540 47.025 442.710 47.195 ;
        RECT 447.830 47.025 448.000 47.195 ;
        RECT 453.120 68.545 453.290 68.715 ;
        RECT 453.120 68.185 453.290 68.355 ;
        RECT 453.120 67.825 453.290 67.995 ;
        RECT 453.120 63.435 453.290 63.605 ;
        RECT 453.120 63.075 453.290 63.245 ;
        RECT 453.120 62.715 453.290 62.885 ;
        RECT 453.120 62.355 453.290 62.525 ;
        RECT 453.120 57.965 453.290 58.135 ;
        RECT 453.120 57.605 453.290 57.775 ;
        RECT 453.120 57.245 453.290 57.415 ;
        RECT 453.120 56.885 453.290 57.055 ;
        RECT 453.120 52.495 453.290 52.665 ;
        RECT 453.120 52.135 453.290 52.305 ;
        RECT 453.120 51.775 453.290 51.945 ;
        RECT 453.120 51.415 453.290 51.585 ;
        RECT 453.120 47.025 453.290 47.195 ;
        RECT 468.990 68.905 469.160 69.075 ;
        RECT 458.410 68.545 458.580 68.715 ;
        RECT 458.410 68.185 458.580 68.355 ;
        RECT 458.410 67.825 458.580 67.995 ;
        RECT 458.410 63.435 458.580 63.605 ;
        RECT 458.410 63.075 458.580 63.245 ;
        RECT 458.410 62.715 458.580 62.885 ;
        RECT 458.410 62.355 458.580 62.525 ;
        RECT 458.410 57.965 458.580 58.135 ;
        RECT 458.410 57.605 458.580 57.775 ;
        RECT 458.410 57.245 458.580 57.415 ;
        RECT 458.410 56.885 458.580 57.055 ;
        RECT 458.410 52.495 458.580 52.665 ;
        RECT 458.410 52.135 458.580 52.305 ;
        RECT 458.410 51.775 458.580 51.945 ;
        RECT 458.410 51.415 458.580 51.585 ;
        RECT 458.410 47.025 458.580 47.195 ;
        RECT 463.700 68.545 463.870 68.715 ;
        RECT 463.700 68.185 463.870 68.355 ;
        RECT 463.700 67.825 463.870 67.995 ;
        RECT 463.700 63.435 463.870 63.605 ;
        RECT 463.700 63.075 463.870 63.245 ;
        RECT 463.700 62.715 463.870 62.885 ;
        RECT 463.700 62.355 463.870 62.525 ;
        RECT 463.700 57.965 463.870 58.135 ;
        RECT 463.700 57.605 463.870 57.775 ;
        RECT 463.700 57.245 463.870 57.415 ;
        RECT 463.700 56.885 463.870 57.055 ;
        RECT 463.700 52.495 463.870 52.665 ;
        RECT 463.700 52.135 463.870 52.305 ;
        RECT 463.700 51.775 463.870 51.945 ;
        RECT 463.700 51.415 463.870 51.585 ;
        RECT 442.540 46.665 442.710 46.835 ;
        RECT 442.540 46.305 442.710 46.475 ;
        RECT 447.830 46.665 448.000 46.835 ;
        RECT 442.540 45.945 442.710 46.115 ;
        RECT 447.830 46.305 448.000 46.475 ;
        RECT 453.120 46.665 453.290 46.835 ;
        RECT 447.830 45.945 448.000 46.115 ;
        RECT 453.120 46.305 453.290 46.475 ;
        RECT 463.700 47.025 463.870 47.195 ;
        RECT 468.990 68.545 469.160 68.715 ;
        RECT 468.990 68.185 469.160 68.355 ;
        RECT 468.990 67.825 469.160 67.995 ;
        RECT 468.990 63.435 469.160 63.605 ;
        RECT 468.990 63.075 469.160 63.245 ;
        RECT 468.990 62.715 469.160 62.885 ;
        RECT 468.990 62.355 469.160 62.525 ;
        RECT 468.990 57.965 469.160 58.135 ;
        RECT 468.990 57.605 469.160 57.775 ;
        RECT 468.990 57.245 469.160 57.415 ;
        RECT 468.990 56.885 469.160 57.055 ;
        RECT 468.990 52.495 469.160 52.665 ;
        RECT 468.990 52.135 469.160 52.305 ;
        RECT 468.990 51.775 469.160 51.945 ;
        RECT 468.990 51.415 469.160 51.585 ;
        RECT 458.410 46.665 458.580 46.835 ;
        RECT 458.410 46.305 458.580 46.475 ;
        RECT 468.990 47.025 469.160 47.195 ;
        RECT 474.860 98.255 475.030 98.425 ;
        RECT 474.860 97.895 475.030 98.065 ;
        RECT 480.150 98.255 480.320 98.425 ;
        RECT 485.440 98.255 485.610 98.425 ;
        RECT 490.730 98.255 490.900 98.425 ;
        RECT 496.020 98.255 496.190 98.425 ;
        RECT 474.860 97.535 475.030 97.705 ;
        RECT 474.860 97.175 475.030 97.345 ;
        RECT 480.150 97.895 480.320 98.065 ;
        RECT 480.150 97.535 480.320 97.705 ;
        RECT 480.150 97.175 480.320 97.345 ;
        RECT 474.860 92.785 475.030 92.955 ;
        RECT 474.860 92.425 475.030 92.595 ;
        RECT 474.860 92.065 475.030 92.235 ;
        RECT 474.860 91.705 475.030 91.875 ;
        RECT 480.150 92.785 480.320 92.955 ;
        RECT 480.150 92.425 480.320 92.595 ;
        RECT 480.150 92.065 480.320 92.235 ;
        RECT 480.150 91.705 480.320 91.875 ;
        RECT 474.860 87.315 475.030 87.485 ;
        RECT 474.860 86.955 475.030 87.125 ;
        RECT 474.860 86.595 475.030 86.765 ;
        RECT 474.860 86.235 475.030 86.405 ;
        RECT 480.150 87.315 480.320 87.485 ;
        RECT 480.150 86.955 480.320 87.125 ;
        RECT 480.150 86.595 480.320 86.765 ;
        RECT 480.150 86.235 480.320 86.405 ;
        RECT 474.860 81.845 475.030 82.015 ;
        RECT 474.860 81.485 475.030 81.655 ;
        RECT 474.860 81.125 475.030 81.295 ;
        RECT 474.860 80.765 475.030 80.935 ;
        RECT 480.150 81.845 480.320 82.015 ;
        RECT 480.150 81.485 480.320 81.655 ;
        RECT 480.150 81.125 480.320 81.295 ;
        RECT 480.150 80.765 480.320 80.935 ;
        RECT 474.860 76.375 475.030 76.545 ;
        RECT 480.150 76.375 480.320 76.545 ;
        RECT 485.440 97.895 485.610 98.065 ;
        RECT 485.440 97.535 485.610 97.705 ;
        RECT 485.440 97.175 485.610 97.345 ;
        RECT 485.440 92.785 485.610 92.955 ;
        RECT 485.440 92.425 485.610 92.595 ;
        RECT 485.440 92.065 485.610 92.235 ;
        RECT 485.440 91.705 485.610 91.875 ;
        RECT 485.440 87.315 485.610 87.485 ;
        RECT 485.440 86.955 485.610 87.125 ;
        RECT 485.440 86.595 485.610 86.765 ;
        RECT 485.440 86.235 485.610 86.405 ;
        RECT 485.440 81.845 485.610 82.015 ;
        RECT 485.440 81.485 485.610 81.655 ;
        RECT 485.440 81.125 485.610 81.295 ;
        RECT 485.440 80.765 485.610 80.935 ;
        RECT 485.440 76.375 485.610 76.545 ;
        RECT 501.310 98.255 501.480 98.425 ;
        RECT 490.730 97.895 490.900 98.065 ;
        RECT 490.730 97.535 490.900 97.705 ;
        RECT 490.730 97.175 490.900 97.345 ;
        RECT 490.730 92.785 490.900 92.955 ;
        RECT 490.730 92.425 490.900 92.595 ;
        RECT 490.730 92.065 490.900 92.235 ;
        RECT 490.730 91.705 490.900 91.875 ;
        RECT 490.730 87.315 490.900 87.485 ;
        RECT 490.730 86.955 490.900 87.125 ;
        RECT 490.730 86.595 490.900 86.765 ;
        RECT 490.730 86.235 490.900 86.405 ;
        RECT 490.730 81.845 490.900 82.015 ;
        RECT 490.730 81.485 490.900 81.655 ;
        RECT 490.730 81.125 490.900 81.295 ;
        RECT 490.730 80.765 490.900 80.935 ;
        RECT 490.730 76.375 490.900 76.545 ;
        RECT 496.020 97.895 496.190 98.065 ;
        RECT 496.020 97.535 496.190 97.705 ;
        RECT 496.020 97.175 496.190 97.345 ;
        RECT 496.020 92.785 496.190 92.955 ;
        RECT 496.020 92.425 496.190 92.595 ;
        RECT 496.020 92.065 496.190 92.235 ;
        RECT 496.020 91.705 496.190 91.875 ;
        RECT 496.020 87.315 496.190 87.485 ;
        RECT 496.020 86.955 496.190 87.125 ;
        RECT 496.020 86.595 496.190 86.765 ;
        RECT 496.020 86.235 496.190 86.405 ;
        RECT 496.020 81.845 496.190 82.015 ;
        RECT 496.020 81.485 496.190 81.655 ;
        RECT 496.020 81.125 496.190 81.295 ;
        RECT 496.020 80.765 496.190 80.935 ;
        RECT 474.860 76.015 475.030 76.185 ;
        RECT 474.860 75.655 475.030 75.825 ;
        RECT 480.150 76.015 480.320 76.185 ;
        RECT 474.860 75.295 475.030 75.465 ;
        RECT 480.150 75.655 480.320 75.825 ;
        RECT 485.440 76.015 485.610 76.185 ;
        RECT 480.150 75.295 480.320 75.465 ;
        RECT 485.440 75.655 485.610 75.825 ;
        RECT 496.020 76.375 496.190 76.545 ;
        RECT 501.310 97.895 501.480 98.065 ;
        RECT 501.310 97.535 501.480 97.705 ;
        RECT 501.310 97.175 501.480 97.345 ;
        RECT 501.310 92.785 501.480 92.955 ;
        RECT 501.310 92.425 501.480 92.595 ;
        RECT 501.310 92.065 501.480 92.235 ;
        RECT 501.310 91.705 501.480 91.875 ;
        RECT 501.310 87.315 501.480 87.485 ;
        RECT 501.310 86.955 501.480 87.125 ;
        RECT 501.310 86.595 501.480 86.765 ;
        RECT 501.310 86.235 501.480 86.405 ;
        RECT 501.310 81.845 501.480 82.015 ;
        RECT 501.310 81.485 501.480 81.655 ;
        RECT 501.310 81.125 501.480 81.295 ;
        RECT 501.310 80.765 501.480 80.935 ;
        RECT 490.730 76.015 490.900 76.185 ;
        RECT 490.730 75.655 490.900 75.825 ;
        RECT 501.310 76.375 501.480 76.545 ;
        RECT 503.850 77.015 505.460 94.825 ;
        RECT 496.020 76.015 496.190 76.185 ;
        RECT 496.020 75.655 496.190 75.825 ;
        RECT 501.310 76.015 501.480 76.185 ;
        RECT 485.440 75.295 485.610 75.465 ;
        RECT 490.730 75.295 490.900 75.465 ;
        RECT 496.020 75.295 496.190 75.465 ;
        RECT 501.310 75.655 501.480 75.825 ;
        RECT 501.310 75.295 501.480 75.465 ;
        RECT 471.870 61.305 472.040 61.475 ;
        RECT 471.870 60.945 472.040 61.115 ;
        RECT 471.870 60.585 472.040 60.755 ;
        RECT 471.870 60.225 472.040 60.395 ;
        RECT 471.870 59.865 472.040 60.035 ;
        RECT 471.870 59.505 472.040 59.675 ;
        RECT 471.870 59.145 472.040 59.315 ;
        RECT 471.870 58.785 472.040 58.955 ;
        RECT 471.870 58.425 472.040 58.595 ;
        RECT 471.870 58.065 472.040 58.235 ;
        RECT 471.870 57.705 472.040 57.875 ;
        RECT 471.870 57.345 472.040 57.515 ;
        RECT 471.870 56.985 472.040 57.155 ;
        RECT 471.870 56.625 472.040 56.795 ;
        RECT 471.870 56.265 472.040 56.435 ;
        RECT 471.870 55.905 472.040 56.075 ;
        RECT 471.870 55.545 472.040 55.715 ;
        RECT 463.700 46.665 463.870 46.835 ;
        RECT 463.700 46.305 463.870 46.475 ;
        RECT 468.990 46.665 469.160 46.835 ;
        RECT 453.120 45.945 453.290 46.115 ;
        RECT 458.410 45.945 458.580 46.115 ;
        RECT 463.700 45.945 463.870 46.115 ;
        RECT 468.990 46.305 469.160 46.475 ;
        RECT 468.990 45.945 469.160 46.115 ;
        RECT 439.530 32.025 439.700 32.195 ;
        RECT 439.530 31.665 439.700 31.835 ;
        RECT 439.530 31.305 439.700 31.475 ;
        RECT 439.530 30.945 439.700 31.115 ;
        RECT 439.530 30.585 439.700 30.755 ;
        RECT 439.530 30.225 439.700 30.395 ;
        RECT 439.530 29.865 439.700 30.035 ;
        RECT 439.530 29.505 439.700 29.675 ;
        RECT 439.530 29.145 439.700 29.315 ;
        RECT 439.530 28.785 439.700 28.955 ;
        RECT 439.530 28.425 439.700 28.595 ;
        RECT 439.530 28.065 439.700 28.235 ;
        RECT 439.530 27.705 439.700 27.875 ;
        RECT 439.530 27.345 439.700 27.515 ;
        RECT 439.530 26.985 439.700 27.155 ;
        RECT 439.530 26.625 439.700 26.795 ;
        RECT 439.530 26.265 439.700 26.435 ;
        RECT 442.540 39.615 442.710 39.785 ;
        RECT 442.540 39.255 442.710 39.425 ;
        RECT 447.830 39.615 448.000 39.785 ;
        RECT 453.120 39.615 453.290 39.785 ;
        RECT 458.410 39.615 458.580 39.785 ;
        RECT 463.700 39.615 463.870 39.785 ;
        RECT 442.540 38.895 442.710 39.065 ;
        RECT 442.540 38.535 442.710 38.705 ;
        RECT 447.830 39.255 448.000 39.425 ;
        RECT 447.830 38.895 448.000 39.065 ;
        RECT 447.830 38.535 448.000 38.705 ;
        RECT 442.540 34.145 442.710 34.315 ;
        RECT 442.540 33.785 442.710 33.955 ;
        RECT 442.540 33.425 442.710 33.595 ;
        RECT 442.540 33.065 442.710 33.235 ;
        RECT 447.830 34.145 448.000 34.315 ;
        RECT 447.830 33.785 448.000 33.955 ;
        RECT 447.830 33.425 448.000 33.595 ;
        RECT 447.830 33.065 448.000 33.235 ;
        RECT 442.540 28.675 442.710 28.845 ;
        RECT 442.540 28.315 442.710 28.485 ;
        RECT 442.540 27.955 442.710 28.125 ;
        RECT 442.540 27.595 442.710 27.765 ;
        RECT 447.830 28.675 448.000 28.845 ;
        RECT 447.830 28.315 448.000 28.485 ;
        RECT 447.830 27.955 448.000 28.125 ;
        RECT 447.830 27.595 448.000 27.765 ;
        RECT 442.540 23.205 442.710 23.375 ;
        RECT 442.540 22.845 442.710 23.015 ;
        RECT 442.540 22.485 442.710 22.655 ;
        RECT 442.540 22.125 442.710 22.295 ;
        RECT 447.830 23.205 448.000 23.375 ;
        RECT 447.830 22.845 448.000 23.015 ;
        RECT 447.830 22.485 448.000 22.655 ;
        RECT 447.830 22.125 448.000 22.295 ;
        RECT 414.020 17.405 414.190 17.575 ;
        RECT 402.820 17.055 402.990 17.225 ;
        RECT 381.660 16.695 381.830 16.865 ;
        RECT 392.240 16.695 392.410 16.865 ;
        RECT 402.820 16.695 402.990 16.865 ;
        RECT 414.020 17.045 414.190 17.215 ;
        RECT 424.600 17.405 424.770 17.575 ;
        RECT 424.600 17.045 424.770 17.215 ;
        RECT 442.540 17.735 442.710 17.905 ;
        RECT 435.180 17.405 435.350 17.575 ;
        RECT 435.180 17.045 435.350 17.215 ;
        RECT 447.830 17.735 448.000 17.905 ;
        RECT 453.120 39.255 453.290 39.425 ;
        RECT 453.120 38.895 453.290 39.065 ;
        RECT 453.120 38.535 453.290 38.705 ;
        RECT 453.120 34.145 453.290 34.315 ;
        RECT 453.120 33.785 453.290 33.955 ;
        RECT 453.120 33.425 453.290 33.595 ;
        RECT 453.120 33.065 453.290 33.235 ;
        RECT 453.120 28.675 453.290 28.845 ;
        RECT 453.120 28.315 453.290 28.485 ;
        RECT 453.120 27.955 453.290 28.125 ;
        RECT 453.120 27.595 453.290 27.765 ;
        RECT 453.120 23.205 453.290 23.375 ;
        RECT 453.120 22.845 453.290 23.015 ;
        RECT 453.120 22.485 453.290 22.655 ;
        RECT 453.120 22.125 453.290 22.295 ;
        RECT 453.120 17.735 453.290 17.905 ;
        RECT 468.990 39.615 469.160 39.785 ;
        RECT 458.410 39.255 458.580 39.425 ;
        RECT 458.410 38.895 458.580 39.065 ;
        RECT 458.410 38.535 458.580 38.705 ;
        RECT 458.410 34.145 458.580 34.315 ;
        RECT 458.410 33.785 458.580 33.955 ;
        RECT 458.410 33.425 458.580 33.595 ;
        RECT 458.410 33.065 458.580 33.235 ;
        RECT 458.410 28.675 458.580 28.845 ;
        RECT 458.410 28.315 458.580 28.485 ;
        RECT 458.410 27.955 458.580 28.125 ;
        RECT 458.410 27.595 458.580 27.765 ;
        RECT 458.410 23.205 458.580 23.375 ;
        RECT 458.410 22.845 458.580 23.015 ;
        RECT 458.410 22.485 458.580 22.655 ;
        RECT 458.410 22.125 458.580 22.295 ;
        RECT 458.410 17.735 458.580 17.905 ;
        RECT 463.700 39.255 463.870 39.425 ;
        RECT 463.700 38.895 463.870 39.065 ;
        RECT 463.700 38.535 463.870 38.705 ;
        RECT 463.700 34.145 463.870 34.315 ;
        RECT 463.700 33.785 463.870 33.955 ;
        RECT 463.700 33.425 463.870 33.595 ;
        RECT 463.700 33.065 463.870 33.235 ;
        RECT 463.700 28.675 463.870 28.845 ;
        RECT 463.700 28.315 463.870 28.485 ;
        RECT 463.700 27.955 463.870 28.125 ;
        RECT 463.700 27.595 463.870 27.765 ;
        RECT 463.700 23.205 463.870 23.375 ;
        RECT 463.700 22.845 463.870 23.015 ;
        RECT 463.700 22.485 463.870 22.655 ;
        RECT 463.700 22.125 463.870 22.295 ;
        RECT 442.540 17.375 442.710 17.545 ;
        RECT 414.020 16.685 414.190 16.855 ;
        RECT 424.600 16.685 424.770 16.855 ;
        RECT 435.180 16.685 435.350 16.855 ;
        RECT 442.540 17.015 442.710 17.185 ;
        RECT 447.830 17.375 448.000 17.545 ;
        RECT 442.540 16.655 442.710 16.825 ;
        RECT 447.830 17.015 448.000 17.185 ;
        RECT 453.120 17.375 453.290 17.545 ;
        RECT 447.830 16.655 448.000 16.825 ;
        RECT 453.120 17.015 453.290 17.185 ;
        RECT 463.700 17.735 463.870 17.905 ;
        RECT 468.990 39.255 469.160 39.425 ;
        RECT 468.990 38.895 469.160 39.065 ;
        RECT 468.990 38.535 469.160 38.705 ;
        RECT 468.990 34.145 469.160 34.315 ;
        RECT 468.990 33.785 469.160 33.955 ;
        RECT 468.990 33.425 469.160 33.595 ;
        RECT 468.990 33.065 469.160 33.235 ;
        RECT 468.990 28.675 469.160 28.845 ;
        RECT 468.990 28.315 469.160 28.485 ;
        RECT 468.990 27.955 469.160 28.125 ;
        RECT 468.990 27.595 469.160 27.765 ;
        RECT 468.990 23.205 469.160 23.375 ;
        RECT 468.990 22.845 469.160 23.015 ;
        RECT 468.990 22.485 469.160 22.655 ;
        RECT 468.990 22.125 469.160 22.295 ;
        RECT 474.880 68.895 475.050 69.065 ;
        RECT 474.880 68.535 475.050 68.705 ;
        RECT 480.170 68.895 480.340 69.065 ;
        RECT 485.460 68.895 485.630 69.065 ;
        RECT 490.750 68.895 490.920 69.065 ;
        RECT 496.040 68.895 496.210 69.065 ;
        RECT 474.880 68.175 475.050 68.345 ;
        RECT 474.880 67.815 475.050 67.985 ;
        RECT 480.170 68.535 480.340 68.705 ;
        RECT 480.170 68.175 480.340 68.345 ;
        RECT 480.170 67.815 480.340 67.985 ;
        RECT 474.880 63.425 475.050 63.595 ;
        RECT 474.880 63.065 475.050 63.235 ;
        RECT 474.880 62.705 475.050 62.875 ;
        RECT 474.880 62.345 475.050 62.515 ;
        RECT 480.170 63.425 480.340 63.595 ;
        RECT 480.170 63.065 480.340 63.235 ;
        RECT 480.170 62.705 480.340 62.875 ;
        RECT 480.170 62.345 480.340 62.515 ;
        RECT 474.880 57.955 475.050 58.125 ;
        RECT 474.880 57.595 475.050 57.765 ;
        RECT 474.880 57.235 475.050 57.405 ;
        RECT 474.880 56.875 475.050 57.045 ;
        RECT 480.170 57.955 480.340 58.125 ;
        RECT 480.170 57.595 480.340 57.765 ;
        RECT 480.170 57.235 480.340 57.405 ;
        RECT 480.170 56.875 480.340 57.045 ;
        RECT 474.880 52.485 475.050 52.655 ;
        RECT 474.880 52.125 475.050 52.295 ;
        RECT 474.880 51.765 475.050 51.935 ;
        RECT 474.880 51.405 475.050 51.575 ;
        RECT 480.170 52.485 480.340 52.655 ;
        RECT 480.170 52.125 480.340 52.295 ;
        RECT 480.170 51.765 480.340 51.935 ;
        RECT 480.170 51.405 480.340 51.575 ;
        RECT 474.880 47.015 475.050 47.185 ;
        RECT 480.170 47.015 480.340 47.185 ;
        RECT 485.460 68.535 485.630 68.705 ;
        RECT 485.460 68.175 485.630 68.345 ;
        RECT 485.460 67.815 485.630 67.985 ;
        RECT 485.460 63.425 485.630 63.595 ;
        RECT 485.460 63.065 485.630 63.235 ;
        RECT 485.460 62.705 485.630 62.875 ;
        RECT 485.460 62.345 485.630 62.515 ;
        RECT 485.460 57.955 485.630 58.125 ;
        RECT 485.460 57.595 485.630 57.765 ;
        RECT 485.460 57.235 485.630 57.405 ;
        RECT 485.460 56.875 485.630 57.045 ;
        RECT 485.460 52.485 485.630 52.655 ;
        RECT 485.460 52.125 485.630 52.295 ;
        RECT 485.460 51.765 485.630 51.935 ;
        RECT 485.460 51.405 485.630 51.575 ;
        RECT 485.460 47.015 485.630 47.185 ;
        RECT 501.330 68.895 501.500 69.065 ;
        RECT 490.750 68.535 490.920 68.705 ;
        RECT 490.750 68.175 490.920 68.345 ;
        RECT 490.750 67.815 490.920 67.985 ;
        RECT 490.750 63.425 490.920 63.595 ;
        RECT 490.750 63.065 490.920 63.235 ;
        RECT 490.750 62.705 490.920 62.875 ;
        RECT 490.750 62.345 490.920 62.515 ;
        RECT 490.750 57.955 490.920 58.125 ;
        RECT 490.750 57.595 490.920 57.765 ;
        RECT 490.750 57.235 490.920 57.405 ;
        RECT 490.750 56.875 490.920 57.045 ;
        RECT 490.750 52.485 490.920 52.655 ;
        RECT 490.750 52.125 490.920 52.295 ;
        RECT 490.750 51.765 490.920 51.935 ;
        RECT 490.750 51.405 490.920 51.575 ;
        RECT 490.750 47.015 490.920 47.185 ;
        RECT 496.040 68.535 496.210 68.705 ;
        RECT 496.040 68.175 496.210 68.345 ;
        RECT 496.040 67.815 496.210 67.985 ;
        RECT 496.040 63.425 496.210 63.595 ;
        RECT 496.040 63.065 496.210 63.235 ;
        RECT 496.040 62.705 496.210 62.875 ;
        RECT 496.040 62.345 496.210 62.515 ;
        RECT 496.040 57.955 496.210 58.125 ;
        RECT 496.040 57.595 496.210 57.765 ;
        RECT 496.040 57.235 496.210 57.405 ;
        RECT 496.040 56.875 496.210 57.045 ;
        RECT 496.040 52.485 496.210 52.655 ;
        RECT 496.040 52.125 496.210 52.295 ;
        RECT 496.040 51.765 496.210 51.935 ;
        RECT 496.040 51.405 496.210 51.575 ;
        RECT 474.880 46.655 475.050 46.825 ;
        RECT 474.880 46.295 475.050 46.465 ;
        RECT 480.170 46.655 480.340 46.825 ;
        RECT 474.880 45.935 475.050 46.105 ;
        RECT 480.170 46.295 480.340 46.465 ;
        RECT 485.460 46.655 485.630 46.825 ;
        RECT 480.170 45.935 480.340 46.105 ;
        RECT 485.460 46.295 485.630 46.465 ;
        RECT 496.040 47.015 496.210 47.185 ;
        RECT 501.330 68.535 501.500 68.705 ;
        RECT 501.330 68.175 501.500 68.345 ;
        RECT 501.330 67.815 501.500 67.985 ;
        RECT 501.330 63.425 501.500 63.595 ;
        RECT 501.330 63.065 501.500 63.235 ;
        RECT 501.330 62.705 501.500 62.875 ;
        RECT 501.330 62.345 501.500 62.515 ;
        RECT 501.330 57.955 501.500 58.125 ;
        RECT 501.330 57.595 501.500 57.765 ;
        RECT 501.330 57.235 501.500 57.405 ;
        RECT 501.330 56.875 501.500 57.045 ;
        RECT 501.330 52.485 501.500 52.655 ;
        RECT 501.330 52.125 501.500 52.295 ;
        RECT 501.330 51.765 501.500 51.935 ;
        RECT 501.330 51.405 501.500 51.575 ;
        RECT 490.750 46.655 490.920 46.825 ;
        RECT 490.750 46.295 490.920 46.465 ;
        RECT 501.330 47.015 501.500 47.185 ;
        RECT 504.490 48.955 505.380 67.125 ;
        RECT 496.040 46.655 496.210 46.825 ;
        RECT 496.040 46.295 496.210 46.465 ;
        RECT 501.330 46.655 501.500 46.825 ;
        RECT 485.460 45.935 485.630 46.105 ;
        RECT 490.750 45.935 490.920 46.105 ;
        RECT 496.040 45.935 496.210 46.105 ;
        RECT 501.330 46.295 501.500 46.465 ;
        RECT 501.330 45.935 501.500 46.105 ;
        RECT 471.890 32.015 472.060 32.185 ;
        RECT 471.890 31.655 472.060 31.825 ;
        RECT 471.890 31.295 472.060 31.465 ;
        RECT 471.890 30.935 472.060 31.105 ;
        RECT 471.890 30.575 472.060 30.745 ;
        RECT 471.890 30.215 472.060 30.385 ;
        RECT 471.890 29.855 472.060 30.025 ;
        RECT 471.890 29.495 472.060 29.665 ;
        RECT 471.890 29.135 472.060 29.305 ;
        RECT 471.890 28.775 472.060 28.945 ;
        RECT 471.890 28.415 472.060 28.585 ;
        RECT 471.890 28.055 472.060 28.225 ;
        RECT 471.890 27.695 472.060 27.865 ;
        RECT 471.890 27.335 472.060 27.505 ;
        RECT 471.890 26.975 472.060 27.145 ;
        RECT 471.890 26.615 472.060 26.785 ;
        RECT 471.890 26.255 472.060 26.425 ;
        RECT 474.900 39.605 475.070 39.775 ;
        RECT 474.900 39.245 475.070 39.415 ;
        RECT 480.190 39.605 480.360 39.775 ;
        RECT 485.480 39.605 485.650 39.775 ;
        RECT 490.770 39.605 490.940 39.775 ;
        RECT 496.060 39.605 496.230 39.775 ;
        RECT 474.900 38.885 475.070 39.055 ;
        RECT 474.900 38.525 475.070 38.695 ;
        RECT 480.190 39.245 480.360 39.415 ;
        RECT 480.190 38.885 480.360 39.055 ;
        RECT 480.190 38.525 480.360 38.695 ;
        RECT 474.900 34.135 475.070 34.305 ;
        RECT 474.900 33.775 475.070 33.945 ;
        RECT 474.900 33.415 475.070 33.585 ;
        RECT 474.900 33.055 475.070 33.225 ;
        RECT 480.190 34.135 480.360 34.305 ;
        RECT 480.190 33.775 480.360 33.945 ;
        RECT 480.190 33.415 480.360 33.585 ;
        RECT 480.190 33.055 480.360 33.225 ;
        RECT 474.900 28.665 475.070 28.835 ;
        RECT 474.900 28.305 475.070 28.475 ;
        RECT 474.900 27.945 475.070 28.115 ;
        RECT 474.900 27.585 475.070 27.755 ;
        RECT 480.190 28.665 480.360 28.835 ;
        RECT 480.190 28.305 480.360 28.475 ;
        RECT 480.190 27.945 480.360 28.115 ;
        RECT 480.190 27.585 480.360 27.755 ;
        RECT 474.900 23.195 475.070 23.365 ;
        RECT 474.900 22.835 475.070 23.005 ;
        RECT 474.900 22.475 475.070 22.645 ;
        RECT 474.900 22.115 475.070 22.285 ;
        RECT 480.190 23.195 480.360 23.365 ;
        RECT 480.190 22.835 480.360 23.005 ;
        RECT 480.190 22.475 480.360 22.645 ;
        RECT 480.190 22.115 480.360 22.285 ;
        RECT 458.410 17.375 458.580 17.545 ;
        RECT 458.410 17.015 458.580 17.185 ;
        RECT 468.990 17.735 469.160 17.905 ;
        RECT 474.900 17.725 475.070 17.895 ;
        RECT 463.700 17.375 463.870 17.545 ;
        RECT 463.700 17.015 463.870 17.185 ;
        RECT 468.990 17.375 469.160 17.545 ;
        RECT 453.120 16.655 453.290 16.825 ;
        RECT 458.410 16.655 458.580 16.825 ;
        RECT 463.700 16.655 463.870 16.825 ;
        RECT 468.990 17.015 469.160 17.185 ;
        RECT 480.190 17.725 480.360 17.895 ;
        RECT 485.480 39.245 485.650 39.415 ;
        RECT 485.480 38.885 485.650 39.055 ;
        RECT 485.480 38.525 485.650 38.695 ;
        RECT 485.480 34.135 485.650 34.305 ;
        RECT 485.480 33.775 485.650 33.945 ;
        RECT 485.480 33.415 485.650 33.585 ;
        RECT 485.480 33.055 485.650 33.225 ;
        RECT 485.480 28.665 485.650 28.835 ;
        RECT 485.480 28.305 485.650 28.475 ;
        RECT 485.480 27.945 485.650 28.115 ;
        RECT 485.480 27.585 485.650 27.755 ;
        RECT 485.480 23.195 485.650 23.365 ;
        RECT 485.480 22.835 485.650 23.005 ;
        RECT 485.480 22.475 485.650 22.645 ;
        RECT 485.480 22.115 485.650 22.285 ;
        RECT 485.480 17.725 485.650 17.895 ;
        RECT 501.350 39.605 501.520 39.775 ;
        RECT 490.770 39.245 490.940 39.415 ;
        RECT 490.770 38.885 490.940 39.055 ;
        RECT 490.770 38.525 490.940 38.695 ;
        RECT 490.770 34.135 490.940 34.305 ;
        RECT 490.770 33.775 490.940 33.945 ;
        RECT 490.770 33.415 490.940 33.585 ;
        RECT 490.770 33.055 490.940 33.225 ;
        RECT 490.770 28.665 490.940 28.835 ;
        RECT 490.770 28.305 490.940 28.475 ;
        RECT 490.770 27.945 490.940 28.115 ;
        RECT 490.770 27.585 490.940 27.755 ;
        RECT 490.770 23.195 490.940 23.365 ;
        RECT 490.770 22.835 490.940 23.005 ;
        RECT 490.770 22.475 490.940 22.645 ;
        RECT 490.770 22.115 490.940 22.285 ;
        RECT 490.770 17.725 490.940 17.895 ;
        RECT 496.060 39.245 496.230 39.415 ;
        RECT 496.060 38.885 496.230 39.055 ;
        RECT 496.060 38.525 496.230 38.695 ;
        RECT 496.060 34.135 496.230 34.305 ;
        RECT 496.060 33.775 496.230 33.945 ;
        RECT 496.060 33.415 496.230 33.585 ;
        RECT 496.060 33.055 496.230 33.225 ;
        RECT 496.060 28.665 496.230 28.835 ;
        RECT 496.060 28.305 496.230 28.475 ;
        RECT 496.060 27.945 496.230 28.115 ;
        RECT 496.060 27.585 496.230 27.755 ;
        RECT 496.060 23.195 496.230 23.365 ;
        RECT 496.060 22.835 496.230 23.005 ;
        RECT 496.060 22.475 496.230 22.645 ;
        RECT 496.060 22.115 496.230 22.285 ;
        RECT 474.900 17.365 475.070 17.535 ;
        RECT 468.990 16.655 469.160 16.825 ;
        RECT 474.900 17.005 475.070 17.175 ;
        RECT 480.190 17.365 480.360 17.535 ;
        RECT 474.900 16.645 475.070 16.815 ;
        RECT 480.190 17.005 480.360 17.175 ;
        RECT 485.480 17.365 485.650 17.535 ;
        RECT 480.190 16.645 480.360 16.815 ;
        RECT 485.480 17.005 485.650 17.175 ;
        RECT 496.060 17.725 496.230 17.895 ;
        RECT 501.350 39.245 501.520 39.415 ;
        RECT 501.350 38.885 501.520 39.055 ;
        RECT 501.350 38.525 501.520 38.695 ;
        RECT 501.350 34.135 501.520 34.305 ;
        RECT 501.350 33.775 501.520 33.945 ;
        RECT 501.350 33.415 501.520 33.585 ;
        RECT 501.350 33.055 501.520 33.225 ;
        RECT 501.350 28.665 501.520 28.835 ;
        RECT 501.350 28.305 501.520 28.475 ;
        RECT 501.350 27.945 501.520 28.115 ;
        RECT 501.350 27.585 501.520 27.755 ;
        RECT 501.350 23.195 501.520 23.365 ;
        RECT 501.350 22.835 501.520 23.005 ;
        RECT 501.350 22.475 501.520 22.645 ;
        RECT 501.350 22.115 501.520 22.285 ;
        RECT 490.770 17.365 490.940 17.535 ;
        RECT 490.770 17.005 490.940 17.175 ;
        RECT 501.350 17.725 501.520 17.895 ;
        RECT 504.545 18.070 505.435 36.240 ;
        RECT 496.060 17.365 496.230 17.535 ;
        RECT 496.060 17.005 496.230 17.175 ;
        RECT 501.350 17.365 501.520 17.535 ;
        RECT 485.480 16.645 485.650 16.815 ;
        RECT 490.770 16.645 490.940 16.815 ;
        RECT 496.060 16.645 496.230 16.815 ;
        RECT 501.350 17.005 501.520 17.175 ;
        RECT 501.350 16.645 501.520 16.815 ;
        RECT 199.260 -6.060 207.710 -2.650 ;
        RECT 297.680 -3.330 302.890 -1.000 ;
        RECT 368.500 -0.985 379.110 3.865 ;
      LAYER met1 ;
        RECT -97.390 354.515 -97.160 355.730 ;
        RECT -94.810 354.515 -94.580 355.730 ;
        RECT -92.230 354.555 -92.000 355.730 ;
        RECT -89.650 354.575 -89.420 355.730 ;
        RECT -87.070 354.645 -86.840 355.730 ;
        RECT -97.395 354.150 -97.160 354.515 ;
        RECT -94.855 354.150 -94.580 354.515 ;
        RECT -92.255 354.150 -92.000 354.555 ;
        RECT -89.685 354.150 -89.420 354.575 ;
        RECT -87.105 354.150 -86.840 354.645 ;
        RECT -84.490 354.555 -84.260 355.730 ;
        RECT -84.505 354.150 -84.260 354.555 ;
        RECT -81.910 354.645 -81.680 355.730 ;
        RECT -81.910 354.150 -81.675 354.645 ;
        RECT -79.330 354.575 -79.100 355.730 ;
        RECT -76.750 354.575 -76.520 355.730 ;
        RECT -74.170 354.605 -73.940 355.730 ;
        RECT -79.330 354.150 -79.075 354.575 ;
        RECT -76.750 354.150 -76.485 354.575 ;
        RECT -97.395 353.255 -97.165 354.150 ;
        RECT -94.855 353.255 -94.625 354.150 ;
        RECT -92.255 353.255 -92.025 354.150 ;
        RECT -89.685 353.255 -89.455 354.150 ;
        RECT -87.105 353.255 -86.875 354.150 ;
        RECT -84.505 353.255 -84.275 354.150 ;
        RECT -81.905 353.255 -81.675 354.150 ;
        RECT -79.305 353.255 -79.075 354.150 ;
        RECT -76.715 353.255 -76.485 354.150 ;
        RECT -74.215 354.150 -73.940 354.605 ;
        RECT -71.590 354.555 -71.360 355.730 ;
        RECT -71.595 354.150 -71.360 354.555 ;
        RECT -74.215 353.255 -73.985 354.150 ;
        RECT -71.595 353.255 -71.365 354.150 ;
        RECT -97.415 352.955 -71.365 353.255 ;
        RECT -97.395 352.935 -97.165 352.955 ;
        RECT -94.855 352.935 -94.625 352.955 ;
        RECT -82.565 352.280 -82.375 352.955 ;
        RECT -96.900 352.050 -96.360 352.280 ;
        RECT -95.610 352.050 -95.070 352.280 ;
        RECT -94.320 352.050 -93.780 352.280 ;
        RECT -93.030 352.050 -92.490 352.280 ;
        RECT -91.740 352.050 -91.200 352.280 ;
        RECT -90.450 352.050 -89.910 352.280 ;
        RECT -89.160 352.050 -88.620 352.280 ;
        RECT -87.870 352.050 -87.330 352.280 ;
        RECT -86.580 352.050 -86.040 352.280 ;
        RECT -85.290 352.050 -84.750 352.280 ;
        RECT -84.000 352.050 -83.460 352.280 ;
        RECT -82.710 352.050 -82.170 352.280 ;
        RECT -81.420 352.050 -80.880 352.280 ;
        RECT -80.130 352.050 -79.590 352.280 ;
        RECT -78.840 352.050 -78.300 352.280 ;
        RECT -77.550 352.050 -77.010 352.280 ;
        RECT -76.260 352.050 -75.720 352.280 ;
        RECT -74.970 352.050 -74.430 352.280 ;
        RECT -73.680 352.050 -73.140 352.280 ;
        RECT -72.390 352.050 -71.850 352.280 ;
        RECT -91.040 349.600 -77.450 351.780 ;
        RECT 653.970 351.340 655.410 351.485 ;
        RECT 653.910 351.270 655.410 351.340 ;
        RECT 657.550 351.270 672.910 351.475 ;
        RECT 653.910 351.250 672.910 351.270 ;
        RECT 675.600 351.260 690.960 351.435 ;
        RECT 693.190 351.260 708.550 351.455 ;
        RECT 675.600 351.250 708.550 351.260 ;
        RECT 653.910 351.210 708.550 351.250 ;
        RECT 711.040 351.230 726.400 351.455 ;
        RECT 729.300 351.250 744.660 351.455 ;
        RECT 747.070 351.250 762.430 351.425 ;
        RECT 729.300 351.230 762.430 351.250 ;
        RECT 711.040 351.210 762.430 351.230 ;
        RECT 653.910 351.120 762.430 351.210 ;
        RECT 765.110 351.150 780.470 351.345 ;
        RECT 783.270 351.160 798.630 351.385 ;
        RECT 801.650 351.190 817.010 351.395 ;
        RECT 820.450 351.190 835.810 351.375 ;
        RECT 801.650 351.160 835.810 351.190 ;
        RECT 783.270 351.150 835.810 351.160 ;
        RECT 765.110 351.120 835.810 351.150 ;
        RECT 653.910 351.105 835.810 351.120 ;
        RECT 653.910 350.965 657.970 351.105 ;
        RECT 671.630 351.085 835.810 351.105 ;
        RECT 671.630 351.065 693.840 351.085 ;
        RECT 671.630 350.965 676.270 351.065 ;
        RECT 653.910 350.925 676.270 350.965 ;
        RECT 689.200 350.945 693.840 351.065 ;
        RECT 707.050 350.945 711.690 351.085 ;
        RECT 725.410 350.945 730.050 351.085 ;
        RECT 742.840 351.055 835.810 351.085 ;
        RECT 742.840 350.945 747.480 351.055 ;
        RECT 689.200 350.925 747.480 350.945 ;
        RECT 653.910 350.915 747.480 350.925 ;
        RECT 760.980 351.025 835.810 351.055 ;
        RECT 760.980 351.015 802.020 351.025 ;
        RECT 760.980 350.975 785.070 351.015 ;
        RECT 760.980 350.915 765.620 350.975 ;
        RECT 653.910 350.850 765.620 350.915 ;
        RECT 653.910 350.840 690.960 350.850 ;
        RECT 653.910 350.820 672.910 350.840 ;
        RECT 653.910 350.770 655.410 350.820 ;
        RECT 653.970 350.745 655.410 350.770 ;
        RECT 657.550 350.735 672.910 350.820 ;
        RECT 675.600 350.695 690.960 350.840 ;
        RECT 693.190 350.840 765.620 350.850 ;
        RECT 693.190 350.820 744.660 350.840 ;
        RECT 693.190 350.800 726.400 350.820 ;
        RECT 693.190 350.715 708.550 350.800 ;
        RECT 711.040 350.715 726.400 350.800 ;
        RECT 729.300 350.715 744.660 350.820 ;
        RECT 747.070 350.835 765.620 350.840 ;
        RECT 779.340 350.875 785.070 350.975 ;
        RECT 797.380 350.885 802.020 351.015 ;
        RECT 816.260 351.005 835.810 351.025 ;
        RECT 816.260 350.885 820.900 351.005 ;
        RECT 838.920 350.985 840.360 351.355 ;
        RECT 797.380 350.875 820.900 350.885 ;
        RECT 779.340 350.865 820.900 350.875 ;
        RECT 779.340 350.835 835.810 350.865 ;
        RECT 839.510 350.845 840.030 350.985 ;
        RECT 747.070 350.780 835.810 350.835 ;
        RECT 747.070 350.750 817.010 350.780 ;
        RECT 747.070 350.740 798.630 350.750 ;
        RECT 747.070 350.710 780.470 350.740 ;
        RECT 747.070 350.685 762.430 350.710 ;
        RECT 765.110 350.605 780.470 350.710 ;
        RECT 781.790 343.100 782.420 350.740 ;
        RECT 783.270 350.645 798.630 350.740 ;
        RECT 801.650 350.655 817.010 350.750 ;
        RECT 820.450 350.750 835.810 350.780 ;
        RECT 838.920 350.750 840.360 350.845 ;
        RECT 784.360 350.070 785.070 350.645 ;
        RECT 820.450 350.635 840.360 350.750 ;
        RECT 835.540 350.615 840.360 350.635 ;
        RECT 835.540 350.540 839.150 350.615 ;
        RECT 783.830 343.150 787.190 343.215 ;
        RECT 790.390 343.150 791.830 343.245 ;
        RECT 793.850 343.150 809.210 343.305 ;
        RECT 783.830 343.100 809.210 343.150 ;
        RECT 781.790 343.040 809.210 343.100 ;
        RECT 813.210 343.040 828.570 343.215 ;
        RECT 781.790 342.935 828.570 343.040 ;
        RECT 781.790 342.845 794.650 342.935 ;
        RECT 781.790 342.705 784.150 342.845 ;
        RECT 785.150 342.795 794.650 342.845 ;
        RECT 807.920 342.845 828.570 342.935 ;
        RECT 807.920 342.795 813.780 342.845 ;
        RECT 785.150 342.705 813.780 342.795 ;
        RECT 781.790 342.690 828.570 342.705 ;
        RECT 781.790 342.490 787.190 342.690 ;
        RECT 790.390 342.505 791.830 342.690 ;
        RECT 793.850 342.580 828.570 342.690 ;
        RECT 793.850 342.565 809.210 342.580 ;
        RECT 783.830 342.475 787.190 342.490 ;
        RECT 813.210 342.475 828.570 342.580 ;
        RECT 853.880 337.820 854.110 337.920 ;
        RECT 853.880 337.540 854.150 337.820 ;
        RECT 853.900 336.450 854.150 337.540 ;
        RECT 853.880 336.070 854.150 336.450 ;
        RECT 853.900 334.980 854.150 336.070 ;
        RECT 853.880 334.600 854.150 334.980 ;
        RECT 853.900 333.510 854.150 334.600 ;
        RECT 853.880 333.130 854.150 333.510 ;
        RECT 853.900 332.040 854.150 333.130 ;
        RECT 853.880 331.660 854.150 332.040 ;
        RECT 853.900 330.570 854.150 331.660 ;
        RECT 853.880 330.190 854.150 330.570 ;
        RECT 678.350 329.160 679.130 329.690 ;
        RECT 663.190 328.755 666.550 329.125 ;
        RECT 668.820 328.755 672.180 329.125 ;
        RECT 677.800 329.025 679.130 329.160 ;
        RECT 853.900 329.100 854.150 330.190 ;
        RECT 674.580 328.970 679.130 329.025 ;
        RECT 664.460 328.615 666.010 328.755 ;
        RECT 670.460 328.615 671.220 328.755 ;
        RECT 674.580 328.655 677.940 328.970 ;
        RECT 678.350 328.920 679.130 328.970 ;
        RECT 681.610 328.695 685.450 329.065 ;
        RECT 687.470 328.705 690.830 329.075 ;
        RECT 853.880 328.720 854.150 329.100 ;
        RECT 635.260 327.415 636.700 327.785 ;
        RECT 639.450 327.505 640.890 327.875 ;
        RECT 595.370 326.965 596.810 327.335 ;
        RECT 635.390 327.275 635.570 327.415 ;
        RECT 639.550 327.365 639.690 327.505 ;
        RECT 643.550 327.485 644.990 327.855 ;
        RECT 635.260 327.250 636.700 327.275 ;
        RECT 639.450 327.250 640.890 327.365 ;
        RECT 643.970 327.345 644.210 327.485 ;
        RECT 643.550 327.260 644.990 327.345 ;
        RECT 645.940 327.260 646.590 328.510 ;
        RECT 663.190 328.385 666.550 328.615 ;
        RECT 668.820 328.385 672.180 328.615 ;
        RECT 675.810 328.515 676.570 328.655 ;
        RECT 683.490 328.555 684.250 328.695 ;
        RECT 689.220 328.565 689.980 328.705 ;
        RECT 670.770 328.370 671.040 328.385 ;
        RECT 674.580 328.285 677.940 328.515 ;
        RECT 681.610 328.325 685.450 328.555 ;
        RECT 687.470 328.335 690.830 328.565 ;
        RECT 853.900 327.630 854.150 328.720 ;
        RECT 635.260 327.240 643.180 327.250 ;
        RECT 643.550 327.240 646.590 327.260 ;
        RECT 635.260 327.200 646.590 327.240 ;
        RECT 596.610 326.825 596.750 326.965 ;
        RECT 595.370 326.595 596.810 326.825 ;
        RECT 596.610 326.170 596.750 326.595 ;
        RECT 596.550 325.810 597.240 326.170 ;
        RECT 605.330 322.580 606.220 327.050 ;
        RECT 614.990 324.320 615.220 324.700 ;
        RECT 616.570 324.320 616.800 324.700 ;
        RECT 615.010 323.230 615.170 324.320 ;
        RECT 616.590 323.230 616.750 324.320 ;
        RECT 614.990 322.850 615.220 323.230 ;
        RECT 616.570 322.850 616.800 323.230 ;
        RECT 625.510 323.050 626.430 327.180 ;
        RECT 635.260 327.135 646.320 327.200 ;
        RECT 635.260 327.045 639.750 327.135 ;
        RECT 635.310 326.450 635.540 327.045 ;
        RECT 636.440 327.030 639.750 327.045 ;
        RECT 640.650 327.030 646.320 327.135 ;
        RECT 643.150 327.020 644.720 327.030 ;
        RECT 645.100 327.020 646.320 327.030 ;
        RECT 635.080 326.100 635.580 326.450 ;
        RECT 640.340 323.430 640.570 323.810 ;
        RECT 644.390 323.570 644.620 323.860 ;
        RECT 644.390 323.480 644.640 323.570 ;
        RECT 627.010 323.050 627.560 323.140 ;
        RECT 615.010 322.680 615.180 322.850 ;
        RECT 616.620 322.680 616.790 322.850 ;
        RECT 625.510 322.740 627.560 323.050 ;
        RECT 625.510 322.680 626.430 322.740 ;
        RECT 605.430 321.530 605.900 322.580 ;
        RECT 614.950 322.540 616.810 322.680 ;
        RECT 615.700 321.530 616.040 322.540 ;
        RECT 625.700 321.530 626.170 322.680 ;
        RECT 627.010 322.600 627.560 322.740 ;
        RECT 640.380 321.540 640.560 323.430 ;
        RECT 644.400 321.540 644.640 323.480 ;
        RECT 658.760 322.455 660.200 322.825 ;
        RECT 658.980 322.315 659.720 322.455 ;
        RECT 663.660 322.415 665.100 322.785 ;
        RECT 668.250 322.780 669.690 322.815 ;
        RECT 670.710 322.780 671.290 323.210 ;
        RECT 668.250 322.480 671.290 322.780 ;
        RECT 668.250 322.445 669.690 322.480 ;
        RECT 658.760 322.085 660.200 322.315 ;
        RECT 663.950 322.275 664.690 322.415 ;
        RECT 668.810 322.305 669.080 322.445 ;
        RECT 670.710 322.370 671.290 322.480 ;
        RECT 672.790 322.425 674.230 322.795 ;
        RECT 676.220 322.435 680.060 322.805 ;
        RECT 681.990 322.435 685.350 322.805 ;
        RECT 687.440 322.750 690.800 322.805 ;
        RECT 691.410 322.750 692.140 323.200 ;
        RECT 687.440 322.530 692.140 322.750 ;
        RECT 687.440 322.435 690.800 322.530 ;
        RECT 691.410 322.460 692.140 322.530 ;
        RECT 692.750 322.455 696.110 322.825 ;
        RECT 663.660 322.045 665.100 322.275 ;
        RECT 668.250 322.180 669.690 322.305 ;
        RECT 673.200 322.285 673.470 322.425 ;
        RECT 677.620 322.295 677.890 322.435 ;
        RECT 684.250 322.295 684.520 322.435 ;
        RECT 688.930 322.295 689.930 322.435 ;
        RECT 694.890 322.315 695.160 322.455 ;
        RECT 692.750 322.300 696.110 322.315 ;
        RECT 697.870 322.300 698.240 322.340 ;
        RECT 672.790 322.280 674.230 322.285 ;
        RECT 676.220 322.280 680.060 322.295 ;
        RECT 672.790 322.240 680.060 322.280 ;
        RECT 681.990 322.260 685.350 322.295 ;
        RECT 687.440 322.260 690.800 322.295 ;
        RECT 681.990 322.240 690.800 322.260 ;
        RECT 672.790 322.210 690.800 322.240 ;
        RECT 692.750 322.210 698.240 322.300 ;
        RECT 672.790 322.180 698.240 322.210 ;
        RECT 668.250 322.085 698.240 322.180 ;
        RECT 668.250 322.075 693.340 322.085 ;
        RECT 669.570 322.070 693.340 322.075 ;
        RECT 669.570 322.055 674.230 322.070 ;
        RECT 676.220 322.065 693.340 322.070 ;
        RECT 669.570 322.030 672.940 322.055 ;
        RECT 679.760 322.030 682.710 322.065 ;
        RECT 685.030 322.050 687.980 322.065 ;
        RECT 690.390 322.000 693.340 322.065 ;
        RECT 646.180 321.540 649.390 322.000 ;
        RECT 695.920 321.970 698.240 322.085 ;
        RECT 632.020 321.530 643.570 321.540 ;
        RECT 643.810 321.530 649.390 321.540 ;
        RECT 600.330 320.370 649.390 321.530 ;
        RECT 632.020 320.340 649.390 320.370 ;
        RECT 646.180 319.610 649.390 320.340 ;
        RECT 661.400 316.575 665.240 316.945 ;
        RECT 667.220 316.890 670.580 316.955 ;
        RECT 671.050 316.890 671.780 317.180 ;
        RECT 667.220 316.620 671.780 316.890 ;
        RECT 667.220 316.585 670.580 316.620 ;
        RECT 661.690 316.435 663.730 316.575 ;
        RECT 668.830 316.445 669.100 316.585 ;
        RECT 671.050 316.510 671.780 316.620 ;
        RECT 672.660 316.595 676.020 316.965 ;
        RECT 677.980 316.960 681.340 316.965 ;
        RECT 681.900 316.960 682.670 317.130 ;
        RECT 677.980 316.670 682.670 316.960 ;
        RECT 677.980 316.595 681.340 316.670 ;
        RECT 674.450 316.455 674.720 316.595 ;
        RECT 679.330 316.455 680.170 316.595 ;
        RECT 681.900 316.490 682.670 316.670 ;
        RECT 683.330 316.595 686.690 316.965 ;
        RECT 689.150 316.910 691.550 316.945 ;
        RECT 692.160 316.910 693.000 317.140 ;
        RECT 685.340 316.455 685.610 316.595 ;
        RECT 689.150 316.590 693.000 316.910 ;
        RECT 689.150 316.575 691.550 316.590 ;
        RECT 661.400 316.360 665.240 316.435 ;
        RECT 667.220 316.360 670.580 316.445 ;
        RECT 661.400 316.340 670.580 316.360 ;
        RECT 672.660 316.340 676.020 316.455 ;
        RECT 677.980 316.350 681.340 316.455 ;
        RECT 683.330 316.350 686.690 316.455 ;
        RECT 690.380 316.435 690.650 316.575 ;
        RECT 692.160 316.530 693.000 316.590 ;
        RECT 693.550 316.575 695.950 316.945 ;
        RECT 694.820 316.435 695.090 316.575 ;
        RECT 661.400 316.330 676.020 316.340 ;
        RECT 677.010 316.330 677.400 316.340 ;
        RECT 677.980 316.330 686.690 316.350 ;
        RECT 661.400 316.310 686.690 316.330 ;
        RECT 689.150 316.360 691.550 316.435 ;
        RECT 693.550 316.380 695.950 316.435 ;
        RECT 697.870 316.380 698.240 321.970 ;
        RECT 693.550 316.360 698.240 316.380 ;
        RECT 689.150 316.310 698.240 316.360 ;
        RECT 661.400 316.225 698.240 316.310 ;
        RECT 661.400 316.215 672.760 316.225 ;
        RECT 661.400 316.205 667.450 316.215 ;
        RECT 665.060 316.170 667.450 316.205 ;
        RECT 670.370 316.150 672.760 316.215 ;
        RECT 675.740 316.140 678.130 316.225 ;
        RECT 681.070 316.160 683.460 316.225 ;
        RECT 686.470 316.205 698.240 316.225 ;
        RECT 635.110 309.245 636.550 309.615 ;
        RECT 639.300 309.335 640.740 309.705 ;
        RECT 595.220 308.795 596.660 309.165 ;
        RECT 635.240 309.105 635.420 309.245 ;
        RECT 639.400 309.195 639.540 309.335 ;
        RECT 643.400 309.315 644.840 309.685 ;
        RECT 635.110 309.080 636.550 309.105 ;
        RECT 639.300 309.080 640.740 309.195 ;
        RECT 643.820 309.175 644.060 309.315 ;
        RECT 643.400 309.080 644.840 309.175 ;
        RECT 646.040 309.080 646.680 310.320 ;
        RECT 635.110 309.070 643.030 309.080 ;
        RECT 643.400 309.070 646.680 309.080 ;
        RECT 596.460 308.655 596.600 308.795 ;
        RECT 595.220 308.425 596.660 308.655 ;
        RECT 596.460 308.000 596.600 308.425 ;
        RECT 596.400 307.640 597.090 308.000 ;
        RECT 605.180 304.410 606.070 308.880 ;
        RECT 614.840 306.150 615.070 306.530 ;
        RECT 616.420 306.150 616.650 306.530 ;
        RECT 614.860 305.060 615.020 306.150 ;
        RECT 616.440 305.060 616.600 306.150 ;
        RECT 614.840 304.680 615.070 305.060 ;
        RECT 616.420 304.680 616.650 305.060 ;
        RECT 625.360 304.880 626.280 309.010 ;
        RECT 635.110 308.965 646.680 309.070 ;
        RECT 635.110 308.875 639.600 308.965 ;
        RECT 635.160 308.280 635.390 308.875 ;
        RECT 636.290 308.860 639.600 308.875 ;
        RECT 640.500 308.960 646.680 308.965 ;
        RECT 640.500 308.860 646.320 308.960 ;
        RECT 643.000 308.850 644.570 308.860 ;
        RECT 645.100 308.840 646.320 308.860 ;
        RECT 634.930 307.930 635.430 308.280 ;
        RECT 640.190 305.260 640.420 305.640 ;
        RECT 644.240 305.400 644.470 305.690 ;
        RECT 644.240 305.310 644.490 305.400 ;
        RECT 626.860 304.880 627.410 304.970 ;
        RECT 614.860 304.510 615.030 304.680 ;
        RECT 616.470 304.510 616.640 304.680 ;
        RECT 625.360 304.570 627.410 304.880 ;
        RECT 625.360 304.510 626.280 304.570 ;
        RECT 605.280 303.360 605.750 304.410 ;
        RECT 614.800 304.370 616.660 304.510 ;
        RECT 615.550 303.360 615.890 304.370 ;
        RECT 625.550 303.360 626.020 304.510 ;
        RECT 626.860 304.430 627.410 304.570 ;
        RECT 640.230 303.370 640.410 305.260 ;
        RECT 644.250 303.370 644.490 305.310 ;
        RECT 646.060 303.370 649.270 303.990 ;
        RECT 631.870 303.360 643.420 303.370 ;
        RECT 643.660 303.360 649.270 303.370 ;
        RECT 600.180 302.200 649.270 303.360 ;
        RECT 631.870 302.170 649.270 302.200 ;
        RECT 646.060 301.600 649.270 302.170 ;
        RECT 677.010 298.860 677.400 316.140 ;
        RECT 686.470 316.100 689.420 316.205 ;
        RECT 691.300 316.150 694.250 316.205 ;
        RECT 695.670 316.050 698.240 316.205 ;
        RECT 695.670 315.990 698.220 316.050 ;
        RECT 851.510 315.680 852.180 327.420 ;
        RECT 853.880 327.250 854.150 327.630 ;
        RECT 853.900 326.160 854.150 327.250 ;
        RECT 853.880 325.780 854.150 326.160 ;
        RECT 853.900 324.690 854.150 325.780 ;
        RECT 853.880 324.310 854.150 324.690 ;
        RECT 853.900 323.220 854.150 324.310 ;
        RECT 853.880 322.840 854.150 323.220 ;
        RECT 853.900 321.750 854.150 322.840 ;
        RECT 853.880 321.370 854.150 321.750 ;
        RECT 853.900 320.280 854.150 321.370 ;
        RECT 874.480 320.550 874.710 320.780 ;
        RECT 853.880 319.900 854.150 320.280 ;
        RECT 853.900 318.810 854.150 319.900 ;
        RECT 853.880 318.430 854.150 318.810 ;
        RECT 853.900 317.340 854.150 318.430 ;
        RECT 853.880 316.960 854.150 317.340 ;
        RECT 853.900 315.870 854.150 316.960 ;
        RECT 851.640 312.970 851.980 315.680 ;
        RECT 853.880 315.490 854.150 315.870 ;
        RECT 853.900 314.400 854.150 315.490 ;
        RECT 874.470 314.930 874.720 320.550 ;
        RECT 876.590 316.360 877.440 320.440 ;
        RECT 853.880 314.330 854.150 314.400 ;
        RECT 853.870 314.210 854.150 314.330 ;
        RECT 874.430 314.660 874.720 314.930 ;
        RECT 874.430 314.520 874.710 314.660 ;
        RECT 876.560 314.620 877.440 316.360 ;
        RECT 853.870 314.020 854.110 314.210 ;
        RECT 853.870 312.970 854.090 314.020 ;
        RECT 874.430 312.970 874.690 314.520 ;
        RECT 876.560 312.970 877.370 314.620 ;
        RECT 851.640 310.890 877.810 312.970 ;
        RECT 796.480 304.490 811.840 304.655 ;
        RECT 814.240 304.490 829.600 304.655 ;
        RECT 796.480 304.470 829.600 304.490 ;
        RECT 831.780 304.470 833.220 304.625 ;
        RECT 835.420 304.490 840.700 304.685 ;
        RECT 842.690 304.490 844.130 304.685 ;
        RECT 835.420 304.470 844.130 304.490 ;
        RECT 796.480 304.315 844.130 304.470 ;
        RECT 796.480 304.285 836.240 304.315 ;
        RECT 810.940 304.145 814.700 304.285 ;
        RECT 828.490 304.175 836.240 304.285 ;
        RECT 840.440 304.175 844.110 304.315 ;
        RECT 828.490 304.145 844.130 304.175 ;
        RECT 796.480 304.030 844.130 304.145 ;
        RECT 796.480 303.970 840.700 304.030 ;
        RECT 796.480 303.915 811.840 303.970 ;
        RECT 814.240 303.950 840.700 303.970 ;
        RECT 814.240 303.915 829.600 303.950 ;
        RECT 831.780 303.885 833.220 303.950 ;
        RECT 835.420 303.945 840.700 303.950 ;
        RECT 842.690 303.945 844.130 304.030 ;
        RECT 669.220 296.820 669.930 296.880 ;
        RECT 676.970 296.820 677.440 298.860 ;
        RECT 669.220 296.800 677.440 296.820 ;
        RECT 669.220 296.060 677.400 296.800 ;
        RECT 635.060 290.065 636.500 290.435 ;
        RECT 639.250 290.155 640.690 290.525 ;
        RECT 595.170 289.615 596.610 289.985 ;
        RECT 635.190 289.925 635.370 290.065 ;
        RECT 639.350 290.015 639.490 290.155 ;
        RECT 643.350 290.135 644.790 290.505 ;
        RECT 635.060 289.900 636.500 289.925 ;
        RECT 639.250 289.900 640.690 290.015 ;
        RECT 643.770 289.995 644.010 290.135 ;
        RECT 643.350 289.950 644.790 289.995 ;
        RECT 645.730 289.950 646.380 291.070 ;
        RECT 635.060 289.890 642.980 289.900 ;
        RECT 643.350 289.890 646.380 289.950 ;
        RECT 596.410 289.475 596.550 289.615 ;
        RECT 595.170 289.245 596.610 289.475 ;
        RECT 596.410 288.820 596.550 289.245 ;
        RECT 596.350 288.460 597.040 288.820 ;
        RECT 118.110 287.200 119.090 287.430 ;
        RECT 121.580 287.200 122.560 287.430 ;
        RECT 125.050 287.200 126.030 287.430 ;
        RECT 128.520 287.200 129.500 287.430 ;
        RECT 131.990 287.200 132.970 287.430 ;
        RECT 135.460 287.200 136.440 287.430 ;
        RECT 138.930 287.200 139.910 287.430 ;
        RECT 142.400 287.200 143.380 287.430 ;
        RECT 145.870 287.200 146.850 287.430 ;
        RECT 149.340 287.200 150.320 287.430 ;
        RECT 605.130 285.230 606.020 289.700 ;
        RECT 614.790 286.970 615.020 287.350 ;
        RECT 616.370 286.970 616.600 287.350 ;
        RECT 614.810 285.880 614.970 286.970 ;
        RECT 616.390 285.880 616.550 286.970 ;
        RECT 614.790 285.500 615.020 285.880 ;
        RECT 616.370 285.500 616.600 285.880 ;
        RECT 625.310 285.700 626.230 289.830 ;
        RECT 635.060 289.785 646.380 289.890 ;
        RECT 635.060 289.695 639.550 289.785 ;
        RECT 635.110 289.100 635.340 289.695 ;
        RECT 636.240 289.680 639.550 289.695 ;
        RECT 640.450 289.760 646.380 289.785 ;
        RECT 640.450 289.720 646.000 289.760 ;
        RECT 640.450 289.680 645.160 289.720 ;
        RECT 642.950 289.670 644.520 289.680 ;
        RECT 634.880 288.750 635.380 289.100 ;
        RECT 640.140 286.080 640.370 286.460 ;
        RECT 644.190 286.220 644.420 286.510 ;
        RECT 644.190 286.130 644.440 286.220 ;
        RECT 626.810 285.700 627.360 285.790 ;
        RECT 614.810 285.330 614.980 285.500 ;
        RECT 616.420 285.330 616.590 285.500 ;
        RECT 625.310 285.390 627.360 285.700 ;
        RECT 625.310 285.330 626.230 285.390 ;
        RECT 118.110 283.910 119.090 284.140 ;
        RECT 121.580 283.910 122.560 284.140 ;
        RECT 125.050 283.910 126.030 284.140 ;
        RECT 128.520 283.910 129.500 284.140 ;
        RECT 131.990 283.910 132.970 284.140 ;
        RECT 135.460 283.910 136.440 284.140 ;
        RECT 138.930 283.910 139.910 284.140 ;
        RECT 142.400 283.910 143.380 284.140 ;
        RECT 145.870 283.910 146.850 284.140 ;
        RECT 149.340 283.910 150.320 284.140 ;
        RECT 151.610 283.750 152.080 284.350 ;
        RECT 605.230 284.180 605.700 285.230 ;
        RECT 614.750 285.190 616.610 285.330 ;
        RECT 615.500 284.180 615.840 285.190 ;
        RECT 625.500 284.180 625.970 285.330 ;
        RECT 626.810 285.250 627.360 285.390 ;
        RECT 640.180 284.190 640.360 286.080 ;
        RECT 644.200 284.190 644.440 286.130 ;
        RECT 645.860 284.190 649.070 284.900 ;
        RECT 631.820 284.180 643.370 284.190 ;
        RECT 643.610 284.180 649.070 284.190 ;
        RECT 600.130 283.020 649.070 284.180 ;
        RECT 631.820 282.990 649.070 283.020 ;
        RECT 645.860 282.510 649.070 282.990 ;
        RECT 118.110 280.620 119.090 280.850 ;
        RECT 121.580 280.620 122.560 280.850 ;
        RECT 125.050 280.620 126.030 280.850 ;
        RECT 128.520 280.620 129.500 280.850 ;
        RECT 131.990 280.620 132.970 280.850 ;
        RECT 135.460 280.620 136.440 280.850 ;
        RECT 138.930 280.620 139.910 280.850 ;
        RECT 142.400 280.620 143.380 280.850 ;
        RECT 145.870 280.620 146.850 280.850 ;
        RECT 149.340 280.620 150.320 280.850 ;
        RECT 121.370 278.660 125.810 279.540 ;
        RECT 143.430 279.240 147.880 279.950 ;
        RECT 114.580 274.300 116.010 276.880 ;
        RECT 118.140 274.460 119.120 274.690 ;
        RECT 121.610 274.460 122.590 274.690 ;
        RECT 125.080 274.460 126.060 274.690 ;
        RECT 128.550 274.460 129.530 274.690 ;
        RECT 132.020 274.460 133.000 274.690 ;
        RECT 135.490 274.460 136.470 274.690 ;
        RECT 138.960 274.460 139.940 274.690 ;
        RECT 142.430 274.460 143.410 274.690 ;
        RECT 145.900 274.460 146.880 274.690 ;
        RECT 149.370 274.460 150.350 274.690 ;
        RECT 634.980 271.595 636.420 271.965 ;
        RECT 639.170 271.685 640.610 272.055 ;
        RECT 595.090 271.145 596.530 271.515 ;
        RECT 635.110 271.455 635.290 271.595 ;
        RECT 639.270 271.545 639.410 271.685 ;
        RECT 643.270 271.665 644.710 272.035 ;
        RECT 634.980 271.430 636.420 271.455 ;
        RECT 639.170 271.430 640.610 271.545 ;
        RECT 643.690 271.525 643.930 271.665 ;
        RECT 643.270 271.430 644.710 271.525 ;
        RECT 645.850 271.470 646.500 272.630 ;
        RECT 644.930 271.430 646.500 271.470 ;
        RECT 634.980 271.420 642.900 271.430 ;
        RECT 643.270 271.420 646.500 271.430 ;
        RECT 596.330 271.005 596.470 271.145 ;
        RECT 595.090 270.775 596.530 271.005 ;
        RECT 121.400 269.210 125.840 270.090 ;
        RECT 143.460 269.790 147.910 270.500 ;
        RECT 596.330 270.350 596.470 270.775 ;
        RECT 596.270 269.990 596.960 270.350 ;
        RECT 118.220 268.040 119.200 268.270 ;
        RECT 121.690 268.040 122.670 268.270 ;
        RECT 125.160 268.040 126.140 268.270 ;
        RECT 128.630 268.040 129.610 268.270 ;
        RECT 132.100 268.040 133.080 268.270 ;
        RECT 135.570 268.040 136.550 268.270 ;
        RECT 139.040 268.040 140.020 268.270 ;
        RECT 142.510 268.040 143.490 268.270 ;
        RECT 145.980 268.040 146.960 268.270 ;
        RECT 149.450 268.040 150.430 268.270 ;
        RECT 605.050 266.760 605.940 271.230 ;
        RECT 614.710 268.500 614.940 268.880 ;
        RECT 616.290 268.500 616.520 268.880 ;
        RECT 614.730 267.410 614.890 268.500 ;
        RECT 616.310 267.410 616.470 268.500 ;
        RECT 614.710 267.030 614.940 267.410 ;
        RECT 616.290 267.030 616.520 267.410 ;
        RECT 625.230 267.230 626.150 271.360 ;
        RECT 634.980 271.320 646.500 271.420 ;
        RECT 634.980 271.315 646.030 271.320 ;
        RECT 634.980 271.225 639.470 271.315 ;
        RECT 635.030 270.630 635.260 271.225 ;
        RECT 636.160 271.210 639.470 271.225 ;
        RECT 640.370 271.240 646.030 271.315 ;
        RECT 640.370 271.210 645.080 271.240 ;
        RECT 642.870 271.200 644.440 271.210 ;
        RECT 634.800 270.280 635.300 270.630 ;
        RECT 640.060 267.610 640.290 267.990 ;
        RECT 644.110 267.750 644.340 268.040 ;
        RECT 644.110 267.660 644.360 267.750 ;
        RECT 626.730 267.230 627.280 267.320 ;
        RECT 614.730 266.860 614.900 267.030 ;
        RECT 616.340 266.860 616.510 267.030 ;
        RECT 625.230 266.920 627.280 267.230 ;
        RECT 625.230 266.860 626.150 266.920 ;
        RECT 605.150 265.710 605.620 266.760 ;
        RECT 614.670 266.720 616.530 266.860 ;
        RECT 615.420 265.710 615.760 266.720 ;
        RECT 625.420 265.710 625.890 266.860 ;
        RECT 626.730 266.780 627.280 266.920 ;
        RECT 640.100 265.720 640.280 267.610 ;
        RECT 644.120 265.720 644.360 267.660 ;
        RECT 669.220 267.330 669.930 296.060 ;
        RECT 677.010 295.100 677.400 296.060 ;
        RECT 680.060 295.480 695.420 295.595 ;
        RECT 697.550 295.480 712.910 295.555 ;
        RECT 680.060 295.410 712.910 295.480 ;
        RECT 715.160 295.470 730.520 295.615 ;
        RECT 732.860 295.470 748.220 295.565 ;
        RECT 715.160 295.450 748.220 295.470 ;
        RECT 750.600 295.450 765.960 295.555 ;
        RECT 715.160 295.410 765.960 295.450 ;
        RECT 680.060 295.245 765.960 295.410 ;
        RECT 680.060 295.225 716.080 295.245 ;
        RECT 694.060 295.185 716.080 295.225 ;
        RECT 677.010 295.030 679.860 295.100 ;
        RECT 694.060 295.085 698.310 295.185 ;
        RECT 680.060 295.045 698.310 295.085 ;
        RECT 711.830 295.105 716.080 295.185 ;
        RECT 729.560 295.195 765.960 295.245 ;
        RECT 729.560 295.105 733.810 295.195 ;
        RECT 711.830 295.055 733.810 295.105 ;
        RECT 746.990 295.185 765.960 295.195 ;
        RECT 746.990 295.055 751.240 295.185 ;
        RECT 711.830 295.045 751.240 295.055 ;
        RECT 680.060 295.030 765.960 295.045 ;
        RECT 677.010 294.960 765.960 295.030 ;
        RECT 677.010 294.890 695.420 294.960 ;
        RECT 677.010 294.760 679.860 294.890 ;
        RECT 680.060 294.855 695.420 294.890 ;
        RECT 697.550 294.950 765.960 294.960 ;
        RECT 697.550 294.890 730.520 294.950 ;
        RECT 697.550 294.815 712.910 294.890 ;
        RECT 715.160 294.875 730.520 294.890 ;
        RECT 732.860 294.930 765.960 294.950 ;
        RECT 732.860 294.825 748.220 294.930 ;
        RECT 750.600 294.815 765.960 294.930 ;
        RECT 855.800 294.545 859.160 294.915 ;
        RECT 857.650 294.405 858.360 294.545 ;
        RECT 855.800 294.175 859.160 294.405 ;
        RECT 839.390 292.565 842.750 292.935 ;
        RECT 839.570 292.425 840.230 292.565 ;
        RECT 841.440 292.425 841.660 292.565 ;
        RECT 839.390 292.195 842.750 292.425 ;
        RECT 845.090 290.915 848.450 291.285 ;
        RECT 847.260 290.775 847.480 290.915 ;
        RECT 861.180 290.830 864.540 291.015 ;
        RECT 870.170 290.830 870.770 310.890 ;
        RECT 845.090 290.700 848.450 290.775 ;
        RECT 845.090 290.680 851.120 290.700 ;
        RECT 845.090 290.545 851.210 290.680 ;
        RECT 861.180 290.645 870.770 290.830 ;
        RECT 818.940 289.555 822.300 289.925 ;
        RECT 820.620 289.415 822.020 289.555 ;
        RECT 818.940 289.185 822.300 289.415 ;
        RECT 824.390 287.385 827.750 287.755 ;
        RECT 829.930 287.405 835.210 287.775 ;
        RECT 839.400 287.445 842.760 287.815 ;
        RECT 824.700 287.245 825.860 287.385 ;
        RECT 831.950 287.265 832.170 287.405 ;
        RECT 833.900 287.265 834.120 287.405 ;
        RECT 839.600 287.305 840.260 287.445 ;
        RECT 841.390 287.305 841.610 287.445 ;
        RECT 845.210 287.440 845.480 290.545 ;
        RECT 848.120 290.340 851.210 290.545 ;
        RECT 861.990 290.505 862.650 290.645 ;
        RECT 864.270 290.505 870.770 290.645 ;
        RECT 850.870 288.760 851.210 290.340 ;
        RECT 861.180 290.470 870.770 290.505 ;
        RECT 861.180 290.430 870.760 290.470 ;
        RECT 861.180 290.275 864.540 290.430 ;
        RECT 855.840 289.015 859.200 289.385 ;
        RECT 857.590 288.875 858.500 289.015 ;
        RECT 855.840 288.760 859.200 288.875 ;
        RECT 850.870 288.645 859.200 288.760 ;
        RECT 850.870 288.390 856.170 288.645 ;
        RECT 850.870 288.370 851.750 288.390 ;
        RECT 824.390 287.180 827.750 287.245 ;
        RECT 829.930 287.210 835.210 287.265 ;
        RECT 839.400 287.240 842.760 287.305 ;
        RECT 844.610 287.240 845.480 287.440 ;
        RECT 839.400 287.210 845.500 287.240 ;
        RECT 829.930 287.180 845.500 287.210 ;
        RECT 824.390 287.075 845.500 287.180 ;
        RECT 824.390 287.035 839.650 287.075 ;
        RECT 824.390 287.015 830.880 287.035 ;
        RECT 827.500 286.870 830.880 287.015 ;
        RECT 835.100 286.890 839.650 287.035 ;
        RECT 842.500 286.970 845.500 287.075 ;
        RECT 844.610 286.650 845.380 286.970 ;
        RECT 818.910 284.395 822.270 284.765 ;
        RECT 821.560 284.255 822.130 284.395 ;
        RECT 818.910 284.025 822.270 284.255 ;
        RECT 855.910 283.615 859.270 283.985 ;
        RECT 857.560 283.475 858.130 283.615 ;
        RECT 855.910 283.245 859.270 283.475 ;
        RECT 861.260 281.595 864.620 281.965 ;
        RECT 861.920 281.455 862.720 281.595 ;
        RECT 861.260 281.225 864.620 281.455 ;
        RECT 799.530 279.930 800.970 280.075 ;
        RECT 799.250 279.705 800.970 279.930 ;
        RECT 799.250 279.565 799.870 279.705 ;
        RECT 799.250 279.335 800.970 279.565 ;
        RECT 819.350 279.365 824.630 279.735 ;
        RECT 799.250 279.240 799.870 279.335 ;
        RECT 821.640 279.225 822.210 279.365 ;
        RECT 827.960 279.275 831.320 279.645 ;
        RECT 833.250 279.275 838.530 279.645 ;
        RECT 840.460 279.275 844.300 279.645 ;
        RECT 819.350 279.100 824.630 279.225 ;
        RECT 829.570 279.135 829.750 279.275 ;
        RECT 834.870 279.135 835.050 279.275 ;
        RECT 842.870 279.135 843.090 279.275 ;
        RECT 827.960 279.100 831.320 279.135 ;
        RECT 819.350 279.070 831.320 279.100 ;
        RECT 833.250 279.070 838.530 279.135 ;
        RECT 819.350 278.995 838.530 279.070 ;
        RECT 824.310 278.905 838.530 278.995 ;
        RECT 840.460 279.010 844.300 279.135 ;
        RECT 845.040 279.010 845.610 279.390 ;
        RECT 846.300 279.275 851.580 279.645 ;
        RECT 848.280 279.135 848.500 279.275 ;
        RECT 846.300 279.010 851.580 279.135 ;
        RECT 840.460 278.905 851.580 279.010 ;
        RECT 824.310 278.890 828.220 278.905 ;
        RECT 679.390 278.485 684.670 278.855 ;
        RECT 696.670 278.495 701.950 278.865 ;
        RECT 714.440 278.495 719.720 278.865 ;
        RECT 731.680 278.495 736.960 278.865 ;
        RECT 749.160 278.505 754.440 278.875 ;
        RECT 831.070 278.860 834.980 278.905 ;
        RECT 844.030 278.740 846.530 278.905 ;
        RECT 682.530 278.345 682.710 278.485 ;
        RECT 679.390 278.270 684.670 278.345 ;
        RECT 694.480 278.270 695.160 278.460 ;
        RECT 698.000 278.355 698.180 278.495 ;
        RECT 699.550 278.355 699.850 278.495 ;
        RECT 717.180 278.355 717.480 278.495 ;
        RECT 733.380 278.355 733.640 278.495 ;
        RECT 751.490 278.365 751.770 278.505 ;
        RECT 696.670 278.270 701.950 278.355 ;
        RECT 679.390 278.240 701.950 278.270 ;
        RECT 714.440 278.250 719.720 278.355 ;
        RECT 731.680 278.250 736.960 278.355 ;
        RECT 714.440 278.240 736.960 278.250 ;
        RECT 679.390 278.220 736.960 278.240 ;
        RECT 749.160 278.220 754.440 278.365 ;
        RECT 679.390 278.135 754.440 278.220 ;
        RECT 855.930 278.155 859.290 278.525 ;
        RECT 679.390 278.125 749.500 278.135 ;
        RECT 679.390 278.115 697.140 278.125 ;
        RECT 684.300 278.000 697.140 278.115 ;
        RECT 694.480 277.680 695.160 278.000 ;
        RECT 701.680 277.970 714.520 278.125 ;
        RECT 719.400 277.980 732.240 278.125 ;
        RECT 736.660 277.950 749.500 278.125 ;
        RECT 857.630 278.015 858.360 278.155 ;
        RECT 855.930 277.785 859.290 278.015 ;
        RECT 748.150 274.870 748.370 274.880 ;
        RECT 748.140 274.860 749.090 274.870 ;
        RECT 749.570 274.860 750.130 275.100 ;
        RECT 751.620 274.860 751.880 274.990 ;
        RECT 748.140 274.690 751.880 274.860 ;
        RECT 748.140 274.670 749.090 274.690 ;
        RECT 748.140 274.640 748.750 274.670 ;
        RECT 679.800 272.825 685.080 273.195 ;
        RECT 682.310 272.685 682.550 272.825 ;
        RECT 687.040 272.785 692.320 273.155 ;
        RECT 679.800 272.530 685.080 272.685 ;
        RECT 688.720 272.645 690.160 272.785 ;
        RECT 687.040 272.610 692.320 272.645 ;
        RECT 694.710 272.610 695.390 273.060 ;
        RECT 697.030 272.845 702.310 273.215 ;
        RECT 699.540 272.705 699.780 272.845 ;
        RECT 704.270 272.805 709.550 273.175 ;
        RECT 714.600 272.945 719.880 273.315 ;
        RECT 717.110 272.805 717.350 272.945 ;
        RECT 721.840 272.905 727.120 273.275 ;
        RECT 731.770 272.975 737.050 273.345 ;
        RECT 697.030 272.610 702.310 272.705 ;
        RECT 705.950 272.665 707.390 272.805 ;
        RECT 714.600 272.680 719.880 272.805 ;
        RECT 723.520 272.765 724.960 272.905 ;
        RECT 734.280 272.835 734.520 272.975 ;
        RECT 739.010 272.935 744.290 273.305 ;
        RECT 687.040 272.550 702.310 272.610 ;
        RECT 704.270 272.620 709.550 272.665 ;
        RECT 709.690 272.650 719.880 272.680 ;
        RECT 721.840 272.740 727.120 272.765 ;
        RECT 731.770 272.740 737.050 272.835 ;
        RECT 740.690 272.795 742.130 272.935 ;
        RECT 748.150 272.800 748.370 274.640 ;
        RECT 749.570 274.600 750.130 274.690 ;
        RECT 751.620 274.620 751.880 274.690 ;
        RECT 798.800 274.250 799.570 274.940 ;
        RECT 749.580 273.035 754.860 273.405 ;
        RECT 752.090 272.895 752.330 273.035 ;
        RECT 756.820 272.995 762.100 273.365 ;
        RECT 749.580 272.800 754.860 272.895 ;
        RECT 758.500 272.855 759.940 272.995 ;
        RECT 721.840 272.680 737.050 272.740 ;
        RECT 739.010 272.730 744.290 272.795 ;
        RECT 744.440 272.740 754.860 272.800 ;
        RECT 756.820 272.740 762.100 272.855 ;
        RECT 744.440 272.730 762.100 272.740 ;
        RECT 739.010 272.680 762.100 272.730 ;
        RECT 721.840 272.665 762.100 272.680 ;
        RECT 721.840 272.650 749.740 272.665 ;
        RECT 709.690 272.620 749.740 272.650 ;
        RECT 704.270 272.605 749.740 272.620 ;
        RECT 704.270 272.575 731.950 272.605 ;
        RECT 704.270 272.550 714.710 272.575 ;
        RECT 687.040 272.530 714.710 272.550 ;
        RECT 679.800 272.475 714.710 272.530 ;
        RECT 679.800 272.455 697.220 272.475 ;
        RECT 684.500 272.415 697.220 272.455 ;
        RECT 684.500 272.340 687.440 272.415 ;
        RECT 691.940 272.260 697.220 272.415 ;
        RECT 701.730 272.435 714.710 272.475 ;
        RECT 719.300 272.535 731.950 272.575 ;
        RECT 719.300 272.460 722.240 272.535 ;
        RECT 726.790 272.500 731.950 272.535 ;
        RECT 736.470 272.565 749.740 272.605 ;
        RECT 736.470 272.490 739.410 272.565 ;
        RECT 701.730 272.360 704.670 272.435 ;
        RECT 709.370 272.390 714.710 272.435 ;
        RECT 743.990 272.410 749.740 272.565 ;
        RECT 754.280 272.625 762.100 272.665 ;
        RECT 754.280 272.550 757.220 272.625 ;
        RECT 748.150 272.400 748.370 272.410 ;
        RECT 780.960 271.665 796.320 272.035 ;
        RECT 794.950 271.525 795.190 271.665 ;
        RECT 780.960 271.380 796.320 271.525 ;
        RECT 799.040 271.380 799.300 274.250 ;
        RECT 799.850 271.655 815.210 272.025 ;
        RECT 813.920 271.515 814.160 271.655 ;
        RECT 818.700 271.625 834.060 271.995 ;
        RECT 838.420 271.665 842.260 272.035 ;
        RECT 799.850 271.380 815.210 271.515 ;
        RECT 821.240 271.485 821.480 271.625 ;
        RECT 841.430 271.525 841.610 271.665 ;
        RECT 855.930 271.615 859.290 271.985 ;
        RECT 818.700 271.410 834.060 271.485 ;
        RECT 838.420 271.410 842.260 271.525 ;
        RECT 857.580 271.475 858.160 271.615 ;
        RECT 818.700 271.380 842.260 271.410 ;
        RECT 780.960 271.295 842.260 271.380 ;
        RECT 796.010 271.285 838.660 271.295 ;
        RECT 796.010 271.200 800.110 271.285 ;
        RECT 814.910 271.255 838.660 271.285 ;
        RECT 814.910 271.200 819.010 271.255 ;
        RECT 749.760 268.430 750.270 268.870 ;
        RECT 749.830 268.410 750.190 268.430 ;
        RECT 679.920 267.390 683.280 267.515 ;
        RECT 674.600 267.330 683.280 267.390 ;
        RECT 669.220 267.145 683.280 267.330 ;
        RECT 685.580 267.155 688.940 267.525 ;
        RECT 690.930 267.175 694.290 267.545 ;
        RECT 669.220 267.005 681.430 267.145 ;
        RECT 687.240 267.015 687.500 267.155 ;
        RECT 669.220 266.900 683.280 267.005 ;
        RECT 685.580 266.960 688.940 267.015 ;
        RECT 689.750 266.960 690.430 267.150 ;
        RECT 692.430 267.035 692.670 267.175 ;
        RECT 697.150 267.165 700.510 267.535 ;
        RECT 702.810 267.175 706.170 267.545 ;
        RECT 708.160 267.195 711.520 267.565 ;
        RECT 714.720 267.265 718.080 267.635 ;
        RECT 720.380 267.275 723.740 267.645 ;
        RECT 725.730 267.295 729.090 267.665 ;
        RECT 731.890 267.295 735.250 267.665 ;
        RECT 737.550 267.305 740.910 267.675 ;
        RECT 742.900 267.325 746.260 267.695 ;
        RECT 749.700 267.355 753.060 267.725 ;
        RECT 755.360 267.365 758.720 267.735 ;
        RECT 760.710 267.600 764.070 267.755 ;
        RECT 760.710 267.385 764.220 267.600 ;
        RECT 690.930 267.000 694.290 267.035 ;
        RECT 698.410 267.025 698.660 267.165 ;
        RECT 704.470 267.035 704.730 267.175 ;
        RECT 697.150 267.000 700.510 267.025 ;
        RECT 690.930 266.960 700.510 267.000 ;
        RECT 685.580 266.920 700.510 266.960 ;
        RECT 702.810 266.980 706.170 267.035 ;
        RECT 706.980 266.980 707.660 267.170 ;
        RECT 709.660 267.055 709.900 267.195 ;
        RECT 715.980 267.125 716.230 267.265 ;
        RECT 722.040 267.135 722.300 267.275 ;
        RECT 708.160 267.030 711.520 267.055 ;
        RECT 714.720 267.030 718.080 267.125 ;
        RECT 708.160 267.020 718.080 267.030 ;
        RECT 720.380 267.080 723.740 267.135 ;
        RECT 724.550 267.080 725.230 267.270 ;
        RECT 727.230 267.155 727.470 267.295 ;
        RECT 733.150 267.155 733.400 267.295 ;
        RECT 739.210 267.165 739.470 267.305 ;
        RECT 725.730 267.080 729.090 267.155 ;
        RECT 720.380 267.020 729.090 267.080 ;
        RECT 708.160 267.010 729.090 267.020 ;
        RECT 731.890 267.050 735.250 267.155 ;
        RECT 737.550 267.110 740.910 267.165 ;
        RECT 741.720 267.110 742.400 267.300 ;
        RECT 744.400 267.185 744.640 267.325 ;
        RECT 750.960 267.215 751.210 267.355 ;
        RECT 757.020 267.225 757.280 267.365 ;
        RECT 742.900 267.130 746.260 267.185 ;
        RECT 749.700 267.130 753.060 267.215 ;
        RECT 742.900 267.110 753.060 267.130 ;
        RECT 755.360 267.170 758.720 267.225 ;
        RECT 759.530 267.170 760.210 267.360 ;
        RECT 762.210 267.245 762.450 267.385 ;
        RECT 763.620 267.245 764.220 267.385 ;
        RECT 760.710 267.170 764.220 267.245 ;
        RECT 755.360 267.110 764.220 267.170 ;
        RECT 737.550 267.050 764.220 267.110 ;
        RECT 731.890 267.015 764.070 267.050 ;
        RECT 731.890 267.010 761.170 267.015 ;
        RECT 708.160 266.995 761.170 267.010 ;
        RECT 708.160 266.985 755.510 266.995 ;
        RECT 708.160 266.980 750.000 266.985 ;
        RECT 702.810 266.955 750.000 266.980 ;
        RECT 702.810 266.935 743.360 266.955 ;
        RECT 702.810 266.925 737.700 266.935 ;
        RECT 702.810 266.920 726.190 266.925 ;
        RECT 685.580 266.905 726.190 266.920 ;
        RECT 685.580 266.900 720.530 266.905 ;
        RECT 669.220 266.895 720.530 266.900 ;
        RECT 669.220 266.825 714.830 266.895 ;
        RECT 717.590 266.830 720.530 266.895 ;
        RECT 723.250 266.890 726.190 266.905 ;
        RECT 669.220 266.805 708.620 266.825 ;
        RECT 669.220 266.800 691.390 266.805 ;
        RECT 669.220 266.740 675.000 266.800 ;
        RECT 679.920 266.785 691.390 266.800 ;
        RECT 679.920 266.775 685.730 266.785 ;
        RECT 682.790 266.710 685.730 266.775 ;
        RECT 688.450 266.770 691.390 266.785 ;
        RECT 693.830 266.795 702.960 266.805 ;
        RECT 689.750 266.610 690.430 266.770 ;
        RECT 693.830 266.690 697.260 266.795 ;
        RECT 700.020 266.730 702.960 266.795 ;
        RECT 705.680 266.790 708.620 266.805 ;
        RECT 706.980 266.630 707.660 266.790 ;
        RECT 711.400 266.720 714.830 266.825 ;
        RECT 724.550 266.730 725.230 266.890 ;
        RECT 728.890 266.800 732.790 266.925 ;
        RECT 734.760 266.860 737.700 266.925 ;
        RECT 740.420 266.920 743.360 266.935 ;
        RECT 746.100 266.920 750.000 266.955 ;
        RECT 752.570 266.920 755.510 266.985 ;
        RECT 758.230 266.980 761.170 266.995 ;
        RECT 741.720 266.760 742.400 266.920 ;
        RECT 759.530 266.820 760.210 266.980 ;
        RECT 645.900 265.720 649.110 266.210 ;
        RECT 631.740 265.710 643.290 265.720 ;
        RECT 643.530 265.710 649.110 265.720 ;
        RECT 118.220 264.750 119.200 264.980 ;
        RECT 121.690 264.750 122.670 264.980 ;
        RECT 125.160 264.750 126.140 264.980 ;
        RECT 128.630 264.750 129.610 264.980 ;
        RECT 132.100 264.750 133.080 264.980 ;
        RECT 135.570 264.750 136.550 264.980 ;
        RECT 139.040 264.750 140.020 264.980 ;
        RECT 142.510 264.750 143.490 264.980 ;
        RECT 145.980 264.750 146.960 264.980 ;
        RECT 149.450 264.750 150.430 264.980 ;
        RECT 151.800 264.460 152.550 265.530 ;
        RECT 600.050 264.550 649.110 265.710 ;
        RECT 631.740 264.520 649.110 264.550 ;
        RECT 645.900 263.820 649.110 264.520 ;
        RECT 780.970 264.390 796.330 264.475 ;
        RECT 780.680 264.105 796.330 264.390 ;
        RECT 799.500 264.165 814.860 264.535 ;
        RECT 780.680 263.965 781.430 264.105 ;
        RECT 792.120 263.965 792.360 264.105 ;
        RECT 813.530 264.025 813.770 264.165 ;
        RECT 799.500 263.990 814.860 264.025 ;
        RECT 818.220 263.990 818.550 271.200 ;
        RECT 833.830 271.190 838.660 271.255 ;
        RECT 855.930 271.245 859.290 271.475 ;
        RECT 835.200 265.870 835.600 271.190 ;
        RECT 844.670 269.405 848.030 269.775 ;
        RECT 850.080 269.415 851.520 269.785 ;
        RECT 846.720 269.265 846.910 269.405 ;
        RECT 850.280 269.275 850.470 269.415 ;
        RECT 844.670 269.230 848.030 269.265 ;
        RECT 850.080 269.230 851.520 269.275 ;
        RECT 844.670 269.090 851.520 269.230 ;
        RECT 844.670 269.035 848.030 269.090 ;
        RECT 850.080 269.045 851.520 269.090 ;
        RECT 838.430 266.105 841.790 266.475 ;
        RECT 845.570 266.200 845.850 269.035 ;
        RECT 861.250 268.225 864.610 268.595 ;
        RECT 861.900 268.085 863.500 268.225 ;
        RECT 861.250 267.855 864.610 268.085 ;
        RECT 840.480 265.965 840.660 266.105 ;
        RECT 838.430 265.870 841.790 265.965 ;
        RECT 835.200 265.840 841.790 265.870 ;
        RECT 845.140 265.840 846.240 266.200 ;
        RECT 835.200 265.735 846.240 265.840 ;
        RECT 835.200 265.650 840.030 265.735 ;
        RECT 841.400 265.640 846.240 265.735 ;
        RECT 845.140 265.160 846.240 265.640 ;
        RECT 856.010 264.945 859.370 265.315 ;
        RECT 857.560 264.805 858.590 264.945 ;
        RECT 856.010 264.575 859.370 264.805 ;
        RECT 780.680 263.930 796.330 263.965 ;
        RECT 799.500 263.930 818.550 263.990 ;
        RECT 780.680 263.810 818.550 263.930 ;
        RECT 780.680 263.795 814.860 263.810 ;
        RECT 780.680 263.750 799.790 263.795 ;
        RECT 818.220 263.790 818.550 263.810 ;
        RECT 780.680 263.735 796.330 263.750 ;
        RECT 780.680 263.700 781.430 263.735 ;
        RECT 118.220 261.460 119.200 261.690 ;
        RECT 121.690 261.460 122.670 261.690 ;
        RECT 125.160 261.460 126.140 261.690 ;
        RECT 128.630 261.460 129.610 261.690 ;
        RECT 132.100 261.460 133.080 261.690 ;
        RECT 135.570 261.460 136.550 261.690 ;
        RECT 139.040 261.460 140.020 261.690 ;
        RECT 142.510 261.460 143.490 261.690 ;
        RECT 145.980 261.460 146.960 261.690 ;
        RECT 149.450 261.460 150.430 261.690 ;
        RECT 121.480 259.500 125.920 260.380 ;
        RECT 143.540 260.080 147.990 260.790 ;
        RECT 682.170 258.790 682.620 258.850 ;
        RECT 699.470 258.790 699.920 258.900 ;
        RECT 717.260 258.790 717.710 258.940 ;
        RECT 734.520 258.790 734.970 258.970 ;
        RECT 751.990 258.880 752.440 258.960 ;
        RECT 756.330 258.880 756.990 259.030 ;
        RECT 751.990 258.790 756.990 258.880 ;
        RECT 682.170 258.700 756.990 258.790 ;
        RECT 682.170 258.650 752.440 258.700 ;
        RECT 682.170 258.510 682.620 258.650 ;
        RECT 679.370 256.955 684.650 257.325 ;
        RECT 682.510 256.815 682.690 256.955 ;
        RECT 679.370 256.740 684.650 256.815 ;
        RECT 691.320 256.740 691.730 258.650 ;
        RECT 699.470 258.560 699.920 258.650 ;
        RECT 717.260 258.600 717.710 258.650 ;
        RECT 734.520 258.630 734.970 258.650 ;
        RECT 751.990 258.620 752.440 258.650 ;
        RECT 756.330 258.420 756.990 258.700 ;
        RECT 696.650 256.965 701.930 257.335 ;
        RECT 714.420 256.965 719.700 257.335 ;
        RECT 731.660 256.965 736.940 257.335 ;
        RECT 749.140 256.975 754.420 257.345 ;
        RECT 694.460 256.740 695.140 256.930 ;
        RECT 697.980 256.825 698.160 256.965 ;
        RECT 699.530 256.825 699.830 256.965 ;
        RECT 717.160 256.825 717.460 256.965 ;
        RECT 733.360 256.825 733.620 256.965 ;
        RECT 751.470 256.835 751.750 256.975 ;
        RECT 696.650 256.740 701.930 256.825 ;
        RECT 679.370 256.710 701.930 256.740 ;
        RECT 714.420 256.720 719.700 256.825 ;
        RECT 731.660 256.720 736.940 256.825 ;
        RECT 714.420 256.710 736.940 256.720 ;
        RECT 679.370 256.690 736.940 256.710 ;
        RECT 749.140 256.690 754.420 256.835 ;
        RECT 679.370 256.605 754.420 256.690 ;
        RECT 679.370 256.595 749.480 256.605 ;
        RECT 679.370 256.585 697.120 256.595 ;
        RECT 684.280 256.470 697.120 256.585 ;
        RECT 694.460 256.150 695.140 256.470 ;
        RECT 701.660 256.440 714.500 256.595 ;
        RECT 719.380 256.450 732.220 256.595 ;
        RECT 736.640 256.420 749.480 256.595 ;
        RECT 855.880 255.635 859.240 256.005 ;
        RECT 857.520 255.495 858.120 255.635 ;
        RECT 855.880 255.265 859.240 255.495 ;
        RECT 634.830 253.865 636.270 254.235 ;
        RECT 639.020 253.955 640.460 254.325 ;
        RECT 594.940 253.415 596.380 253.785 ;
        RECT 634.960 253.725 635.140 253.865 ;
        RECT 639.120 253.815 639.260 253.955 ;
        RECT 643.120 253.935 644.560 254.305 ;
        RECT 634.830 253.700 636.270 253.725 ;
        RECT 639.020 253.700 640.460 253.815 ;
        RECT 643.540 253.795 643.780 253.935 ;
        RECT 643.120 253.700 644.560 253.795 ;
        RECT 645.650 253.710 646.300 254.940 ;
        RECT 644.790 253.700 646.300 253.710 ;
        RECT 634.830 253.690 642.750 253.700 ;
        RECT 643.120 253.690 646.300 253.700 ;
        RECT 634.830 253.630 646.300 253.690 ;
        RECT 596.180 253.275 596.320 253.415 ;
        RECT 594.940 253.045 596.380 253.275 ;
        RECT 596.180 252.620 596.320 253.045 ;
        RECT 596.120 252.260 596.810 252.620 ;
        RECT 604.900 249.030 605.790 253.500 ;
        RECT 614.560 250.770 614.790 251.150 ;
        RECT 616.140 250.770 616.370 251.150 ;
        RECT 614.580 249.680 614.740 250.770 ;
        RECT 616.160 249.680 616.320 250.770 ;
        RECT 614.560 249.300 614.790 249.680 ;
        RECT 616.140 249.300 616.370 249.680 ;
        RECT 625.080 249.500 626.000 253.630 ;
        RECT 634.830 253.585 645.850 253.630 ;
        RECT 634.830 253.495 639.320 253.585 ;
        RECT 634.880 252.900 635.110 253.495 ;
        RECT 636.010 253.480 639.320 253.495 ;
        RECT 640.220 253.540 645.850 253.585 ;
        RECT 640.220 253.480 644.930 253.540 ;
        RECT 642.720 253.470 644.290 253.480 ;
        RECT 678.770 253.120 679.190 253.130 ;
        RECT 679.770 253.120 680.330 253.360 ;
        RECT 748.400 253.330 749.070 253.340 ;
        RECT 749.550 253.330 750.110 253.570 ;
        RECT 751.600 253.330 751.860 253.460 ;
        RECT 681.820 253.120 682.080 253.250 ;
        RECT 678.770 253.110 682.080 253.120 ;
        RECT 678.710 252.950 682.080 253.110 ;
        RECT 678.710 252.910 679.190 252.950 ;
        RECT 634.650 252.550 635.150 252.900 ;
        RECT 678.710 252.820 679.000 252.910 ;
        RECT 679.770 252.860 680.330 252.950 ;
        RECT 681.820 252.880 682.080 252.950 ;
        RECT 748.400 253.160 751.860 253.330 ;
        RECT 748.400 253.140 749.070 253.160 ;
        RECT 678.710 252.400 678.980 252.820 ;
        RECT 678.710 251.410 679.000 252.400 ;
        RECT 679.780 251.410 685.060 251.665 ;
        RECT 678.710 251.295 685.060 251.410 ;
        RECT 678.710 251.155 680.210 251.295 ;
        RECT 682.290 251.155 682.530 251.295 ;
        RECT 687.020 251.255 692.300 251.625 ;
        RECT 678.710 251.010 685.060 251.155 ;
        RECT 688.700 251.115 690.140 251.255 ;
        RECT 679.780 251.000 685.060 251.010 ;
        RECT 687.020 251.080 692.300 251.115 ;
        RECT 694.690 251.080 695.370 251.530 ;
        RECT 697.010 251.315 702.290 251.685 ;
        RECT 699.520 251.175 699.760 251.315 ;
        RECT 704.250 251.275 709.530 251.645 ;
        RECT 714.580 251.415 719.860 251.785 ;
        RECT 717.090 251.275 717.330 251.415 ;
        RECT 721.820 251.375 727.100 251.745 ;
        RECT 731.750 251.445 737.030 251.815 ;
        RECT 697.010 251.080 702.290 251.175 ;
        RECT 705.930 251.135 707.370 251.275 ;
        RECT 714.580 251.150 719.860 251.275 ;
        RECT 723.500 251.235 724.940 251.375 ;
        RECT 734.260 251.305 734.500 251.445 ;
        RECT 738.990 251.405 744.270 251.775 ;
        RECT 687.020 251.020 702.290 251.080 ;
        RECT 704.250 251.090 709.530 251.135 ;
        RECT 709.670 251.120 719.860 251.150 ;
        RECT 721.820 251.210 727.100 251.235 ;
        RECT 730.510 251.210 730.780 251.290 ;
        RECT 731.750 251.210 737.030 251.305 ;
        RECT 740.670 251.265 742.110 251.405 ;
        RECT 748.400 251.270 748.670 253.140 ;
        RECT 749.550 253.070 750.110 253.160 ;
        RECT 751.600 253.090 751.860 253.160 ;
        RECT 861.190 253.145 864.550 253.515 ;
        RECT 756.280 252.840 756.870 252.940 ;
        RECT 760.260 252.840 760.500 253.060 ;
        RECT 861.940 253.005 862.670 253.145 ;
        RECT 756.140 252.710 760.500 252.840 ;
        RECT 861.190 252.775 864.550 253.005 ;
        RECT 756.140 252.650 760.470 252.710 ;
        RECT 756.280 252.120 756.870 252.650 ;
        RECT 749.560 251.505 754.840 251.875 ;
        RECT 752.070 251.365 752.310 251.505 ;
        RECT 756.800 251.465 762.080 251.835 ;
        RECT 749.560 251.270 754.840 251.365 ;
        RECT 758.480 251.325 759.920 251.465 ;
        RECT 721.820 251.150 737.030 251.210 ;
        RECT 738.990 251.200 744.270 251.265 ;
        RECT 744.420 251.210 754.840 251.270 ;
        RECT 756.800 251.210 762.080 251.325 ;
        RECT 744.420 251.200 762.080 251.210 ;
        RECT 738.990 251.150 762.080 251.200 ;
        RECT 721.820 251.135 762.080 251.150 ;
        RECT 721.820 251.120 749.720 251.135 ;
        RECT 709.670 251.090 749.720 251.120 ;
        RECT 704.250 251.075 749.720 251.090 ;
        RECT 704.250 251.045 731.930 251.075 ;
        RECT 704.250 251.020 714.690 251.045 ;
        RECT 687.020 251.000 714.690 251.020 ;
        RECT 679.780 250.945 714.690 251.000 ;
        RECT 679.780 250.925 697.200 250.945 ;
        RECT 684.480 250.885 697.200 250.925 ;
        RECT 684.480 250.810 687.420 250.885 ;
        RECT 691.920 250.730 697.200 250.885 ;
        RECT 701.710 250.905 714.690 250.945 ;
        RECT 719.280 251.005 731.930 251.045 ;
        RECT 719.280 250.930 722.220 251.005 ;
        RECT 726.770 250.970 731.930 251.005 ;
        RECT 736.450 251.035 749.720 251.075 ;
        RECT 736.450 250.960 739.390 251.035 ;
        RECT 701.710 250.830 704.650 250.905 ;
        RECT 709.350 250.860 714.690 250.905 ;
        RECT 743.970 250.880 749.720 251.035 ;
        RECT 754.260 251.095 762.080 251.135 ;
        RECT 754.260 251.020 757.200 251.095 ;
        RECT 639.910 249.880 640.140 250.260 ;
        RECT 643.960 250.020 644.190 250.310 ;
        RECT 643.960 249.930 644.210 250.020 ;
        RECT 626.580 249.500 627.130 249.590 ;
        RECT 614.580 249.130 614.750 249.300 ;
        RECT 616.190 249.130 616.360 249.300 ;
        RECT 625.080 249.190 627.130 249.500 ;
        RECT 625.080 249.130 626.000 249.190 ;
        RECT 601.550 248.380 602.610 248.820 ;
        RECT 605.000 247.980 605.470 249.030 ;
        RECT 614.520 248.990 616.380 249.130 ;
        RECT 615.270 247.980 615.610 248.990 ;
        RECT 625.270 247.980 625.740 249.130 ;
        RECT 626.580 249.050 627.130 249.190 ;
        RECT 639.950 247.990 640.130 249.880 ;
        RECT 643.970 247.990 644.210 249.930 ;
        RECT 855.940 249.865 859.300 250.235 ;
        RECT 857.490 249.725 858.270 249.865 ;
        RECT 855.940 249.630 859.300 249.725 ;
        RECT 861.600 249.630 861.900 252.775 ;
        RECT 855.940 249.495 861.900 249.630 ;
        RECT 859.150 249.410 861.900 249.495 ;
        RECT 859.150 249.380 861.850 249.410 ;
        RECT 645.980 247.990 649.190 248.480 ;
        RECT 631.590 247.980 643.140 247.990 ;
        RECT 643.380 247.980 649.190 247.990 ;
        RECT 591.480 246.060 591.730 247.355 ;
        RECT 599.900 246.820 649.190 247.980 ;
        RECT 591.130 244.660 592.380 246.060 ;
        RECT 602.620 245.730 603.050 246.820 ;
        RECT 631.590 246.790 649.190 246.820 ;
        RECT 645.980 246.090 649.190 246.790 ;
        RECT 679.960 246.690 680.470 247.130 ;
        RECT 749.740 246.900 750.250 247.340 ;
        RECT 756.410 247.110 756.830 247.170 ;
        RECT 749.810 246.880 750.170 246.900 ;
        RECT 680.030 246.670 680.390 246.690 ;
        RECT 756.390 246.530 756.850 247.110 ;
        RECT 756.410 246.470 756.830 246.530 ;
        RECT 676.450 245.840 678.250 246.450 ;
        RECT 679.900 245.840 683.260 245.985 ;
        RECT 601.670 245.100 603.240 245.730 ;
        RECT 676.450 245.615 683.260 245.840 ;
        RECT 685.560 245.625 688.920 245.995 ;
        RECT 690.910 245.645 694.270 246.015 ;
        RECT 676.450 245.475 681.410 245.615 ;
        RECT 687.220 245.485 687.480 245.625 ;
        RECT 676.450 245.370 683.260 245.475 ;
        RECT 685.560 245.430 688.920 245.485 ;
        RECT 689.730 245.430 690.410 245.620 ;
        RECT 692.410 245.505 692.650 245.645 ;
        RECT 697.130 245.635 700.490 246.005 ;
        RECT 702.790 245.645 706.150 246.015 ;
        RECT 708.140 245.665 711.500 246.035 ;
        RECT 714.700 245.735 718.060 246.105 ;
        RECT 720.360 245.745 723.720 246.115 ;
        RECT 725.710 245.765 729.070 246.135 ;
        RECT 731.870 245.765 735.230 246.135 ;
        RECT 737.530 245.775 740.890 246.145 ;
        RECT 742.880 245.795 746.240 246.165 ;
        RECT 749.680 245.825 753.040 246.195 ;
        RECT 755.340 245.835 758.700 246.205 ;
        RECT 760.690 245.855 764.050 246.225 ;
        RECT 690.910 245.470 694.270 245.505 ;
        RECT 698.390 245.495 698.640 245.635 ;
        RECT 704.450 245.505 704.710 245.645 ;
        RECT 697.130 245.470 700.490 245.495 ;
        RECT 690.910 245.430 700.490 245.470 ;
        RECT 685.560 245.390 700.490 245.430 ;
        RECT 702.790 245.450 706.150 245.505 ;
        RECT 706.960 245.450 707.640 245.640 ;
        RECT 709.640 245.525 709.880 245.665 ;
        RECT 715.960 245.595 716.210 245.735 ;
        RECT 722.020 245.605 722.280 245.745 ;
        RECT 708.140 245.500 711.500 245.525 ;
        RECT 714.700 245.500 718.060 245.595 ;
        RECT 708.140 245.490 718.060 245.500 ;
        RECT 720.360 245.550 723.720 245.605 ;
        RECT 724.530 245.550 725.210 245.740 ;
        RECT 727.210 245.625 727.450 245.765 ;
        RECT 733.130 245.625 733.380 245.765 ;
        RECT 739.190 245.635 739.450 245.775 ;
        RECT 725.710 245.550 729.070 245.625 ;
        RECT 720.360 245.490 729.070 245.550 ;
        RECT 708.140 245.480 729.070 245.490 ;
        RECT 731.870 245.520 735.230 245.625 ;
        RECT 737.530 245.580 740.890 245.635 ;
        RECT 741.700 245.580 742.380 245.770 ;
        RECT 744.380 245.655 744.620 245.795 ;
        RECT 750.940 245.685 751.190 245.825 ;
        RECT 757.000 245.695 757.260 245.835 ;
        RECT 742.880 245.600 746.240 245.655 ;
        RECT 749.680 245.600 753.040 245.685 ;
        RECT 742.880 245.580 753.040 245.600 ;
        RECT 755.340 245.640 758.700 245.695 ;
        RECT 759.510 245.640 760.190 245.830 ;
        RECT 762.190 245.715 762.430 245.855 ;
        RECT 760.690 245.640 764.050 245.715 ;
        RECT 755.340 245.580 764.050 245.640 ;
        RECT 737.530 245.520 764.050 245.580 ;
        RECT 731.870 245.485 764.050 245.520 ;
        RECT 731.870 245.480 761.150 245.485 ;
        RECT 708.140 245.465 761.150 245.480 ;
        RECT 708.140 245.455 755.490 245.465 ;
        RECT 708.140 245.450 749.980 245.455 ;
        RECT 702.790 245.425 749.980 245.450 ;
        RECT 702.790 245.405 743.340 245.425 ;
        RECT 702.790 245.395 737.680 245.405 ;
        RECT 702.790 245.390 726.170 245.395 ;
        RECT 685.560 245.375 726.170 245.390 ;
        RECT 685.560 245.370 720.510 245.375 ;
        RECT 676.450 245.365 720.510 245.370 ;
        RECT 676.450 245.320 714.810 245.365 ;
        RECT 676.450 244.390 678.250 245.320 ;
        RECT 679.900 245.295 714.810 245.320 ;
        RECT 717.570 245.300 720.510 245.365 ;
        RECT 723.230 245.360 726.170 245.375 ;
        RECT 679.900 245.275 708.600 245.295 ;
        RECT 679.900 245.255 691.370 245.275 ;
        RECT 679.900 245.245 685.710 245.255 ;
        RECT 682.770 245.180 685.710 245.245 ;
        RECT 688.430 245.240 691.370 245.255 ;
        RECT 693.810 245.265 702.940 245.275 ;
        RECT 689.730 245.080 690.410 245.240 ;
        RECT 693.810 245.160 697.240 245.265 ;
        RECT 700.000 245.200 702.940 245.265 ;
        RECT 705.660 245.260 708.600 245.275 ;
        RECT 706.960 245.100 707.640 245.260 ;
        RECT 711.380 245.190 714.810 245.295 ;
        RECT 724.530 245.200 725.210 245.360 ;
        RECT 728.870 245.270 732.770 245.395 ;
        RECT 734.740 245.330 737.680 245.395 ;
        RECT 740.400 245.390 743.340 245.405 ;
        RECT 746.080 245.390 749.980 245.425 ;
        RECT 752.550 245.390 755.490 245.455 ;
        RECT 758.210 245.450 761.150 245.465 ;
        RECT 741.700 245.230 742.380 245.390 ;
        RECT 759.510 245.290 760.190 245.450 ;
        RECT 192.070 239.190 198.830 243.820 ;
        RECT -97.880 233.315 -97.650 234.530 ;
        RECT -95.300 233.315 -95.070 234.530 ;
        RECT -92.720 233.355 -92.490 234.530 ;
        RECT -90.140 233.375 -89.910 234.530 ;
        RECT -87.560 233.445 -87.330 234.530 ;
        RECT -97.885 232.950 -97.650 233.315 ;
        RECT -95.345 232.950 -95.070 233.315 ;
        RECT -92.745 232.950 -92.490 233.355 ;
        RECT -90.175 232.950 -89.910 233.375 ;
        RECT -87.595 232.950 -87.330 233.445 ;
        RECT -84.980 233.355 -84.750 234.530 ;
        RECT -84.995 232.950 -84.750 233.355 ;
        RECT -82.400 233.445 -82.170 234.530 ;
        RECT -82.400 232.950 -82.165 233.445 ;
        RECT -79.820 233.375 -79.590 234.530 ;
        RECT -77.240 233.375 -77.010 234.530 ;
        RECT -74.660 233.405 -74.430 234.530 ;
        RECT -79.820 232.950 -79.565 233.375 ;
        RECT -77.240 232.950 -76.975 233.375 ;
        RECT -97.885 232.055 -97.655 232.950 ;
        RECT -95.345 232.055 -95.115 232.950 ;
        RECT -92.745 232.055 -92.515 232.950 ;
        RECT -90.175 232.055 -89.945 232.950 ;
        RECT -87.595 232.055 -87.365 232.950 ;
        RECT -84.995 232.055 -84.765 232.950 ;
        RECT -82.395 232.055 -82.165 232.950 ;
        RECT -79.795 232.055 -79.565 232.950 ;
        RECT -77.205 232.055 -76.975 232.950 ;
        RECT -74.705 232.950 -74.430 233.405 ;
        RECT -72.080 233.355 -71.850 234.530 ;
        RECT -72.085 232.950 -71.850 233.355 ;
        RECT -74.705 232.055 -74.475 232.950 ;
        RECT -72.085 232.055 -71.855 232.950 ;
        RECT -97.905 231.755 -71.855 232.055 ;
        RECT -97.885 231.735 -97.655 231.755 ;
        RECT -95.345 231.735 -95.115 231.755 ;
        RECT -83.055 231.080 -82.865 231.755 ;
        RECT -97.390 230.850 -96.850 231.080 ;
        RECT -96.100 230.850 -95.560 231.080 ;
        RECT -94.810 230.850 -94.270 231.080 ;
        RECT -93.520 230.850 -92.980 231.080 ;
        RECT -92.230 230.850 -91.690 231.080 ;
        RECT -90.940 230.850 -90.400 231.080 ;
        RECT -89.650 230.850 -89.110 231.080 ;
        RECT -88.360 230.850 -87.820 231.080 ;
        RECT -87.070 230.850 -86.530 231.080 ;
        RECT -85.780 230.850 -85.240 231.080 ;
        RECT -84.490 230.850 -83.950 231.080 ;
        RECT -83.200 230.850 -82.660 231.080 ;
        RECT -81.910 230.850 -81.370 231.080 ;
        RECT -80.620 230.850 -80.080 231.080 ;
        RECT -79.330 230.850 -78.790 231.080 ;
        RECT -78.040 230.850 -77.500 231.080 ;
        RECT -76.750 230.850 -76.210 231.080 ;
        RECT -75.460 230.850 -74.920 231.080 ;
        RECT -74.170 230.850 -73.630 231.080 ;
        RECT -72.880 230.850 -72.340 231.080 ;
        RECT -91.670 227.820 -78.060 230.500 ;
        RECT 195.450 225.890 197.480 239.190 ;
        RECT 340.940 237.120 344.470 239.060 ;
        RECT 120.120 222.910 127.210 225.350 ;
        RECT -97.190 221.215 -96.960 222.430 ;
        RECT -94.610 221.215 -94.380 222.430 ;
        RECT -92.030 221.255 -91.800 222.430 ;
        RECT -89.450 221.275 -89.220 222.430 ;
        RECT -86.870 221.345 -86.640 222.430 ;
        RECT -97.195 220.850 -96.960 221.215 ;
        RECT -94.655 220.850 -94.380 221.215 ;
        RECT -92.055 220.850 -91.800 221.255 ;
        RECT -89.485 220.850 -89.220 221.275 ;
        RECT -86.905 220.850 -86.640 221.345 ;
        RECT -84.290 221.255 -84.060 222.430 ;
        RECT -84.305 220.850 -84.060 221.255 ;
        RECT -81.710 221.345 -81.480 222.430 ;
        RECT -81.710 220.850 -81.475 221.345 ;
        RECT -79.130 221.275 -78.900 222.430 ;
        RECT -76.550 221.275 -76.320 222.430 ;
        RECT -73.970 221.305 -73.740 222.430 ;
        RECT -79.130 220.850 -78.875 221.275 ;
        RECT -76.550 220.850 -76.285 221.275 ;
        RECT -97.195 219.955 -96.965 220.850 ;
        RECT -94.655 219.955 -94.425 220.850 ;
        RECT -92.055 219.955 -91.825 220.850 ;
        RECT -89.485 219.955 -89.255 220.850 ;
        RECT -86.905 219.955 -86.675 220.850 ;
        RECT -84.305 219.955 -84.075 220.850 ;
        RECT -81.705 219.955 -81.475 220.850 ;
        RECT -79.105 219.955 -78.875 220.850 ;
        RECT -76.515 219.955 -76.285 220.850 ;
        RECT -74.015 220.850 -73.740 221.305 ;
        RECT -71.390 221.255 -71.160 222.430 ;
        RECT 193.570 221.540 213.970 225.890 ;
        RECT -71.395 220.850 -71.160 221.255 ;
        RECT -74.015 219.955 -73.785 220.850 ;
        RECT -71.395 219.955 -71.165 220.850 ;
        RECT -97.215 219.655 -71.165 219.955 ;
        RECT -97.195 219.635 -96.965 219.655 ;
        RECT -94.655 219.635 -94.425 219.655 ;
        RECT -82.365 218.980 -82.175 219.655 ;
        RECT -96.700 218.750 -96.160 218.980 ;
        RECT -95.410 218.750 -94.870 218.980 ;
        RECT -94.120 218.750 -93.580 218.980 ;
        RECT -92.830 218.750 -92.290 218.980 ;
        RECT -91.540 218.750 -91.000 218.980 ;
        RECT -90.250 218.750 -89.710 218.980 ;
        RECT -88.960 218.750 -88.420 218.980 ;
        RECT -87.670 218.750 -87.130 218.980 ;
        RECT -86.380 218.750 -85.840 218.980 ;
        RECT -85.090 218.750 -84.550 218.980 ;
        RECT -83.800 218.750 -83.260 218.980 ;
        RECT -82.510 218.750 -81.970 218.980 ;
        RECT -81.220 218.750 -80.680 218.980 ;
        RECT -79.930 218.750 -79.390 218.980 ;
        RECT -78.640 218.750 -78.100 218.980 ;
        RECT -77.350 218.750 -76.810 218.980 ;
        RECT -76.060 218.750 -75.520 218.980 ;
        RECT -74.770 218.750 -74.230 218.980 ;
        RECT -73.480 218.750 -72.940 218.980 ;
        RECT -72.190 218.750 -71.650 218.980 ;
        RECT -91.040 215.700 -77.430 218.380 ;
        RECT 55.080 217.830 56.450 218.870 ;
        RECT 247.270 218.070 250.350 220.020 ;
        RECT 342.040 219.920 343.050 237.120 ;
        RECT 341.380 218.910 345.300 219.920 ;
        RECT 318.960 217.220 321.190 218.260 ;
        RECT 357.850 217.130 359.390 218.190 ;
        RECT 9.760 213.740 9.990 215.320 ;
        RECT 15.050 213.740 15.280 215.320 ;
        RECT 20.340 213.740 20.570 215.320 ;
        RECT 25.630 213.740 25.860 215.320 ;
        RECT 30.920 213.740 31.150 215.320 ;
        RECT 36.210 213.740 36.440 215.320 ;
        RECT 42.330 213.780 42.560 215.360 ;
        RECT 47.620 213.780 47.850 215.360 ;
        RECT 52.910 213.780 53.140 215.360 ;
        RECT 58.200 213.780 58.430 215.360 ;
        RECT 63.490 213.780 63.720 215.360 ;
        RECT 68.780 213.780 69.010 215.360 ;
        RECT 74.860 213.820 75.090 215.400 ;
        RECT 80.150 213.820 80.380 215.400 ;
        RECT 85.440 213.820 85.670 215.400 ;
        RECT 90.730 213.820 90.960 215.400 ;
        RECT 96.020 213.820 96.250 215.400 ;
        RECT 101.310 213.820 101.540 215.400 ;
        RECT 9.760 208.270 9.990 209.850 ;
        RECT 15.050 208.270 15.280 209.850 ;
        RECT 20.340 208.270 20.570 209.850 ;
        RECT 25.630 208.270 25.860 209.850 ;
        RECT 30.920 208.270 31.150 209.850 ;
        RECT 36.210 208.270 36.440 209.850 ;
        RECT 6.520 207.080 7.270 208.220 ;
        RECT -97.590 133.465 -97.360 134.680 ;
        RECT -95.010 133.465 -94.780 134.680 ;
        RECT -92.430 133.505 -92.200 134.680 ;
        RECT -89.850 133.525 -89.620 134.680 ;
        RECT -87.270 133.595 -87.040 134.680 ;
        RECT -97.595 133.100 -97.360 133.465 ;
        RECT -95.055 133.100 -94.780 133.465 ;
        RECT -92.455 133.100 -92.200 133.505 ;
        RECT -89.885 133.100 -89.620 133.525 ;
        RECT -87.305 133.100 -87.040 133.595 ;
        RECT -84.690 133.505 -84.460 134.680 ;
        RECT -84.705 133.100 -84.460 133.505 ;
        RECT -82.110 133.595 -81.880 134.680 ;
        RECT -82.110 133.100 -81.875 133.595 ;
        RECT -79.530 133.525 -79.300 134.680 ;
        RECT -76.950 133.525 -76.720 134.680 ;
        RECT -74.370 133.555 -74.140 134.680 ;
        RECT -79.530 133.100 -79.275 133.525 ;
        RECT -76.950 133.100 -76.685 133.525 ;
        RECT -97.595 132.205 -97.365 133.100 ;
        RECT -95.055 132.205 -94.825 133.100 ;
        RECT -92.455 132.205 -92.225 133.100 ;
        RECT -89.885 132.205 -89.655 133.100 ;
        RECT -87.305 132.205 -87.075 133.100 ;
        RECT -84.705 132.205 -84.475 133.100 ;
        RECT -82.105 132.205 -81.875 133.100 ;
        RECT -79.505 132.205 -79.275 133.100 ;
        RECT -76.915 132.205 -76.685 133.100 ;
        RECT -74.415 133.100 -74.140 133.555 ;
        RECT -71.790 133.505 -71.560 134.680 ;
        RECT -71.795 133.100 -71.560 133.505 ;
        RECT -74.415 132.205 -74.185 133.100 ;
        RECT -71.795 132.205 -71.565 133.100 ;
        RECT -97.615 131.905 -71.565 132.205 ;
        RECT -97.595 131.885 -97.365 131.905 ;
        RECT -95.055 131.885 -94.825 131.905 ;
        RECT -82.765 131.230 -82.575 131.905 ;
        RECT -97.100 131.000 -96.560 131.230 ;
        RECT -95.810 131.000 -95.270 131.230 ;
        RECT -94.520 131.000 -93.980 131.230 ;
        RECT -93.230 131.000 -92.690 131.230 ;
        RECT -91.940 131.000 -91.400 131.230 ;
        RECT -90.650 131.000 -90.110 131.230 ;
        RECT -89.360 131.000 -88.820 131.230 ;
        RECT -88.070 131.000 -87.530 131.230 ;
        RECT -86.780 131.000 -86.240 131.230 ;
        RECT -85.490 131.000 -84.950 131.230 ;
        RECT -84.200 131.000 -83.660 131.230 ;
        RECT -82.910 131.000 -82.370 131.230 ;
        RECT -81.620 131.000 -81.080 131.230 ;
        RECT -80.330 131.000 -79.790 131.230 ;
        RECT -79.040 131.000 -78.500 131.230 ;
        RECT -77.750 131.000 -77.210 131.230 ;
        RECT -76.460 131.000 -75.920 131.230 ;
        RECT -75.170 131.000 -74.630 131.230 ;
        RECT -73.880 131.000 -73.340 131.230 ;
        RECT -72.590 131.000 -72.050 131.230 ;
        RECT -91.500 127.860 -77.890 130.540 ;
        RECT -97.160 14.135 -96.930 15.350 ;
        RECT -94.580 14.135 -94.350 15.350 ;
        RECT -92.000 14.175 -91.770 15.350 ;
        RECT -89.420 14.195 -89.190 15.350 ;
        RECT -86.840 14.265 -86.610 15.350 ;
        RECT -97.165 13.770 -96.930 14.135 ;
        RECT -94.625 13.770 -94.350 14.135 ;
        RECT -92.025 13.770 -91.770 14.175 ;
        RECT -89.455 13.770 -89.190 14.195 ;
        RECT -86.875 13.770 -86.610 14.265 ;
        RECT -84.260 14.175 -84.030 15.350 ;
        RECT -84.275 13.770 -84.030 14.175 ;
        RECT -81.680 14.265 -81.450 15.350 ;
        RECT -81.680 13.770 -81.445 14.265 ;
        RECT -79.100 14.195 -78.870 15.350 ;
        RECT -76.520 14.195 -76.290 15.350 ;
        RECT -73.940 14.225 -73.710 15.350 ;
        RECT -79.100 13.770 -78.845 14.195 ;
        RECT -76.520 13.770 -76.255 14.195 ;
        RECT -97.165 12.875 -96.935 13.770 ;
        RECT -94.625 12.875 -94.395 13.770 ;
        RECT -92.025 12.875 -91.795 13.770 ;
        RECT -89.455 12.875 -89.225 13.770 ;
        RECT -86.875 12.875 -86.645 13.770 ;
        RECT -84.275 12.875 -84.045 13.770 ;
        RECT -81.675 12.875 -81.445 13.770 ;
        RECT -79.075 12.875 -78.845 13.770 ;
        RECT -76.485 12.875 -76.255 13.770 ;
        RECT -73.985 13.770 -73.710 14.225 ;
        RECT -71.360 14.175 -71.130 15.350 ;
        RECT -71.365 13.770 -71.130 14.175 ;
        RECT -73.985 12.875 -73.755 13.770 ;
        RECT -71.365 12.875 -71.135 13.770 ;
        RECT -97.185 12.575 -71.135 12.875 ;
        RECT -97.165 12.555 -96.935 12.575 ;
        RECT -94.625 12.555 -94.395 12.575 ;
        RECT -82.335 11.900 -82.145 12.575 ;
        RECT -96.670 11.670 -96.130 11.900 ;
        RECT -95.380 11.670 -94.840 11.900 ;
        RECT -94.090 11.670 -93.550 11.900 ;
        RECT -92.800 11.670 -92.260 11.900 ;
        RECT -91.510 11.670 -90.970 11.900 ;
        RECT -90.220 11.670 -89.680 11.900 ;
        RECT -88.930 11.670 -88.390 11.900 ;
        RECT -87.640 11.670 -87.100 11.900 ;
        RECT -86.350 11.670 -85.810 11.900 ;
        RECT -85.060 11.670 -84.520 11.900 ;
        RECT -83.770 11.670 -83.230 11.900 ;
        RECT -82.480 11.670 -81.940 11.900 ;
        RECT -81.190 11.670 -80.650 11.900 ;
        RECT -79.900 11.670 -79.360 11.900 ;
        RECT -78.610 11.670 -78.070 11.900 ;
        RECT -77.320 11.670 -76.780 11.900 ;
        RECT -76.030 11.670 -75.490 11.900 ;
        RECT -74.740 11.670 -74.200 11.900 ;
        RECT -73.450 11.670 -72.910 11.900 ;
        RECT -72.160 11.670 -71.620 11.900 ;
        RECT -90.760 8.650 -77.150 11.330 ;
        RECT 6.320 -12.700 7.800 207.080 ;
        RECT 9.760 202.800 9.990 204.380 ;
        RECT 15.050 202.800 15.280 204.380 ;
        RECT 20.340 202.800 20.570 204.380 ;
        RECT 25.630 202.800 25.860 204.380 ;
        RECT 30.920 202.800 31.150 204.380 ;
        RECT 36.210 202.800 36.440 204.380 ;
        RECT 37.980 204.190 41.260 210.950 ;
        RECT 42.330 208.310 42.560 209.890 ;
        RECT 47.620 208.310 47.850 209.890 ;
        RECT 52.910 208.310 53.140 209.890 ;
        RECT 58.200 208.310 58.430 209.890 ;
        RECT 63.490 208.310 63.720 209.890 ;
        RECT 68.780 208.310 69.010 209.890 ;
        RECT 42.330 204.190 42.560 204.420 ;
        RECT 37.980 202.840 42.560 204.190 ;
        RECT 47.620 202.840 47.850 204.420 ;
        RECT 52.910 202.840 53.140 204.420 ;
        RECT 58.200 202.840 58.430 204.420 ;
        RECT 63.490 202.840 63.720 204.420 ;
        RECT 68.780 204.380 69.010 204.420 ;
        RECT 70.230 204.380 73.430 208.450 ;
        RECT 74.860 208.350 75.090 209.930 ;
        RECT 80.150 208.350 80.380 209.930 ;
        RECT 85.440 208.350 85.670 209.930 ;
        RECT 90.730 208.350 90.960 209.930 ;
        RECT 96.020 208.350 96.250 209.930 ;
        RECT 101.310 208.350 101.540 209.930 ;
        RECT 68.780 202.870 73.430 204.380 ;
        RECT 74.860 202.880 75.090 204.460 ;
        RECT 80.150 202.880 80.380 204.460 ;
        RECT 85.440 202.880 85.670 204.460 ;
        RECT 90.730 202.880 90.960 204.460 ;
        RECT 96.020 202.880 96.250 204.460 ;
        RECT 101.310 202.880 101.540 204.460 ;
        RECT 102.800 204.200 106.000 209.470 ;
        RECT 68.780 202.840 69.010 202.870 ;
        RECT 37.980 202.680 42.480 202.840 ;
        RECT 9.760 197.330 9.990 198.910 ;
        RECT 15.050 197.330 15.280 198.910 ;
        RECT 20.340 197.330 20.570 198.910 ;
        RECT 25.630 197.330 25.860 198.910 ;
        RECT 30.920 197.330 31.150 198.910 ;
        RECT 36.210 197.330 36.440 198.910 ;
        RECT 9.760 191.860 9.990 193.440 ;
        RECT 15.050 191.860 15.280 193.440 ;
        RECT 20.340 191.860 20.570 193.440 ;
        RECT 25.630 191.860 25.860 193.440 ;
        RECT 30.920 191.860 31.150 193.440 ;
        RECT 36.210 191.860 36.440 193.440 ;
        RECT 9.760 184.660 9.990 186.240 ;
        RECT 15.050 184.660 15.280 186.240 ;
        RECT 20.340 184.660 20.570 186.240 ;
        RECT 25.630 184.660 25.860 186.240 ;
        RECT 30.920 184.660 31.150 186.240 ;
        RECT 36.210 184.660 36.440 186.240 ;
        RECT 9.760 179.190 9.990 180.770 ;
        RECT 15.050 179.190 15.280 180.770 ;
        RECT 20.340 179.190 20.570 180.770 ;
        RECT 25.630 179.190 25.860 180.770 ;
        RECT 30.920 179.190 31.150 180.770 ;
        RECT 36.210 179.190 36.440 180.770 ;
        RECT 9.760 173.720 9.990 175.300 ;
        RECT 15.050 173.720 15.280 175.300 ;
        RECT 20.340 173.720 20.570 175.300 ;
        RECT 25.630 173.720 25.860 175.300 ;
        RECT 30.920 173.720 31.150 175.300 ;
        RECT 36.210 173.720 36.440 175.300 ;
        RECT 9.760 168.250 9.990 169.830 ;
        RECT 15.050 168.250 15.280 169.830 ;
        RECT 20.340 168.250 20.570 169.830 ;
        RECT 25.630 168.250 25.860 169.830 ;
        RECT 30.920 168.250 31.150 169.830 ;
        RECT 36.210 168.250 36.440 169.830 ;
        RECT 9.760 162.780 9.990 164.360 ;
        RECT 15.050 162.780 15.280 164.360 ;
        RECT 20.340 162.780 20.570 164.360 ;
        RECT 25.630 162.780 25.860 164.360 ;
        RECT 30.920 162.780 31.150 164.360 ;
        RECT 36.210 162.780 36.440 164.360 ;
        RECT 9.760 155.490 9.990 157.070 ;
        RECT 15.050 155.490 15.280 157.070 ;
        RECT 20.340 155.490 20.570 157.070 ;
        RECT 25.630 155.490 25.860 157.070 ;
        RECT 30.920 155.490 31.150 157.070 ;
        RECT 36.210 155.490 36.440 157.070 ;
        RECT 9.760 150.020 9.990 151.600 ;
        RECT 15.050 150.020 15.280 151.600 ;
        RECT 20.340 150.020 20.570 151.600 ;
        RECT 25.630 150.020 25.860 151.600 ;
        RECT 30.920 150.020 31.150 151.600 ;
        RECT 36.210 150.020 36.440 151.600 ;
        RECT 9.760 144.550 9.990 146.130 ;
        RECT 15.050 144.550 15.280 146.130 ;
        RECT 20.340 144.550 20.570 146.130 ;
        RECT 25.630 144.550 25.860 146.130 ;
        RECT 30.920 144.550 31.150 146.130 ;
        RECT 36.210 144.550 36.440 146.130 ;
        RECT 9.760 139.080 9.990 140.660 ;
        RECT 15.050 139.080 15.280 140.660 ;
        RECT 20.340 139.080 20.570 140.660 ;
        RECT 25.630 139.080 25.860 140.660 ;
        RECT 30.920 139.080 31.150 140.660 ;
        RECT 36.210 139.080 36.440 140.660 ;
        RECT 9.760 133.610 9.990 135.190 ;
        RECT 15.050 133.610 15.280 135.190 ;
        RECT 20.340 133.610 20.570 135.190 ;
        RECT 25.630 133.610 25.860 135.190 ;
        RECT 30.920 133.610 31.150 135.190 ;
        RECT 36.210 133.610 36.440 135.190 ;
        RECT 9.760 126.310 9.990 127.890 ;
        RECT 15.050 126.310 15.280 127.890 ;
        RECT 20.340 126.310 20.570 127.890 ;
        RECT 25.630 126.310 25.860 127.890 ;
        RECT 30.920 126.310 31.150 127.890 ;
        RECT 36.210 126.310 36.440 127.890 ;
        RECT 9.760 120.840 9.990 122.420 ;
        RECT 15.050 120.840 15.280 122.420 ;
        RECT 20.340 120.840 20.570 122.420 ;
        RECT 25.630 120.840 25.860 122.420 ;
        RECT 30.920 120.840 31.150 122.420 ;
        RECT 36.210 120.840 36.440 122.420 ;
        RECT 9.760 115.370 9.990 116.950 ;
        RECT 15.050 115.370 15.280 116.950 ;
        RECT 20.340 115.370 20.570 116.950 ;
        RECT 25.630 115.370 25.860 116.950 ;
        RECT 30.920 115.370 31.150 116.950 ;
        RECT 36.210 115.370 36.440 116.950 ;
        RECT 9.760 109.900 9.990 111.480 ;
        RECT 15.050 109.900 15.280 111.480 ;
        RECT 20.340 109.900 20.570 111.480 ;
        RECT 25.630 109.900 25.860 111.480 ;
        RECT 30.920 109.900 31.150 111.480 ;
        RECT 36.210 109.900 36.440 111.480 ;
        RECT 9.760 104.430 9.990 106.010 ;
        RECT 15.050 104.430 15.280 106.010 ;
        RECT 20.340 104.430 20.570 106.010 ;
        RECT 25.630 104.430 25.860 106.010 ;
        RECT 30.920 104.430 31.150 106.010 ;
        RECT 36.210 104.430 36.440 106.010 ;
        RECT 9.760 96.990 9.990 98.570 ;
        RECT 15.050 96.990 15.280 98.570 ;
        RECT 20.340 96.990 20.570 98.570 ;
        RECT 25.630 96.990 25.860 98.570 ;
        RECT 30.920 96.990 31.150 98.570 ;
        RECT 36.210 96.990 36.440 98.570 ;
        RECT 9.760 91.520 9.990 93.100 ;
        RECT 15.050 91.520 15.280 93.100 ;
        RECT 20.340 91.520 20.570 93.100 ;
        RECT 25.630 91.520 25.860 93.100 ;
        RECT 30.920 91.520 31.150 93.100 ;
        RECT 36.210 91.520 36.440 93.100 ;
        RECT 9.760 86.050 9.990 87.630 ;
        RECT 15.050 86.050 15.280 87.630 ;
        RECT 20.340 86.050 20.570 87.630 ;
        RECT 25.630 86.050 25.860 87.630 ;
        RECT 30.920 86.050 31.150 87.630 ;
        RECT 36.210 86.050 36.440 87.630 ;
        RECT 9.760 80.580 9.990 82.160 ;
        RECT 15.050 80.580 15.280 82.160 ;
        RECT 20.340 80.580 20.570 82.160 ;
        RECT 25.630 80.580 25.860 82.160 ;
        RECT 30.920 80.580 31.150 82.160 ;
        RECT 36.210 80.580 36.440 82.160 ;
        RECT 9.760 75.110 9.990 76.690 ;
        RECT 15.050 75.110 15.280 76.690 ;
        RECT 20.340 75.110 20.570 76.690 ;
        RECT 25.630 75.110 25.860 76.690 ;
        RECT 30.920 75.110 31.150 76.690 ;
        RECT 36.210 75.110 36.440 76.690 ;
        RECT 9.810 67.710 10.040 69.290 ;
        RECT 15.100 67.710 15.330 69.290 ;
        RECT 20.390 67.710 20.620 69.290 ;
        RECT 25.680 67.710 25.910 69.290 ;
        RECT 30.970 67.710 31.200 69.290 ;
        RECT 36.260 67.710 36.490 69.290 ;
        RECT 9.810 62.240 10.040 63.820 ;
        RECT 15.100 62.240 15.330 63.820 ;
        RECT 20.390 62.240 20.620 63.820 ;
        RECT 25.680 62.240 25.910 63.820 ;
        RECT 30.970 62.240 31.200 63.820 ;
        RECT 36.260 62.240 36.490 63.820 ;
        RECT 9.810 56.770 10.040 58.350 ;
        RECT 15.100 56.770 15.330 58.350 ;
        RECT 20.390 56.770 20.620 58.350 ;
        RECT 25.680 56.770 25.910 58.350 ;
        RECT 30.970 56.770 31.200 58.350 ;
        RECT 36.260 56.770 36.490 58.350 ;
        RECT 9.810 51.300 10.040 52.880 ;
        RECT 15.100 51.300 15.330 52.880 ;
        RECT 20.390 51.300 20.620 52.880 ;
        RECT 25.680 51.300 25.910 52.880 ;
        RECT 30.970 51.300 31.200 52.880 ;
        RECT 36.260 51.300 36.490 52.880 ;
        RECT 9.810 45.830 10.040 47.410 ;
        RECT 15.100 45.830 15.330 47.410 ;
        RECT 20.390 45.830 20.620 47.410 ;
        RECT 25.680 45.830 25.910 47.410 ;
        RECT 30.970 45.830 31.200 47.410 ;
        RECT 36.260 45.830 36.490 47.410 ;
        RECT 9.900 38.170 10.130 39.750 ;
        RECT 15.190 38.170 15.420 39.750 ;
        RECT 20.480 38.170 20.710 39.750 ;
        RECT 25.770 38.170 26.000 39.750 ;
        RECT 31.060 38.170 31.290 39.750 ;
        RECT 36.350 38.170 36.580 39.750 ;
        RECT 9.900 32.700 10.130 34.280 ;
        RECT 15.190 32.700 15.420 34.280 ;
        RECT 20.480 32.700 20.710 34.280 ;
        RECT 25.770 32.700 26.000 34.280 ;
        RECT 31.060 32.700 31.290 34.280 ;
        RECT 36.350 32.700 36.580 34.280 ;
        RECT 9.900 27.230 10.130 28.810 ;
        RECT 15.190 27.230 15.420 28.810 ;
        RECT 20.480 27.230 20.710 28.810 ;
        RECT 25.770 27.230 26.000 28.810 ;
        RECT 31.060 27.230 31.290 28.810 ;
        RECT 36.350 27.230 36.580 28.810 ;
        RECT 37.980 24.860 41.260 202.680 ;
        RECT 42.330 197.370 42.560 198.950 ;
        RECT 47.620 197.370 47.850 198.950 ;
        RECT 52.910 197.370 53.140 198.950 ;
        RECT 58.200 197.370 58.430 198.950 ;
        RECT 63.490 197.370 63.720 198.950 ;
        RECT 68.780 197.370 69.010 198.950 ;
        RECT 42.330 191.900 42.560 193.480 ;
        RECT 47.620 191.900 47.850 193.480 ;
        RECT 52.910 191.900 53.140 193.480 ;
        RECT 58.200 191.900 58.430 193.480 ;
        RECT 63.490 191.900 63.720 193.480 ;
        RECT 68.780 191.900 69.010 193.480 ;
        RECT 42.330 184.700 42.560 186.280 ;
        RECT 47.620 184.700 47.850 186.280 ;
        RECT 52.910 184.700 53.140 186.280 ;
        RECT 58.200 184.700 58.430 186.280 ;
        RECT 63.490 184.700 63.720 186.280 ;
        RECT 68.780 184.700 69.010 186.280 ;
        RECT 42.330 179.230 42.560 180.810 ;
        RECT 47.620 179.230 47.850 180.810 ;
        RECT 52.910 179.230 53.140 180.810 ;
        RECT 58.200 179.230 58.430 180.810 ;
        RECT 63.490 179.230 63.720 180.810 ;
        RECT 68.780 179.230 69.010 180.810 ;
        RECT 42.330 173.760 42.560 175.340 ;
        RECT 47.620 173.760 47.850 175.340 ;
        RECT 52.910 173.760 53.140 175.340 ;
        RECT 58.200 173.760 58.430 175.340 ;
        RECT 63.490 173.760 63.720 175.340 ;
        RECT 68.780 173.760 69.010 175.340 ;
        RECT 42.330 168.290 42.560 169.870 ;
        RECT 47.620 168.290 47.850 169.870 ;
        RECT 52.910 168.290 53.140 169.870 ;
        RECT 58.200 168.290 58.430 169.870 ;
        RECT 63.490 168.290 63.720 169.870 ;
        RECT 68.780 168.290 69.010 169.870 ;
        RECT 42.330 162.820 42.560 164.400 ;
        RECT 47.620 162.820 47.850 164.400 ;
        RECT 52.910 162.820 53.140 164.400 ;
        RECT 58.200 162.820 58.430 164.400 ;
        RECT 63.490 162.820 63.720 164.400 ;
        RECT 68.780 162.820 69.010 164.400 ;
        RECT 42.330 155.530 42.560 157.110 ;
        RECT 47.620 155.530 47.850 157.110 ;
        RECT 52.910 155.530 53.140 157.110 ;
        RECT 58.200 155.530 58.430 157.110 ;
        RECT 63.490 155.530 63.720 157.110 ;
        RECT 68.780 155.530 69.010 157.110 ;
        RECT 42.330 150.060 42.560 151.640 ;
        RECT 47.620 150.060 47.850 151.640 ;
        RECT 52.910 150.060 53.140 151.640 ;
        RECT 58.200 150.060 58.430 151.640 ;
        RECT 63.490 150.060 63.720 151.640 ;
        RECT 68.780 150.060 69.010 151.640 ;
        RECT 42.330 144.590 42.560 146.170 ;
        RECT 47.620 144.590 47.850 146.170 ;
        RECT 52.910 144.590 53.140 146.170 ;
        RECT 58.200 144.590 58.430 146.170 ;
        RECT 63.490 144.590 63.720 146.170 ;
        RECT 68.780 144.590 69.010 146.170 ;
        RECT 42.330 139.120 42.560 140.700 ;
        RECT 47.620 139.120 47.850 140.700 ;
        RECT 52.910 139.120 53.140 140.700 ;
        RECT 58.200 139.120 58.430 140.700 ;
        RECT 63.490 139.120 63.720 140.700 ;
        RECT 68.780 139.120 69.010 140.700 ;
        RECT 42.330 133.650 42.560 135.230 ;
        RECT 47.620 133.650 47.850 135.230 ;
        RECT 52.910 133.650 53.140 135.230 ;
        RECT 58.200 133.650 58.430 135.230 ;
        RECT 63.490 133.650 63.720 135.230 ;
        RECT 68.780 133.650 69.010 135.230 ;
        RECT 42.330 126.350 42.560 127.930 ;
        RECT 47.620 126.350 47.850 127.930 ;
        RECT 52.910 126.350 53.140 127.930 ;
        RECT 58.200 126.350 58.430 127.930 ;
        RECT 63.490 126.350 63.720 127.930 ;
        RECT 68.780 126.350 69.010 127.930 ;
        RECT 42.330 120.880 42.560 122.460 ;
        RECT 47.620 120.880 47.850 122.460 ;
        RECT 52.910 120.880 53.140 122.460 ;
        RECT 58.200 120.880 58.430 122.460 ;
        RECT 63.490 120.880 63.720 122.460 ;
        RECT 68.780 120.880 69.010 122.460 ;
        RECT 42.330 115.410 42.560 116.990 ;
        RECT 47.620 115.410 47.850 116.990 ;
        RECT 52.910 115.410 53.140 116.990 ;
        RECT 58.200 115.410 58.430 116.990 ;
        RECT 63.490 115.410 63.720 116.990 ;
        RECT 68.780 115.410 69.010 116.990 ;
        RECT 42.330 109.940 42.560 111.520 ;
        RECT 47.620 109.940 47.850 111.520 ;
        RECT 52.910 109.940 53.140 111.520 ;
        RECT 58.200 109.940 58.430 111.520 ;
        RECT 63.490 109.940 63.720 111.520 ;
        RECT 68.780 109.940 69.010 111.520 ;
        RECT 42.330 104.470 42.560 106.050 ;
        RECT 47.620 104.470 47.850 106.050 ;
        RECT 52.910 104.470 53.140 106.050 ;
        RECT 58.200 104.470 58.430 106.050 ;
        RECT 63.490 104.470 63.720 106.050 ;
        RECT 68.780 104.470 69.010 106.050 ;
        RECT 42.330 97.030 42.560 98.610 ;
        RECT 47.620 97.030 47.850 98.610 ;
        RECT 52.910 97.030 53.140 98.610 ;
        RECT 58.200 97.030 58.430 98.610 ;
        RECT 63.490 97.030 63.720 98.610 ;
        RECT 68.780 97.030 69.010 98.610 ;
        RECT 42.330 91.560 42.560 93.140 ;
        RECT 47.620 91.560 47.850 93.140 ;
        RECT 52.910 91.560 53.140 93.140 ;
        RECT 58.200 91.560 58.430 93.140 ;
        RECT 63.490 91.560 63.720 93.140 ;
        RECT 68.780 91.560 69.010 93.140 ;
        RECT 42.330 86.090 42.560 87.670 ;
        RECT 47.620 86.090 47.850 87.670 ;
        RECT 52.910 86.090 53.140 87.670 ;
        RECT 58.200 86.090 58.430 87.670 ;
        RECT 63.490 86.090 63.720 87.670 ;
        RECT 68.780 86.090 69.010 87.670 ;
        RECT 42.330 80.620 42.560 82.200 ;
        RECT 47.620 80.620 47.850 82.200 ;
        RECT 52.910 80.620 53.140 82.200 ;
        RECT 58.200 80.620 58.430 82.200 ;
        RECT 63.490 80.620 63.720 82.200 ;
        RECT 68.780 80.620 69.010 82.200 ;
        RECT 42.330 75.150 42.560 76.730 ;
        RECT 47.620 75.150 47.850 76.730 ;
        RECT 52.910 75.150 53.140 76.730 ;
        RECT 58.200 75.150 58.430 76.730 ;
        RECT 63.490 75.150 63.720 76.730 ;
        RECT 68.780 75.150 69.010 76.730 ;
        RECT 42.380 67.750 42.610 69.330 ;
        RECT 47.670 67.750 47.900 69.330 ;
        RECT 52.960 67.750 53.190 69.330 ;
        RECT 58.250 67.750 58.480 69.330 ;
        RECT 63.540 67.750 63.770 69.330 ;
        RECT 68.830 67.750 69.060 69.330 ;
        RECT 42.380 62.280 42.610 63.860 ;
        RECT 47.670 62.280 47.900 63.860 ;
        RECT 52.960 62.280 53.190 63.860 ;
        RECT 58.250 62.280 58.480 63.860 ;
        RECT 63.540 62.280 63.770 63.860 ;
        RECT 68.830 62.280 69.060 63.860 ;
        RECT 42.380 56.810 42.610 58.390 ;
        RECT 47.670 56.810 47.900 58.390 ;
        RECT 52.960 56.810 53.190 58.390 ;
        RECT 58.250 56.810 58.480 58.390 ;
        RECT 63.540 56.810 63.770 58.390 ;
        RECT 68.830 56.810 69.060 58.390 ;
        RECT 42.380 51.340 42.610 52.920 ;
        RECT 47.670 51.340 47.900 52.920 ;
        RECT 52.960 51.340 53.190 52.920 ;
        RECT 58.250 51.340 58.480 52.920 ;
        RECT 63.540 51.340 63.770 52.920 ;
        RECT 68.830 51.340 69.060 52.920 ;
        RECT 42.380 45.870 42.610 47.450 ;
        RECT 47.670 45.870 47.900 47.450 ;
        RECT 52.960 45.870 53.190 47.450 ;
        RECT 58.250 45.870 58.480 47.450 ;
        RECT 63.540 45.870 63.770 47.450 ;
        RECT 68.830 45.870 69.060 47.450 ;
        RECT 42.470 38.210 42.700 39.790 ;
        RECT 47.760 38.210 47.990 39.790 ;
        RECT 53.050 38.210 53.280 39.790 ;
        RECT 58.340 38.210 58.570 39.790 ;
        RECT 63.630 38.210 63.860 39.790 ;
        RECT 68.920 38.210 69.150 39.790 ;
        RECT 42.470 32.740 42.700 34.320 ;
        RECT 47.760 32.740 47.990 34.320 ;
        RECT 53.050 32.740 53.280 34.320 ;
        RECT 58.340 32.740 58.570 34.320 ;
        RECT 63.630 32.740 63.860 34.320 ;
        RECT 68.920 32.740 69.150 34.320 ;
        RECT 42.470 27.270 42.700 28.850 ;
        RECT 47.760 27.270 47.990 28.850 ;
        RECT 53.050 27.270 53.280 28.850 ;
        RECT 58.340 27.270 58.570 28.850 ;
        RECT 63.630 27.270 63.860 28.850 ;
        RECT 68.920 27.270 69.150 28.850 ;
        RECT 9.900 21.760 10.130 23.340 ;
        RECT 15.190 21.760 15.420 23.340 ;
        RECT 20.480 21.760 20.710 23.340 ;
        RECT 25.770 21.760 26.000 23.340 ;
        RECT 31.060 21.760 31.290 23.340 ;
        RECT 36.350 21.760 36.580 23.340 ;
        RECT 9.900 16.290 10.130 17.870 ;
        RECT 15.190 16.290 15.420 17.870 ;
        RECT 20.480 16.290 20.710 17.870 ;
        RECT 25.770 16.290 26.000 17.870 ;
        RECT 31.060 16.290 31.290 17.870 ;
        RECT 36.350 16.290 36.580 17.870 ;
        RECT 5.960 -14.640 7.800 -12.700 ;
        RECT -106.270 -15.670 -64.700 -15.510 ;
        RECT 5.960 -15.670 7.740 -14.640 ;
        RECT 38.610 -15.670 40.090 24.860 ;
        RECT 42.470 21.800 42.700 23.380 ;
        RECT 47.760 21.800 47.990 23.380 ;
        RECT 53.050 21.800 53.280 23.380 ;
        RECT 58.340 21.800 58.570 23.380 ;
        RECT 63.630 21.800 63.860 23.380 ;
        RECT 68.920 21.800 69.150 23.380 ;
        RECT 42.470 16.330 42.700 17.910 ;
        RECT 47.760 16.330 47.990 17.910 ;
        RECT 53.050 16.330 53.280 17.910 ;
        RECT 58.340 16.330 58.570 17.910 ;
        RECT 63.630 16.330 63.860 17.910 ;
        RECT 68.920 16.330 69.150 17.910 ;
        RECT 70.230 16.890 73.430 202.870 ;
        RECT 101.690 202.690 106.000 204.200 ;
        RECT 74.860 197.410 75.090 198.990 ;
        RECT 80.150 197.410 80.380 198.990 ;
        RECT 85.440 197.410 85.670 198.990 ;
        RECT 90.730 197.410 90.960 198.990 ;
        RECT 96.020 197.410 96.250 198.990 ;
        RECT 101.310 197.410 101.540 198.990 ;
        RECT 74.860 191.940 75.090 193.520 ;
        RECT 80.150 191.940 80.380 193.520 ;
        RECT 85.440 191.940 85.670 193.520 ;
        RECT 90.730 191.940 90.960 193.520 ;
        RECT 96.020 191.940 96.250 193.520 ;
        RECT 101.310 191.940 101.540 193.520 ;
        RECT 74.860 184.740 75.090 186.320 ;
        RECT 80.150 184.740 80.380 186.320 ;
        RECT 85.440 184.740 85.670 186.320 ;
        RECT 90.730 184.740 90.960 186.320 ;
        RECT 96.020 184.740 96.250 186.320 ;
        RECT 101.310 184.740 101.540 186.320 ;
        RECT 74.860 179.270 75.090 180.850 ;
        RECT 80.150 179.270 80.380 180.850 ;
        RECT 85.440 179.270 85.670 180.850 ;
        RECT 90.730 179.270 90.960 180.850 ;
        RECT 96.020 179.270 96.250 180.850 ;
        RECT 101.310 179.270 101.540 180.850 ;
        RECT 74.860 173.800 75.090 175.380 ;
        RECT 80.150 173.800 80.380 175.380 ;
        RECT 85.440 173.800 85.670 175.380 ;
        RECT 90.730 173.800 90.960 175.380 ;
        RECT 96.020 173.800 96.250 175.380 ;
        RECT 101.310 173.800 101.540 175.380 ;
        RECT 74.860 168.330 75.090 169.910 ;
        RECT 80.150 168.330 80.380 169.910 ;
        RECT 85.440 168.330 85.670 169.910 ;
        RECT 90.730 168.330 90.960 169.910 ;
        RECT 96.020 168.330 96.250 169.910 ;
        RECT 101.310 168.330 101.540 169.910 ;
        RECT 74.860 162.860 75.090 164.440 ;
        RECT 80.150 162.860 80.380 164.440 ;
        RECT 85.440 162.860 85.670 164.440 ;
        RECT 90.730 162.860 90.960 164.440 ;
        RECT 96.020 162.860 96.250 164.440 ;
        RECT 101.310 162.860 101.540 164.440 ;
        RECT 74.860 155.570 75.090 157.150 ;
        RECT 80.150 155.570 80.380 157.150 ;
        RECT 85.440 155.570 85.670 157.150 ;
        RECT 90.730 155.570 90.960 157.150 ;
        RECT 96.020 155.570 96.250 157.150 ;
        RECT 101.310 155.570 101.540 157.150 ;
        RECT 74.860 150.100 75.090 151.680 ;
        RECT 80.150 150.100 80.380 151.680 ;
        RECT 85.440 150.100 85.670 151.680 ;
        RECT 90.730 150.100 90.960 151.680 ;
        RECT 96.020 150.100 96.250 151.680 ;
        RECT 101.310 150.100 101.540 151.680 ;
        RECT 74.860 144.630 75.090 146.210 ;
        RECT 80.150 144.630 80.380 146.210 ;
        RECT 85.440 144.630 85.670 146.210 ;
        RECT 90.730 144.630 90.960 146.210 ;
        RECT 96.020 144.630 96.250 146.210 ;
        RECT 101.310 144.630 101.540 146.210 ;
        RECT 74.860 139.160 75.090 140.740 ;
        RECT 80.150 139.160 80.380 140.740 ;
        RECT 85.440 139.160 85.670 140.740 ;
        RECT 90.730 139.160 90.960 140.740 ;
        RECT 96.020 139.160 96.250 140.740 ;
        RECT 101.310 139.160 101.540 140.740 ;
        RECT 74.860 133.690 75.090 135.270 ;
        RECT 80.150 133.690 80.380 135.270 ;
        RECT 85.440 133.690 85.670 135.270 ;
        RECT 90.730 133.690 90.960 135.270 ;
        RECT 96.020 133.690 96.250 135.270 ;
        RECT 101.310 133.690 101.540 135.270 ;
        RECT 74.860 126.390 75.090 127.970 ;
        RECT 80.150 126.390 80.380 127.970 ;
        RECT 85.440 126.390 85.670 127.970 ;
        RECT 90.730 126.390 90.960 127.970 ;
        RECT 96.020 126.390 96.250 127.970 ;
        RECT 101.310 126.390 101.540 127.970 ;
        RECT 74.860 120.920 75.090 122.500 ;
        RECT 80.150 120.920 80.380 122.500 ;
        RECT 85.440 120.920 85.670 122.500 ;
        RECT 90.730 120.920 90.960 122.500 ;
        RECT 96.020 120.920 96.250 122.500 ;
        RECT 101.310 120.920 101.540 122.500 ;
        RECT 74.860 115.450 75.090 117.030 ;
        RECT 80.150 115.450 80.380 117.030 ;
        RECT 85.440 115.450 85.670 117.030 ;
        RECT 90.730 115.450 90.960 117.030 ;
        RECT 96.020 115.450 96.250 117.030 ;
        RECT 101.310 115.450 101.540 117.030 ;
        RECT 74.860 109.980 75.090 111.560 ;
        RECT 80.150 109.980 80.380 111.560 ;
        RECT 85.440 109.980 85.670 111.560 ;
        RECT 90.730 109.980 90.960 111.560 ;
        RECT 96.020 109.980 96.250 111.560 ;
        RECT 101.310 109.980 101.540 111.560 ;
        RECT 74.860 104.510 75.090 106.090 ;
        RECT 80.150 104.510 80.380 106.090 ;
        RECT 85.440 104.510 85.670 106.090 ;
        RECT 90.730 104.510 90.960 106.090 ;
        RECT 96.020 104.510 96.250 106.090 ;
        RECT 101.310 104.510 101.540 106.090 ;
        RECT 74.860 97.070 75.090 98.650 ;
        RECT 80.150 97.070 80.380 98.650 ;
        RECT 85.440 97.070 85.670 98.650 ;
        RECT 90.730 97.070 90.960 98.650 ;
        RECT 96.020 97.070 96.250 98.650 ;
        RECT 101.310 97.070 101.540 98.650 ;
        RECT 74.860 91.600 75.090 93.180 ;
        RECT 80.150 91.600 80.380 93.180 ;
        RECT 85.440 91.600 85.670 93.180 ;
        RECT 90.730 91.600 90.960 93.180 ;
        RECT 96.020 91.600 96.250 93.180 ;
        RECT 101.310 91.600 101.540 93.180 ;
        RECT 74.860 86.130 75.090 87.710 ;
        RECT 80.150 86.130 80.380 87.710 ;
        RECT 85.440 86.130 85.670 87.710 ;
        RECT 90.730 86.130 90.960 87.710 ;
        RECT 96.020 86.130 96.250 87.710 ;
        RECT 101.310 86.130 101.540 87.710 ;
        RECT 74.860 80.660 75.090 82.240 ;
        RECT 80.150 80.660 80.380 82.240 ;
        RECT 85.440 80.660 85.670 82.240 ;
        RECT 90.730 80.660 90.960 82.240 ;
        RECT 96.020 80.660 96.250 82.240 ;
        RECT 101.310 80.660 101.540 82.240 ;
        RECT 74.860 75.190 75.090 76.770 ;
        RECT 80.150 75.190 80.380 76.770 ;
        RECT 85.440 75.190 85.670 76.770 ;
        RECT 90.730 75.190 90.960 76.770 ;
        RECT 96.020 75.190 96.250 76.770 ;
        RECT 101.310 75.190 101.540 76.770 ;
        RECT 74.910 67.790 75.140 69.370 ;
        RECT 80.200 67.790 80.430 69.370 ;
        RECT 85.490 67.790 85.720 69.370 ;
        RECT 90.780 67.790 91.010 69.370 ;
        RECT 96.070 67.790 96.300 69.370 ;
        RECT 101.360 67.790 101.590 69.370 ;
        RECT 74.910 62.320 75.140 63.900 ;
        RECT 80.200 62.320 80.430 63.900 ;
        RECT 85.490 62.320 85.720 63.900 ;
        RECT 90.780 62.320 91.010 63.900 ;
        RECT 96.070 62.320 96.300 63.900 ;
        RECT 101.360 62.320 101.590 63.900 ;
        RECT 74.910 56.850 75.140 58.430 ;
        RECT 80.200 56.850 80.430 58.430 ;
        RECT 85.490 56.850 85.720 58.430 ;
        RECT 90.780 56.850 91.010 58.430 ;
        RECT 96.070 56.850 96.300 58.430 ;
        RECT 101.360 56.850 101.590 58.430 ;
        RECT 74.910 51.380 75.140 52.960 ;
        RECT 80.200 51.380 80.430 52.960 ;
        RECT 85.490 51.380 85.720 52.960 ;
        RECT 90.780 51.380 91.010 52.960 ;
        RECT 96.070 51.380 96.300 52.960 ;
        RECT 101.360 51.380 101.590 52.960 ;
        RECT 74.910 45.910 75.140 47.490 ;
        RECT 80.200 45.910 80.430 47.490 ;
        RECT 85.490 45.910 85.720 47.490 ;
        RECT 90.780 45.910 91.010 47.490 ;
        RECT 96.070 45.910 96.300 47.490 ;
        RECT 101.360 45.910 101.590 47.490 ;
        RECT 75.000 38.250 75.230 39.830 ;
        RECT 80.290 38.250 80.520 39.830 ;
        RECT 85.580 38.250 85.810 39.830 ;
        RECT 90.870 38.250 91.100 39.830 ;
        RECT 96.160 38.250 96.390 39.830 ;
        RECT 101.450 38.250 101.680 39.830 ;
        RECT 75.000 32.780 75.230 34.360 ;
        RECT 80.290 32.780 80.520 34.360 ;
        RECT 85.580 32.780 85.810 34.360 ;
        RECT 90.870 32.780 91.100 34.360 ;
        RECT 96.160 32.780 96.390 34.360 ;
        RECT 101.450 32.780 101.680 34.360 ;
        RECT 75.000 27.310 75.230 28.890 ;
        RECT 80.290 27.310 80.520 28.890 ;
        RECT 85.580 27.310 85.810 28.890 ;
        RECT 90.870 27.310 91.100 28.890 ;
        RECT 96.160 27.310 96.390 28.890 ;
        RECT 101.450 27.310 101.680 28.890 ;
        RECT 75.000 21.840 75.230 23.420 ;
        RECT 80.290 21.840 80.520 23.420 ;
        RECT 85.580 21.840 85.810 23.420 ;
        RECT 90.870 21.840 91.100 23.420 ;
        RECT 96.160 21.840 96.390 23.420 ;
        RECT 101.450 21.840 101.680 23.420 ;
        RECT 71.080 -15.670 72.560 16.890 ;
        RECT 75.000 16.370 75.230 17.950 ;
        RECT 80.290 16.370 80.520 17.950 ;
        RECT 85.580 16.370 85.810 17.950 ;
        RECT 90.870 16.370 91.100 17.950 ;
        RECT 96.160 16.370 96.390 17.950 ;
        RECT 101.450 16.370 101.680 17.950 ;
        RECT 102.800 17.910 106.000 202.690 ;
        RECT 103.740 -15.670 105.220 17.910 ;
        RECT 135.410 17.650 138.440 213.850 ;
        RECT 167.950 18.940 171.390 214.110 ;
        RECT 204.920 213.850 205.150 215.430 ;
        RECT 210.210 213.850 210.440 215.430 ;
        RECT 215.500 213.850 215.730 215.430 ;
        RECT 220.790 213.850 221.020 215.430 ;
        RECT 226.080 213.850 226.310 215.430 ;
        RECT 231.370 213.850 231.600 215.430 ;
        RECT 237.860 213.960 238.090 215.540 ;
        RECT 243.150 213.960 243.380 215.540 ;
        RECT 248.440 213.960 248.670 215.540 ;
        RECT 253.730 213.960 253.960 215.540 ;
        RECT 259.020 213.960 259.250 215.540 ;
        RECT 264.310 213.960 264.540 215.540 ;
        RECT 270.430 214.030 270.660 215.610 ;
        RECT 275.720 214.030 275.950 215.610 ;
        RECT 281.010 214.030 281.240 215.610 ;
        RECT 286.300 214.030 286.530 215.610 ;
        RECT 291.590 214.030 291.820 215.610 ;
        RECT 296.880 214.030 297.110 215.610 ;
        RECT 312.510 214.620 312.740 215.600 ;
        RECT 315.800 214.620 316.030 215.600 ;
        RECT 319.090 214.620 319.320 215.600 ;
        RECT 322.380 214.620 322.610 215.600 ;
        RECT 325.670 214.620 325.900 215.600 ;
        RECT 328.960 214.620 329.190 215.600 ;
        RECT 334.770 214.630 335.000 215.610 ;
        RECT 341.350 214.630 341.580 215.610 ;
        RECT 347.930 214.630 348.160 215.610 ;
        RECT 350.520 214.700 350.750 215.680 ;
        RECT 353.810 214.700 354.040 215.680 ;
        RECT 357.100 214.700 357.330 215.680 ;
        RECT 360.390 214.700 360.620 215.680 ;
        RECT 363.680 214.700 363.910 215.680 ;
        RECT 366.970 214.700 367.200 215.680 ;
        RECT 200.460 27.940 203.690 212.830 ;
        RECT 204.920 208.380 205.150 209.960 ;
        RECT 210.210 208.380 210.440 209.960 ;
        RECT 215.500 208.380 215.730 209.960 ;
        RECT 220.790 208.380 221.020 209.960 ;
        RECT 226.080 208.380 226.310 209.960 ;
        RECT 231.370 208.380 231.600 209.960 ;
        RECT 204.920 202.910 205.150 204.490 ;
        RECT 210.210 202.910 210.440 204.490 ;
        RECT 215.500 202.910 215.730 204.490 ;
        RECT 220.790 202.910 221.020 204.490 ;
        RECT 226.080 202.910 226.310 204.490 ;
        RECT 231.370 202.910 231.600 204.490 ;
        RECT 204.920 197.440 205.150 199.020 ;
        RECT 210.210 197.440 210.440 199.020 ;
        RECT 215.500 197.440 215.730 199.020 ;
        RECT 220.790 197.440 221.020 199.020 ;
        RECT 226.080 197.440 226.310 199.020 ;
        RECT 231.370 197.440 231.600 199.020 ;
        RECT 204.920 191.970 205.150 193.550 ;
        RECT 210.210 191.970 210.440 193.550 ;
        RECT 215.500 191.970 215.730 193.550 ;
        RECT 220.790 191.970 221.020 193.550 ;
        RECT 226.080 191.970 226.310 193.550 ;
        RECT 231.370 191.970 231.600 193.550 ;
        RECT 204.920 184.770 205.150 186.350 ;
        RECT 210.210 184.770 210.440 186.350 ;
        RECT 215.500 184.770 215.730 186.350 ;
        RECT 220.790 184.770 221.020 186.350 ;
        RECT 226.080 184.770 226.310 186.350 ;
        RECT 231.370 184.770 231.600 186.350 ;
        RECT 204.920 179.300 205.150 180.880 ;
        RECT 210.210 179.300 210.440 180.880 ;
        RECT 215.500 179.300 215.730 180.880 ;
        RECT 220.790 179.300 221.020 180.880 ;
        RECT 226.080 179.300 226.310 180.880 ;
        RECT 231.370 179.300 231.600 180.880 ;
        RECT 204.920 173.830 205.150 175.410 ;
        RECT 210.210 173.830 210.440 175.410 ;
        RECT 215.500 173.830 215.730 175.410 ;
        RECT 220.790 173.830 221.020 175.410 ;
        RECT 226.080 173.830 226.310 175.410 ;
        RECT 231.370 173.830 231.600 175.410 ;
        RECT 204.920 168.360 205.150 169.940 ;
        RECT 210.210 168.360 210.440 169.940 ;
        RECT 215.500 168.360 215.730 169.940 ;
        RECT 220.790 168.360 221.020 169.940 ;
        RECT 226.080 168.360 226.310 169.940 ;
        RECT 231.370 168.360 231.600 169.940 ;
        RECT 204.920 162.890 205.150 164.470 ;
        RECT 210.210 162.890 210.440 164.470 ;
        RECT 215.500 162.890 215.730 164.470 ;
        RECT 220.790 162.890 221.020 164.470 ;
        RECT 226.080 162.890 226.310 164.470 ;
        RECT 231.370 162.890 231.600 164.470 ;
        RECT 204.920 155.600 205.150 157.180 ;
        RECT 210.210 155.600 210.440 157.180 ;
        RECT 215.500 155.600 215.730 157.180 ;
        RECT 220.790 155.600 221.020 157.180 ;
        RECT 226.080 155.600 226.310 157.180 ;
        RECT 231.370 155.600 231.600 157.180 ;
        RECT 204.920 150.130 205.150 151.710 ;
        RECT 210.210 150.130 210.440 151.710 ;
        RECT 215.500 150.130 215.730 151.710 ;
        RECT 220.790 150.130 221.020 151.710 ;
        RECT 226.080 150.130 226.310 151.710 ;
        RECT 231.370 150.130 231.600 151.710 ;
        RECT 204.920 144.660 205.150 146.240 ;
        RECT 210.210 144.660 210.440 146.240 ;
        RECT 215.500 144.660 215.730 146.240 ;
        RECT 220.790 144.660 221.020 146.240 ;
        RECT 226.080 144.660 226.310 146.240 ;
        RECT 231.370 144.660 231.600 146.240 ;
        RECT 204.920 139.190 205.150 140.770 ;
        RECT 210.210 139.190 210.440 140.770 ;
        RECT 215.500 139.190 215.730 140.770 ;
        RECT 220.790 139.190 221.020 140.770 ;
        RECT 226.080 139.190 226.310 140.770 ;
        RECT 231.370 139.190 231.600 140.770 ;
        RECT 204.920 133.720 205.150 135.300 ;
        RECT 210.210 133.720 210.440 135.300 ;
        RECT 215.500 133.720 215.730 135.300 ;
        RECT 220.790 133.720 221.020 135.300 ;
        RECT 226.080 133.720 226.310 135.300 ;
        RECT 231.370 133.720 231.600 135.300 ;
        RECT 204.920 126.420 205.150 128.000 ;
        RECT 210.210 126.420 210.440 128.000 ;
        RECT 215.500 126.420 215.730 128.000 ;
        RECT 220.790 126.420 221.020 128.000 ;
        RECT 226.080 126.420 226.310 128.000 ;
        RECT 231.370 126.420 231.600 128.000 ;
        RECT 204.920 120.950 205.150 122.530 ;
        RECT 210.210 120.950 210.440 122.530 ;
        RECT 215.500 120.950 215.730 122.530 ;
        RECT 220.790 120.950 221.020 122.530 ;
        RECT 226.080 120.950 226.310 122.530 ;
        RECT 231.370 120.950 231.600 122.530 ;
        RECT 204.920 115.480 205.150 117.060 ;
        RECT 210.210 115.480 210.440 117.060 ;
        RECT 215.500 115.480 215.730 117.060 ;
        RECT 220.790 115.480 221.020 117.060 ;
        RECT 226.080 115.480 226.310 117.060 ;
        RECT 231.370 115.480 231.600 117.060 ;
        RECT 204.920 110.010 205.150 111.590 ;
        RECT 210.210 110.010 210.440 111.590 ;
        RECT 215.500 110.010 215.730 111.590 ;
        RECT 220.790 110.010 221.020 111.590 ;
        RECT 226.080 110.010 226.310 111.590 ;
        RECT 231.370 110.010 231.600 111.590 ;
        RECT 204.920 104.540 205.150 106.120 ;
        RECT 210.210 104.540 210.440 106.120 ;
        RECT 215.500 104.540 215.730 106.120 ;
        RECT 220.790 104.540 221.020 106.120 ;
        RECT 226.080 104.540 226.310 106.120 ;
        RECT 231.370 104.540 231.600 106.120 ;
        RECT 204.920 97.100 205.150 98.680 ;
        RECT 210.210 97.100 210.440 98.680 ;
        RECT 215.500 97.100 215.730 98.680 ;
        RECT 220.790 97.100 221.020 98.680 ;
        RECT 226.080 97.100 226.310 98.680 ;
        RECT 231.370 97.100 231.600 98.680 ;
        RECT 204.920 91.630 205.150 93.210 ;
        RECT 210.210 91.630 210.440 93.210 ;
        RECT 215.500 91.630 215.730 93.210 ;
        RECT 220.790 91.630 221.020 93.210 ;
        RECT 226.080 91.630 226.310 93.210 ;
        RECT 231.370 91.630 231.600 93.210 ;
        RECT 204.920 86.160 205.150 87.740 ;
        RECT 210.210 86.160 210.440 87.740 ;
        RECT 215.500 86.160 215.730 87.740 ;
        RECT 220.790 86.160 221.020 87.740 ;
        RECT 226.080 86.160 226.310 87.740 ;
        RECT 231.370 86.160 231.600 87.740 ;
        RECT 204.920 80.690 205.150 82.270 ;
        RECT 210.210 80.690 210.440 82.270 ;
        RECT 215.500 80.690 215.730 82.270 ;
        RECT 220.790 80.690 221.020 82.270 ;
        RECT 226.080 80.690 226.310 82.270 ;
        RECT 231.370 80.690 231.600 82.270 ;
        RECT 204.920 75.220 205.150 76.800 ;
        RECT 210.210 75.220 210.440 76.800 ;
        RECT 215.500 75.220 215.730 76.800 ;
        RECT 220.790 75.220 221.020 76.800 ;
        RECT 226.080 75.220 226.310 76.800 ;
        RECT 231.370 75.220 231.600 76.800 ;
        RECT 204.970 67.820 205.200 69.400 ;
        RECT 210.260 67.820 210.490 69.400 ;
        RECT 215.550 67.820 215.780 69.400 ;
        RECT 220.840 67.820 221.070 69.400 ;
        RECT 226.130 67.820 226.360 69.400 ;
        RECT 231.420 67.820 231.650 69.400 ;
        RECT 204.970 62.350 205.200 63.930 ;
        RECT 210.260 62.350 210.490 63.930 ;
        RECT 215.550 62.350 215.780 63.930 ;
        RECT 220.840 62.350 221.070 63.930 ;
        RECT 226.130 62.350 226.360 63.930 ;
        RECT 231.420 62.350 231.650 63.930 ;
        RECT 204.970 56.880 205.200 58.460 ;
        RECT 210.260 56.880 210.490 58.460 ;
        RECT 215.550 56.880 215.780 58.460 ;
        RECT 220.840 56.880 221.070 58.460 ;
        RECT 226.130 56.880 226.360 58.460 ;
        RECT 231.420 56.880 231.650 58.460 ;
        RECT 204.970 51.410 205.200 52.990 ;
        RECT 210.260 51.410 210.490 52.990 ;
        RECT 215.550 51.410 215.780 52.990 ;
        RECT 220.840 51.410 221.070 52.990 ;
        RECT 226.130 51.410 226.360 52.990 ;
        RECT 231.420 51.410 231.650 52.990 ;
        RECT 204.970 45.940 205.200 47.520 ;
        RECT 210.260 45.940 210.490 47.520 ;
        RECT 215.550 45.940 215.780 47.520 ;
        RECT 220.840 45.940 221.070 47.520 ;
        RECT 226.130 45.940 226.360 47.520 ;
        RECT 231.420 45.940 231.650 47.520 ;
        RECT 205.060 38.280 205.290 39.860 ;
        RECT 210.350 38.280 210.580 39.860 ;
        RECT 215.640 38.280 215.870 39.860 ;
        RECT 220.930 38.280 221.160 39.860 ;
        RECT 226.220 38.280 226.450 39.860 ;
        RECT 231.510 38.280 231.740 39.860 ;
        RECT 205.060 32.810 205.290 34.390 ;
        RECT 210.350 32.810 210.580 34.390 ;
        RECT 215.640 32.810 215.870 34.390 ;
        RECT 220.930 32.810 221.160 34.390 ;
        RECT 226.220 32.810 226.450 34.390 ;
        RECT 231.510 32.810 231.740 34.390 ;
        RECT 201.820 24.530 202.570 27.940 ;
        RECT 205.060 27.340 205.290 28.920 ;
        RECT 210.350 27.340 210.580 28.920 ;
        RECT 215.640 27.340 215.870 28.920 ;
        RECT 220.930 27.340 221.160 28.920 ;
        RECT 226.220 27.340 226.450 28.920 ;
        RECT 231.510 27.340 231.740 28.920 ;
        RECT 232.980 28.420 236.460 212.120 ;
        RECT 237.860 208.490 238.090 210.070 ;
        RECT 243.150 208.490 243.380 210.070 ;
        RECT 248.440 208.490 248.670 210.070 ;
        RECT 253.730 208.490 253.960 210.070 ;
        RECT 259.020 208.490 259.250 210.070 ;
        RECT 264.310 208.490 264.540 210.070 ;
        RECT 237.860 203.020 238.090 204.600 ;
        RECT 243.150 203.020 243.380 204.600 ;
        RECT 248.440 203.020 248.670 204.600 ;
        RECT 253.730 203.020 253.960 204.600 ;
        RECT 259.020 203.020 259.250 204.600 ;
        RECT 264.310 203.020 264.540 204.600 ;
        RECT 237.860 197.550 238.090 199.130 ;
        RECT 243.150 197.550 243.380 199.130 ;
        RECT 248.440 197.550 248.670 199.130 ;
        RECT 253.730 197.550 253.960 199.130 ;
        RECT 259.020 197.550 259.250 199.130 ;
        RECT 264.310 197.550 264.540 199.130 ;
        RECT 237.860 192.080 238.090 193.660 ;
        RECT 243.150 192.080 243.380 193.660 ;
        RECT 248.440 192.080 248.670 193.660 ;
        RECT 253.730 192.080 253.960 193.660 ;
        RECT 259.020 192.080 259.250 193.660 ;
        RECT 264.310 192.080 264.540 193.660 ;
        RECT 237.860 184.880 238.090 186.460 ;
        RECT 243.150 184.880 243.380 186.460 ;
        RECT 248.440 184.880 248.670 186.460 ;
        RECT 253.730 184.880 253.960 186.460 ;
        RECT 259.020 184.880 259.250 186.460 ;
        RECT 264.310 184.880 264.540 186.460 ;
        RECT 237.860 179.410 238.090 180.990 ;
        RECT 243.150 179.410 243.380 180.990 ;
        RECT 248.440 179.410 248.670 180.990 ;
        RECT 253.730 179.410 253.960 180.990 ;
        RECT 259.020 179.410 259.250 180.990 ;
        RECT 264.310 179.410 264.540 180.990 ;
        RECT 237.860 173.940 238.090 175.520 ;
        RECT 243.150 173.940 243.380 175.520 ;
        RECT 248.440 173.940 248.670 175.520 ;
        RECT 253.730 173.940 253.960 175.520 ;
        RECT 259.020 173.940 259.250 175.520 ;
        RECT 264.310 173.940 264.540 175.520 ;
        RECT 237.860 168.470 238.090 170.050 ;
        RECT 243.150 168.470 243.380 170.050 ;
        RECT 248.440 168.470 248.670 170.050 ;
        RECT 253.730 168.470 253.960 170.050 ;
        RECT 259.020 168.470 259.250 170.050 ;
        RECT 264.310 168.470 264.540 170.050 ;
        RECT 237.860 163.000 238.090 164.580 ;
        RECT 243.150 163.000 243.380 164.580 ;
        RECT 248.440 163.000 248.670 164.580 ;
        RECT 253.730 163.000 253.960 164.580 ;
        RECT 259.020 163.000 259.250 164.580 ;
        RECT 264.310 163.000 264.540 164.580 ;
        RECT 237.860 155.710 238.090 157.290 ;
        RECT 243.150 155.710 243.380 157.290 ;
        RECT 248.440 155.710 248.670 157.290 ;
        RECT 253.730 155.710 253.960 157.290 ;
        RECT 259.020 155.710 259.250 157.290 ;
        RECT 264.310 155.710 264.540 157.290 ;
        RECT 237.860 150.240 238.090 151.820 ;
        RECT 243.150 150.240 243.380 151.820 ;
        RECT 248.440 150.240 248.670 151.820 ;
        RECT 253.730 150.240 253.960 151.820 ;
        RECT 259.020 150.240 259.250 151.820 ;
        RECT 264.310 150.240 264.540 151.820 ;
        RECT 237.860 144.770 238.090 146.350 ;
        RECT 243.150 144.770 243.380 146.350 ;
        RECT 248.440 144.770 248.670 146.350 ;
        RECT 253.730 144.770 253.960 146.350 ;
        RECT 259.020 144.770 259.250 146.350 ;
        RECT 264.310 144.770 264.540 146.350 ;
        RECT 237.860 139.300 238.090 140.880 ;
        RECT 243.150 139.300 243.380 140.880 ;
        RECT 248.440 139.300 248.670 140.880 ;
        RECT 253.730 139.300 253.960 140.880 ;
        RECT 259.020 139.300 259.250 140.880 ;
        RECT 264.310 139.300 264.540 140.880 ;
        RECT 237.860 133.830 238.090 135.410 ;
        RECT 243.150 133.830 243.380 135.410 ;
        RECT 248.440 133.830 248.670 135.410 ;
        RECT 253.730 133.830 253.960 135.410 ;
        RECT 259.020 133.830 259.250 135.410 ;
        RECT 264.310 133.830 264.540 135.410 ;
        RECT 237.860 126.530 238.090 128.110 ;
        RECT 243.150 126.530 243.380 128.110 ;
        RECT 248.440 126.530 248.670 128.110 ;
        RECT 253.730 126.530 253.960 128.110 ;
        RECT 259.020 126.530 259.250 128.110 ;
        RECT 264.310 126.530 264.540 128.110 ;
        RECT 237.860 121.060 238.090 122.640 ;
        RECT 243.150 121.060 243.380 122.640 ;
        RECT 248.440 121.060 248.670 122.640 ;
        RECT 253.730 121.060 253.960 122.640 ;
        RECT 259.020 121.060 259.250 122.640 ;
        RECT 264.310 121.060 264.540 122.640 ;
        RECT 237.860 115.590 238.090 117.170 ;
        RECT 243.150 115.590 243.380 117.170 ;
        RECT 248.440 115.590 248.670 117.170 ;
        RECT 253.730 115.590 253.960 117.170 ;
        RECT 259.020 115.590 259.250 117.170 ;
        RECT 264.310 115.590 264.540 117.170 ;
        RECT 237.860 110.120 238.090 111.700 ;
        RECT 243.150 110.120 243.380 111.700 ;
        RECT 248.440 110.120 248.670 111.700 ;
        RECT 253.730 110.120 253.960 111.700 ;
        RECT 259.020 110.120 259.250 111.700 ;
        RECT 264.310 110.120 264.540 111.700 ;
        RECT 237.860 104.650 238.090 106.230 ;
        RECT 243.150 104.650 243.380 106.230 ;
        RECT 248.440 104.650 248.670 106.230 ;
        RECT 253.730 104.650 253.960 106.230 ;
        RECT 259.020 104.650 259.250 106.230 ;
        RECT 264.310 104.650 264.540 106.230 ;
        RECT 237.860 97.210 238.090 98.790 ;
        RECT 243.150 97.210 243.380 98.790 ;
        RECT 248.440 97.210 248.670 98.790 ;
        RECT 253.730 97.210 253.960 98.790 ;
        RECT 259.020 97.210 259.250 98.790 ;
        RECT 264.310 97.210 264.540 98.790 ;
        RECT 237.860 91.740 238.090 93.320 ;
        RECT 243.150 91.740 243.380 93.320 ;
        RECT 248.440 91.740 248.670 93.320 ;
        RECT 253.730 91.740 253.960 93.320 ;
        RECT 259.020 91.740 259.250 93.320 ;
        RECT 264.310 91.740 264.540 93.320 ;
        RECT 237.860 86.270 238.090 87.850 ;
        RECT 243.150 86.270 243.380 87.850 ;
        RECT 248.440 86.270 248.670 87.850 ;
        RECT 253.730 86.270 253.960 87.850 ;
        RECT 259.020 86.270 259.250 87.850 ;
        RECT 264.310 86.270 264.540 87.850 ;
        RECT 237.860 80.800 238.090 82.380 ;
        RECT 243.150 80.800 243.380 82.380 ;
        RECT 248.440 80.800 248.670 82.380 ;
        RECT 253.730 80.800 253.960 82.380 ;
        RECT 259.020 80.800 259.250 82.380 ;
        RECT 264.310 80.800 264.540 82.380 ;
        RECT 237.860 75.330 238.090 76.910 ;
        RECT 243.150 75.330 243.380 76.910 ;
        RECT 248.440 75.330 248.670 76.910 ;
        RECT 253.730 75.330 253.960 76.910 ;
        RECT 259.020 75.330 259.250 76.910 ;
        RECT 264.310 75.330 264.540 76.910 ;
        RECT 237.910 67.930 238.140 69.510 ;
        RECT 243.200 67.930 243.430 69.510 ;
        RECT 248.490 67.930 248.720 69.510 ;
        RECT 253.780 67.930 254.010 69.510 ;
        RECT 259.070 67.930 259.300 69.510 ;
        RECT 264.360 67.930 264.590 69.510 ;
        RECT 237.910 62.460 238.140 64.040 ;
        RECT 243.200 62.460 243.430 64.040 ;
        RECT 248.490 62.460 248.720 64.040 ;
        RECT 253.780 62.460 254.010 64.040 ;
        RECT 259.070 62.460 259.300 64.040 ;
        RECT 264.360 62.460 264.590 64.040 ;
        RECT 237.910 56.990 238.140 58.570 ;
        RECT 243.200 56.990 243.430 58.570 ;
        RECT 248.490 56.990 248.720 58.570 ;
        RECT 253.780 56.990 254.010 58.570 ;
        RECT 259.070 56.990 259.300 58.570 ;
        RECT 264.360 56.990 264.590 58.570 ;
        RECT 237.910 51.520 238.140 53.100 ;
        RECT 243.200 51.520 243.430 53.100 ;
        RECT 248.490 51.520 248.720 53.100 ;
        RECT 253.780 51.520 254.010 53.100 ;
        RECT 259.070 51.520 259.300 53.100 ;
        RECT 264.360 51.520 264.590 53.100 ;
        RECT 237.910 46.050 238.140 47.630 ;
        RECT 243.200 46.050 243.430 47.630 ;
        RECT 248.490 46.050 248.720 47.630 ;
        RECT 253.780 46.050 254.010 47.630 ;
        RECT 259.070 46.050 259.300 47.630 ;
        RECT 264.360 46.050 264.590 47.630 ;
        RECT 238.000 38.390 238.230 39.970 ;
        RECT 243.290 38.390 243.520 39.970 ;
        RECT 248.580 38.390 248.810 39.970 ;
        RECT 253.870 38.390 254.100 39.970 ;
        RECT 259.160 38.390 259.390 39.970 ;
        RECT 264.450 38.390 264.680 39.970 ;
        RECT 238.000 32.920 238.230 34.500 ;
        RECT 243.290 32.920 243.520 34.500 ;
        RECT 248.580 32.920 248.810 34.500 ;
        RECT 253.870 32.920 254.100 34.500 ;
        RECT 259.160 32.920 259.390 34.500 ;
        RECT 264.450 32.920 264.680 34.500 ;
        RECT 238.000 28.420 238.230 29.030 ;
        RECT 232.980 27.390 238.680 28.420 ;
        RECT 243.290 27.450 243.520 29.030 ;
        RECT 248.580 27.450 248.810 29.030 ;
        RECT 253.870 27.450 254.100 29.030 ;
        RECT 259.160 27.450 259.390 29.030 ;
        RECT 264.450 27.450 264.680 29.030 ;
        RECT 265.680 28.600 269.160 211.970 ;
        RECT 270.430 208.560 270.660 210.140 ;
        RECT 275.720 208.560 275.950 210.140 ;
        RECT 281.010 208.560 281.240 210.140 ;
        RECT 286.300 208.560 286.530 210.140 ;
        RECT 291.590 208.560 291.820 210.140 ;
        RECT 296.880 208.560 297.110 210.140 ;
        RECT 297.650 206.460 299.670 209.760 ;
        RECT 310.740 208.020 311.800 213.500 ;
        RECT 312.510 211.150 312.740 212.130 ;
        RECT 315.800 211.150 316.030 212.130 ;
        RECT 319.090 211.150 319.320 212.130 ;
        RECT 322.380 211.150 322.610 212.130 ;
        RECT 325.670 211.150 325.900 212.130 ;
        RECT 328.960 211.150 329.190 212.130 ;
        RECT 329.710 212.040 330.770 213.510 ;
        RECT 348.750 212.340 349.810 213.580 ;
        RECT 368.050 212.710 369.750 215.010 ;
        RECT 442.710 213.330 449.070 218.420 ;
        RECT 310.580 206.460 311.800 208.020 ;
        RECT 312.510 207.680 312.740 208.660 ;
        RECT 315.800 207.680 316.030 208.660 ;
        RECT 319.090 207.680 319.320 208.660 ;
        RECT 322.380 207.680 322.610 208.660 ;
        RECT 325.670 207.680 325.900 208.660 ;
        RECT 328.960 207.680 329.190 208.660 ;
        RECT 297.650 205.200 311.800 206.460 ;
        RECT 270.430 203.090 270.660 204.670 ;
        RECT 275.720 203.090 275.950 204.670 ;
        RECT 281.010 203.090 281.240 204.670 ;
        RECT 286.300 203.090 286.530 204.670 ;
        RECT 291.590 203.090 291.820 204.670 ;
        RECT 296.880 203.090 297.110 204.670 ;
        RECT 297.650 200.330 300.060 205.200 ;
        RECT 270.430 197.620 270.660 199.200 ;
        RECT 275.720 197.620 275.950 199.200 ;
        RECT 281.010 197.620 281.240 199.200 ;
        RECT 286.300 197.620 286.530 199.200 ;
        RECT 291.590 197.620 291.820 199.200 ;
        RECT 296.880 197.620 297.110 199.200 ;
        RECT 270.430 192.150 270.660 193.730 ;
        RECT 275.720 192.150 275.950 193.730 ;
        RECT 281.010 192.150 281.240 193.730 ;
        RECT 286.300 192.150 286.530 193.730 ;
        RECT 291.590 192.150 291.820 193.730 ;
        RECT 296.880 192.150 297.110 193.730 ;
        RECT 270.430 184.950 270.660 186.530 ;
        RECT 275.720 184.950 275.950 186.530 ;
        RECT 281.010 184.950 281.240 186.530 ;
        RECT 286.300 184.950 286.530 186.530 ;
        RECT 291.590 184.950 291.820 186.530 ;
        RECT 296.880 184.950 297.110 186.530 ;
        RECT 270.430 179.480 270.660 181.060 ;
        RECT 275.720 179.480 275.950 181.060 ;
        RECT 281.010 179.480 281.240 181.060 ;
        RECT 286.300 179.480 286.530 181.060 ;
        RECT 291.590 179.480 291.820 181.060 ;
        RECT 296.880 179.480 297.110 181.060 ;
        RECT 298.400 180.420 300.060 200.330 ;
        RECT 310.580 203.950 311.800 205.200 ;
        RECT 312.510 204.210 312.740 205.190 ;
        RECT 315.800 204.210 316.030 205.190 ;
        RECT 319.090 204.210 319.320 205.190 ;
        RECT 322.380 204.210 322.610 205.190 ;
        RECT 325.670 204.210 325.900 205.190 ;
        RECT 328.960 204.210 329.190 205.190 ;
        RECT 329.710 203.960 331.140 212.040 ;
        RECT 334.770 211.160 335.000 212.140 ;
        RECT 341.350 211.160 341.580 212.140 ;
        RECT 347.930 211.160 348.160 212.140 ;
        RECT 334.770 207.690 335.000 208.670 ;
        RECT 341.350 207.690 341.580 208.670 ;
        RECT 347.930 207.690 348.160 208.670 ;
        RECT 334.770 204.220 335.000 205.200 ;
        RECT 341.350 204.220 341.580 205.200 ;
        RECT 347.930 204.220 348.160 205.200 ;
        RECT 310.580 198.110 311.480 203.950 ;
        RECT 312.510 200.740 312.740 201.720 ;
        RECT 315.800 200.740 316.030 201.720 ;
        RECT 319.090 200.740 319.320 201.720 ;
        RECT 322.380 200.740 322.610 201.720 ;
        RECT 325.670 200.740 325.900 201.720 ;
        RECT 328.960 200.740 329.190 201.720 ;
        RECT 329.760 198.110 331.140 203.960 ;
        RECT 334.770 200.750 335.000 201.730 ;
        RECT 341.350 200.750 341.580 201.730 ;
        RECT 347.930 200.750 348.160 201.730 ;
        RECT 348.540 198.110 349.920 212.340 ;
        RECT 350.520 211.230 350.750 212.210 ;
        RECT 353.810 211.230 354.040 212.210 ;
        RECT 357.100 211.230 357.330 212.210 ;
        RECT 360.390 211.230 360.620 212.210 ;
        RECT 363.680 211.230 363.910 212.210 ;
        RECT 366.970 211.230 367.200 212.210 ;
        RECT 350.520 207.760 350.750 208.740 ;
        RECT 353.810 207.760 354.040 208.740 ;
        RECT 357.100 207.760 357.330 208.740 ;
        RECT 360.390 207.760 360.620 208.740 ;
        RECT 363.680 207.760 363.910 208.740 ;
        RECT 366.970 207.760 367.200 208.740 ;
        RECT 350.520 204.290 350.750 205.270 ;
        RECT 353.810 204.290 354.040 205.270 ;
        RECT 357.100 204.290 357.330 205.270 ;
        RECT 360.390 204.290 360.620 205.270 ;
        RECT 363.680 204.290 363.910 205.270 ;
        RECT 366.970 204.290 367.200 205.270 ;
        RECT 367.990 203.340 369.750 212.710 ;
        RECT 433.440 204.430 435.770 204.540 ;
        RECT 444.230 204.430 447.070 213.330 ;
        RECT 350.520 200.820 350.750 201.800 ;
        RECT 353.810 200.820 354.040 201.800 ;
        RECT 357.100 200.820 357.330 201.800 ;
        RECT 360.390 200.820 360.620 201.800 ;
        RECT 363.680 200.820 363.910 201.800 ;
        RECT 366.970 200.820 367.200 201.800 ;
        RECT 367.990 198.170 369.370 203.340 ;
        RECT 433.130 201.980 447.070 204.430 ;
        RECT 383.270 198.170 384.770 198.230 ;
        RECT 367.540 198.110 384.770 198.170 ;
        RECT 310.580 197.270 384.770 198.110 ;
        RECT 310.700 197.090 369.350 197.270 ;
        RECT 329.760 196.850 331.140 197.090 ;
        RECT 383.270 195.410 384.770 197.270 ;
        RECT 392.480 196.930 394.170 197.640 ;
        RECT 425.140 197.010 426.860 197.710 ;
        RECT 270.430 174.010 270.660 175.590 ;
        RECT 275.720 174.010 275.950 175.590 ;
        RECT 281.010 174.010 281.240 175.590 ;
        RECT 286.300 174.010 286.530 175.590 ;
        RECT 291.590 174.010 291.820 175.590 ;
        RECT 296.880 174.010 297.110 175.590 ;
        RECT 298.000 170.780 300.060 180.420 ;
        RECT 383.170 177.650 384.890 195.410 ;
        RECT 385.820 194.550 386.050 195.530 ;
        RECT 389.110 194.550 389.340 195.530 ;
        RECT 392.400 194.550 392.630 195.530 ;
        RECT 395.690 194.550 395.920 195.530 ;
        RECT 398.980 194.550 399.210 195.530 ;
        RECT 385.820 191.080 386.050 192.060 ;
        RECT 389.110 191.080 389.340 192.060 ;
        RECT 392.400 191.080 392.630 192.060 ;
        RECT 395.690 191.080 395.920 192.060 ;
        RECT 398.980 191.080 399.210 192.060 ;
        RECT 385.820 187.610 386.050 188.590 ;
        RECT 389.110 187.610 389.340 188.590 ;
        RECT 392.400 187.610 392.630 188.590 ;
        RECT 395.690 187.610 395.920 188.590 ;
        RECT 398.980 187.610 399.210 188.590 ;
        RECT 385.820 184.140 386.050 185.120 ;
        RECT 389.110 184.140 389.340 185.120 ;
        RECT 392.400 184.140 392.630 185.120 ;
        RECT 395.690 184.140 395.920 185.120 ;
        RECT 398.980 184.140 399.210 185.120 ;
        RECT 385.820 180.670 386.050 181.650 ;
        RECT 389.110 180.670 389.340 181.650 ;
        RECT 392.400 180.670 392.630 181.650 ;
        RECT 395.690 180.670 395.920 181.650 ;
        RECT 398.980 180.670 399.210 181.650 ;
        RECT 383.400 174.370 384.660 177.650 ;
        RECT 385.820 177.200 386.050 178.180 ;
        RECT 389.110 177.200 389.340 178.180 ;
        RECT 392.400 177.200 392.630 178.180 ;
        RECT 395.690 177.200 395.920 178.180 ;
        RECT 398.980 177.200 399.210 178.180 ;
        RECT 399.800 177.620 401.520 195.380 ;
        RECT 405.740 194.520 405.970 195.500 ;
        RECT 412.320 194.520 412.550 195.500 ;
        RECT 405.740 191.050 405.970 192.030 ;
        RECT 412.320 191.050 412.550 192.030 ;
        RECT 405.740 187.580 405.970 188.560 ;
        RECT 412.320 187.580 412.550 188.560 ;
        RECT 405.740 184.110 405.970 185.090 ;
        RECT 412.320 184.110 412.550 185.090 ;
        RECT 405.740 180.640 405.970 181.620 ;
        RECT 412.320 180.640 412.550 181.620 ;
        RECT 405.740 177.770 405.970 178.150 ;
        RECT 400.080 174.370 401.340 177.620 ;
        RECT 405.470 174.370 406.130 177.770 ;
        RECT 412.320 177.170 412.550 178.150 ;
        RECT 416.350 177.620 418.070 195.380 ;
        RECT 419.000 194.520 419.230 195.500 ;
        RECT 422.290 194.520 422.520 195.500 ;
        RECT 425.580 194.520 425.810 195.500 ;
        RECT 428.870 194.520 429.100 195.500 ;
        RECT 432.160 194.520 432.390 195.500 ;
        RECT 433.440 193.810 435.770 201.980 ;
        RECT 444.230 201.880 447.070 201.980 ;
        RECT 419.000 191.050 419.230 192.030 ;
        RECT 422.290 191.050 422.520 192.030 ;
        RECT 425.580 191.050 425.810 192.030 ;
        RECT 428.870 191.050 429.100 192.030 ;
        RECT 432.160 191.050 432.390 192.030 ;
        RECT 419.000 187.580 419.230 188.560 ;
        RECT 422.290 187.580 422.520 188.560 ;
        RECT 425.580 187.580 425.810 188.560 ;
        RECT 428.870 187.580 429.100 188.560 ;
        RECT 432.160 187.580 432.390 188.560 ;
        RECT 419.000 184.110 419.230 185.090 ;
        RECT 422.290 184.110 422.520 185.090 ;
        RECT 425.580 184.110 425.810 185.090 ;
        RECT 428.870 184.110 429.100 185.090 ;
        RECT 432.160 184.110 432.390 185.090 ;
        RECT 419.000 180.640 419.230 181.620 ;
        RECT 422.290 180.640 422.520 181.620 ;
        RECT 425.580 180.640 425.810 181.620 ;
        RECT 428.870 180.640 429.100 181.620 ;
        RECT 432.160 180.640 432.390 181.620 ;
        RECT 416.680 174.370 417.940 177.620 ;
        RECT 419.000 177.170 419.230 178.150 ;
        RECT 422.290 177.170 422.520 178.150 ;
        RECT 425.580 177.170 425.810 178.150 ;
        RECT 428.870 177.170 429.100 178.150 ;
        RECT 432.160 177.170 432.390 178.150 ;
        RECT 433.480 176.210 435.040 193.810 ;
        RECT 433.550 174.370 434.810 176.210 ;
        RECT 383.400 173.350 434.820 174.370 ;
        RECT 416.680 173.140 417.940 173.350 ;
        RECT 270.430 168.540 270.660 170.120 ;
        RECT 275.720 168.540 275.950 170.120 ;
        RECT 281.010 168.540 281.240 170.120 ;
        RECT 286.300 168.540 286.530 170.120 ;
        RECT 291.590 168.540 291.820 170.120 ;
        RECT 296.880 168.540 297.110 170.120 ;
        RECT 270.430 163.070 270.660 164.650 ;
        RECT 275.720 163.070 275.950 164.650 ;
        RECT 281.010 163.070 281.240 164.650 ;
        RECT 286.300 163.070 286.530 164.650 ;
        RECT 291.590 163.070 291.820 164.650 ;
        RECT 296.880 163.070 297.110 164.650 ;
        RECT 270.430 155.780 270.660 157.360 ;
        RECT 275.720 155.780 275.950 157.360 ;
        RECT 281.010 155.780 281.240 157.360 ;
        RECT 286.300 155.780 286.530 157.360 ;
        RECT 291.590 155.780 291.820 157.360 ;
        RECT 296.880 155.780 297.110 157.360 ;
        RECT 270.430 150.310 270.660 151.890 ;
        RECT 275.720 150.310 275.950 151.890 ;
        RECT 281.010 150.310 281.240 151.890 ;
        RECT 286.300 150.310 286.530 151.890 ;
        RECT 291.590 150.310 291.820 151.890 ;
        RECT 296.880 150.310 297.110 151.890 ;
        RECT 298.400 150.450 300.060 170.780 ;
        RECT 270.430 144.840 270.660 146.420 ;
        RECT 275.720 144.840 275.950 146.420 ;
        RECT 281.010 144.840 281.240 146.420 ;
        RECT 286.300 144.840 286.530 146.420 ;
        RECT 291.590 144.840 291.820 146.420 ;
        RECT 296.880 144.840 297.110 146.420 ;
        RECT 270.430 139.370 270.660 140.950 ;
        RECT 275.720 139.370 275.950 140.950 ;
        RECT 281.010 139.370 281.240 140.950 ;
        RECT 286.300 139.370 286.530 140.950 ;
        RECT 291.590 139.370 291.820 140.950 ;
        RECT 296.880 139.370 297.110 140.950 ;
        RECT 297.930 140.670 300.150 150.450 ;
        RECT 270.430 133.900 270.660 135.480 ;
        RECT 275.720 133.900 275.950 135.480 ;
        RECT 281.010 133.900 281.240 135.480 ;
        RECT 286.300 133.900 286.530 135.480 ;
        RECT 291.590 133.900 291.820 135.480 ;
        RECT 296.880 133.900 297.110 135.480 ;
        RECT 270.430 126.600 270.660 128.180 ;
        RECT 275.720 126.600 275.950 128.180 ;
        RECT 281.010 126.600 281.240 128.180 ;
        RECT 286.300 126.600 286.530 128.180 ;
        RECT 291.590 126.600 291.820 128.180 ;
        RECT 296.880 126.600 297.110 128.180 ;
        RECT 270.430 121.130 270.660 122.710 ;
        RECT 275.720 121.130 275.950 122.710 ;
        RECT 281.010 121.130 281.240 122.710 ;
        RECT 286.300 121.130 286.530 122.710 ;
        RECT 291.590 121.130 291.820 122.710 ;
        RECT 296.880 121.130 297.110 122.710 ;
        RECT 298.400 122.570 300.060 140.670 ;
        RECT 337.730 130.800 341.560 131.740 ;
        RECT 469.740 130.670 472.390 131.580 ;
        RECT 310.530 126.320 310.760 127.900 ;
        RECT 315.820 126.320 316.050 127.900 ;
        RECT 321.110 126.320 321.340 127.900 ;
        RECT 326.400 126.320 326.630 127.900 ;
        RECT 331.690 126.320 331.920 127.900 ;
        RECT 336.980 126.320 337.210 127.900 ;
        RECT 270.430 115.660 270.660 117.240 ;
        RECT 275.720 115.660 275.950 117.240 ;
        RECT 281.010 115.660 281.240 117.240 ;
        RECT 286.300 115.660 286.530 117.240 ;
        RECT 291.590 115.660 291.820 117.240 ;
        RECT 296.880 115.660 297.110 117.240 ;
        RECT 297.860 112.090 300.060 122.570 ;
        RECT 310.530 120.850 310.760 122.430 ;
        RECT 315.820 120.850 316.050 122.430 ;
        RECT 321.110 120.850 321.340 122.430 ;
        RECT 326.400 120.850 326.630 122.430 ;
        RECT 331.690 120.850 331.920 122.430 ;
        RECT 336.980 120.850 337.210 122.430 ;
        RECT 307.290 116.400 308.040 120.800 ;
        RECT 338.460 118.950 341.620 126.810 ;
        RECT 342.840 126.310 343.070 127.890 ;
        RECT 348.130 126.310 348.360 127.890 ;
        RECT 353.420 126.310 353.650 127.890 ;
        RECT 358.710 126.310 358.940 127.890 ;
        RECT 364.000 126.310 364.230 127.890 ;
        RECT 369.290 126.310 369.520 127.890 ;
        RECT 381.600 126.180 381.830 127.760 ;
        RECT 392.180 126.180 392.410 127.760 ;
        RECT 402.760 126.180 402.990 127.760 ;
        RECT 413.910 126.170 414.140 127.750 ;
        RECT 424.490 126.170 424.720 127.750 ;
        RECT 435.070 126.170 435.300 127.750 ;
        RECT 442.480 126.140 442.710 127.720 ;
        RECT 447.770 126.140 448.000 127.720 ;
        RECT 453.060 126.140 453.290 127.720 ;
        RECT 458.350 126.140 458.580 127.720 ;
        RECT 463.640 126.140 463.870 127.720 ;
        RECT 468.930 126.140 469.160 127.720 ;
        RECT 474.790 126.130 475.020 127.710 ;
        RECT 480.080 126.130 480.310 127.710 ;
        RECT 485.370 126.130 485.600 127.710 ;
        RECT 490.660 126.130 490.890 127.710 ;
        RECT 495.950 126.130 496.180 127.710 ;
        RECT 501.240 126.130 501.470 127.710 ;
        RECT 438.100 125.520 441.120 125.530 ;
        RECT 342.840 120.840 343.070 122.420 ;
        RECT 348.130 120.840 348.360 122.420 ;
        RECT 353.420 120.840 353.650 122.420 ;
        RECT 358.710 120.840 358.940 122.420 ;
        RECT 364.000 120.840 364.230 122.420 ;
        RECT 369.290 120.840 369.520 122.420 ;
        RECT 310.530 116.400 310.760 116.960 ;
        RECT 307.290 115.770 310.760 116.400 ;
        RECT 307.290 112.570 308.040 115.770 ;
        RECT 310.530 115.380 310.760 115.770 ;
        RECT 315.820 115.380 316.050 116.960 ;
        RECT 321.110 115.380 321.340 116.960 ;
        RECT 326.400 115.380 326.630 116.960 ;
        RECT 331.690 115.380 331.920 116.960 ;
        RECT 336.980 115.380 337.210 116.960 ;
        RECT 270.430 110.190 270.660 111.770 ;
        RECT 275.720 110.190 275.950 111.770 ;
        RECT 281.010 110.190 281.240 111.770 ;
        RECT 286.300 110.190 286.530 111.770 ;
        RECT 291.590 110.190 291.820 111.770 ;
        RECT 296.880 110.190 297.110 111.770 ;
        RECT 270.430 104.720 270.660 106.300 ;
        RECT 275.720 104.720 275.950 106.300 ;
        RECT 281.010 104.720 281.240 106.300 ;
        RECT 286.300 104.720 286.530 106.300 ;
        RECT 291.590 104.720 291.820 106.300 ;
        RECT 296.880 104.720 297.110 106.300 ;
        RECT 270.430 97.280 270.660 98.860 ;
        RECT 275.720 97.280 275.950 98.860 ;
        RECT 281.010 97.280 281.240 98.860 ;
        RECT 286.300 97.280 286.530 98.860 ;
        RECT 291.590 97.280 291.820 98.860 ;
        RECT 296.880 97.280 297.110 98.860 ;
        RECT 298.400 93.430 300.060 112.090 ;
        RECT 310.530 109.910 310.760 111.490 ;
        RECT 315.820 109.910 316.050 111.490 ;
        RECT 321.110 109.910 321.340 111.490 ;
        RECT 326.400 109.910 326.630 111.490 ;
        RECT 331.690 109.910 331.920 111.490 ;
        RECT 336.980 109.910 337.210 111.490 ;
        RECT 310.530 105.060 310.760 106.020 ;
        RECT 310.400 97.800 310.900 105.060 ;
        RECT 315.820 104.440 316.050 106.020 ;
        RECT 321.110 104.440 321.340 106.020 ;
        RECT 326.400 104.440 326.630 106.020 ;
        RECT 331.690 104.440 331.920 106.020 ;
        RECT 336.980 105.220 337.210 106.020 ;
        RECT 310.560 97.130 310.790 97.800 ;
        RECT 315.850 97.130 316.080 98.710 ;
        RECT 321.140 97.130 321.370 98.710 ;
        RECT 326.430 97.130 326.660 98.710 ;
        RECT 331.720 97.130 331.950 98.710 ;
        RECT 336.870 97.960 337.370 105.220 ;
        RECT 337.010 97.130 337.240 97.960 ;
        RECT 270.430 91.810 270.660 93.390 ;
        RECT 275.720 91.810 275.950 93.390 ;
        RECT 281.010 91.810 281.240 93.390 ;
        RECT 286.300 91.810 286.530 93.390 ;
        RECT 291.590 91.810 291.820 93.390 ;
        RECT 296.880 91.810 297.110 93.390 ;
        RECT 270.430 86.340 270.660 87.920 ;
        RECT 275.720 86.340 275.950 87.920 ;
        RECT 281.010 86.340 281.240 87.920 ;
        RECT 286.300 86.340 286.530 87.920 ;
        RECT 291.590 86.340 291.820 87.920 ;
        RECT 296.880 86.340 297.110 87.920 ;
        RECT 298.140 83.510 300.060 93.430 ;
        RECT 310.560 91.660 310.790 93.240 ;
        RECT 315.850 91.660 316.080 93.240 ;
        RECT 321.140 91.660 321.370 93.240 ;
        RECT 326.430 91.660 326.660 93.240 ;
        RECT 331.720 91.660 331.950 93.240 ;
        RECT 337.010 91.660 337.240 93.240 ;
        RECT 270.430 80.870 270.660 82.450 ;
        RECT 275.720 80.870 275.950 82.450 ;
        RECT 281.010 80.870 281.240 82.450 ;
        RECT 286.300 80.870 286.530 82.450 ;
        RECT 291.590 80.870 291.820 82.450 ;
        RECT 296.880 80.870 297.110 82.450 ;
        RECT 270.430 75.400 270.660 76.980 ;
        RECT 275.720 75.400 275.950 76.980 ;
        RECT 281.010 75.400 281.240 76.980 ;
        RECT 286.300 75.400 286.530 76.980 ;
        RECT 291.590 75.400 291.820 76.980 ;
        RECT 296.880 75.400 297.110 76.980 ;
        RECT 270.480 68.000 270.710 69.580 ;
        RECT 275.770 68.000 276.000 69.580 ;
        RECT 281.060 68.000 281.290 69.580 ;
        RECT 286.350 68.000 286.580 69.580 ;
        RECT 291.640 68.000 291.870 69.580 ;
        RECT 296.930 68.000 297.160 69.580 ;
        RECT 270.480 62.530 270.710 64.110 ;
        RECT 275.770 62.530 276.000 64.110 ;
        RECT 281.060 62.530 281.290 64.110 ;
        RECT 286.350 62.530 286.580 64.110 ;
        RECT 291.640 62.530 291.870 64.110 ;
        RECT 296.930 62.530 297.160 64.110 ;
        RECT 298.400 63.470 300.060 83.510 ;
        RECT 307.320 83.380 308.070 91.610 ;
        RECT 310.560 86.190 310.790 87.770 ;
        RECT 315.850 86.190 316.080 87.770 ;
        RECT 321.140 86.190 321.370 87.770 ;
        RECT 326.430 86.190 326.660 87.770 ;
        RECT 331.720 86.190 331.950 87.770 ;
        RECT 337.010 86.190 337.240 87.770 ;
        RECT 310.560 80.720 310.790 82.300 ;
        RECT 315.850 80.720 316.080 82.300 ;
        RECT 321.140 80.720 321.370 82.300 ;
        RECT 326.430 80.720 326.660 82.300 ;
        RECT 331.720 80.720 331.950 82.300 ;
        RECT 337.010 80.720 337.240 82.300 ;
        RECT 310.560 75.730 310.790 76.830 ;
        RECT 310.400 68.470 310.900 75.730 ;
        RECT 315.850 75.250 316.080 76.830 ;
        RECT 321.140 75.250 321.370 76.830 ;
        RECT 326.430 75.250 326.660 76.830 ;
        RECT 331.720 75.250 331.950 76.830 ;
        RECT 337.010 76.060 337.240 76.830 ;
        RECT 310.560 67.840 310.790 68.470 ;
        RECT 315.850 67.840 316.080 69.420 ;
        RECT 321.140 67.840 321.370 69.420 ;
        RECT 326.430 67.840 326.660 69.420 ;
        RECT 331.720 67.840 331.950 69.420 ;
        RECT 336.870 68.800 337.370 76.060 ;
        RECT 337.010 67.840 337.240 68.800 ;
        RECT 270.480 57.060 270.710 58.640 ;
        RECT 275.770 57.060 276.000 58.640 ;
        RECT 281.060 57.060 281.290 58.640 ;
        RECT 286.350 57.060 286.580 58.640 ;
        RECT 291.640 57.060 291.870 58.640 ;
        RECT 296.930 57.060 297.160 58.640 ;
        RECT 298.210 55.010 300.060 63.470 ;
        RECT 310.560 62.370 310.790 63.950 ;
        RECT 315.850 62.370 316.080 63.950 ;
        RECT 321.140 62.370 321.370 63.950 ;
        RECT 326.430 62.370 326.660 63.950 ;
        RECT 331.720 62.370 331.950 63.950 ;
        RECT 337.010 62.370 337.240 63.950 ;
        RECT 270.480 51.590 270.710 53.170 ;
        RECT 275.770 51.590 276.000 53.170 ;
        RECT 281.060 51.590 281.290 53.170 ;
        RECT 286.350 51.590 286.580 53.170 ;
        RECT 291.640 51.590 291.870 53.170 ;
        RECT 296.930 51.590 297.160 53.170 ;
        RECT 270.480 46.120 270.710 47.700 ;
        RECT 275.770 46.120 276.000 47.700 ;
        RECT 281.060 46.120 281.290 47.700 ;
        RECT 286.350 46.120 286.580 47.700 ;
        RECT 291.640 46.120 291.870 47.700 ;
        RECT 296.930 46.120 297.160 47.700 ;
        RECT 270.570 38.460 270.800 40.040 ;
        RECT 275.860 38.460 276.090 40.040 ;
        RECT 281.150 38.460 281.380 40.040 ;
        RECT 286.440 38.460 286.670 40.040 ;
        RECT 291.730 38.460 291.960 40.040 ;
        RECT 297.020 38.460 297.250 40.040 ;
        RECT 270.570 32.990 270.800 34.570 ;
        RECT 275.860 32.990 276.090 34.570 ;
        RECT 281.150 32.990 281.380 34.570 ;
        RECT 286.440 32.990 286.670 34.570 ;
        RECT 291.730 32.990 291.960 34.570 ;
        RECT 297.020 32.990 297.250 34.570 ;
        RECT 298.400 34.060 300.060 55.010 ;
        RECT 307.320 54.090 308.070 62.320 ;
        RECT 310.560 56.900 310.790 58.480 ;
        RECT 315.850 56.900 316.080 58.480 ;
        RECT 321.140 56.900 321.370 58.480 ;
        RECT 326.430 56.900 326.660 58.480 ;
        RECT 331.720 56.900 331.950 58.480 ;
        RECT 337.010 56.900 337.240 58.480 ;
        RECT 310.560 51.430 310.790 53.010 ;
        RECT 315.850 51.430 316.080 53.010 ;
        RECT 321.140 51.430 321.370 53.010 ;
        RECT 326.430 51.430 326.660 53.010 ;
        RECT 331.720 51.430 331.950 53.010 ;
        RECT 337.010 51.430 337.240 53.010 ;
        RECT 310.560 46.460 310.790 47.540 ;
        RECT 310.460 39.200 310.960 46.460 ;
        RECT 315.850 45.960 316.080 47.540 ;
        RECT 321.140 45.960 321.370 47.540 ;
        RECT 326.430 45.960 326.660 47.540 ;
        RECT 331.720 45.960 331.950 47.540 ;
        RECT 337.010 46.630 337.240 47.540 ;
        RECT 310.560 38.550 310.790 39.200 ;
        RECT 315.850 38.550 316.080 40.130 ;
        RECT 321.140 38.550 321.370 40.130 ;
        RECT 326.430 38.550 326.660 40.130 ;
        RECT 331.720 38.550 331.950 40.130 ;
        RECT 336.810 39.370 337.310 46.630 ;
        RECT 337.010 38.550 337.240 39.370 ;
        RECT 270.570 28.600 270.800 29.100 ;
        RECT 265.680 27.570 270.980 28.600 ;
        RECT 232.980 27.030 236.460 27.390 ;
        RECT 234.180 26.720 235.850 27.030 ;
        RECT 265.680 26.880 269.160 27.570 ;
        RECT 270.570 27.520 270.800 27.570 ;
        RECT 275.860 27.520 276.090 29.100 ;
        RECT 281.150 27.520 281.380 29.100 ;
        RECT 286.440 27.520 286.670 29.100 ;
        RECT 291.730 27.520 291.960 29.100 ;
        RECT 297.020 28.510 297.250 29.100 ;
        RECT 298.000 28.510 300.060 34.060 ;
        RECT 310.560 33.080 310.790 34.660 ;
        RECT 315.850 33.080 316.080 34.660 ;
        RECT 321.140 33.080 321.370 34.660 ;
        RECT 326.430 33.080 326.660 34.660 ;
        RECT 331.720 33.080 331.950 34.660 ;
        RECT 337.010 33.080 337.240 34.660 ;
        RECT 296.820 27.390 300.060 28.510 ;
        RECT 234.760 24.640 235.510 26.720 ;
        RECT 267.330 24.710 268.080 26.880 ;
        RECT 298.000 25.870 300.060 27.390 ;
        RECT 205.060 21.870 205.290 23.450 ;
        RECT 210.350 21.870 210.580 23.450 ;
        RECT 215.640 21.870 215.870 23.450 ;
        RECT 220.930 21.870 221.160 23.450 ;
        RECT 226.220 21.870 226.450 23.450 ;
        RECT 231.510 21.870 231.740 23.450 ;
        RECT 238.000 21.980 238.230 23.560 ;
        RECT 243.290 21.980 243.520 23.560 ;
        RECT 248.580 21.980 248.810 23.560 ;
        RECT 253.870 21.980 254.100 23.560 ;
        RECT 259.160 21.980 259.390 23.560 ;
        RECT 264.450 21.980 264.680 23.560 ;
        RECT 270.570 22.050 270.800 23.630 ;
        RECT 275.860 22.050 276.090 23.630 ;
        RECT 281.150 22.050 281.380 23.630 ;
        RECT 286.440 22.050 286.670 23.630 ;
        RECT 291.730 22.050 291.960 23.630 ;
        RECT 297.020 22.050 297.250 23.630 ;
        RECT 136.390 -15.670 137.870 17.650 ;
        RECT 169.240 -15.670 170.720 18.940 ;
        RECT 205.060 16.400 205.290 17.980 ;
        RECT 210.350 16.400 210.580 17.980 ;
        RECT 215.640 16.400 215.870 17.980 ;
        RECT 220.930 16.400 221.160 17.980 ;
        RECT 226.220 16.400 226.450 17.980 ;
        RECT 231.510 16.400 231.740 17.980 ;
        RECT 238.000 16.510 238.230 18.090 ;
        RECT 243.290 16.510 243.520 18.090 ;
        RECT 248.580 16.510 248.810 18.090 ;
        RECT 253.870 16.510 254.100 18.090 ;
        RECT 259.160 16.510 259.390 18.090 ;
        RECT 264.450 16.510 264.680 18.090 ;
        RECT 270.570 16.580 270.800 18.160 ;
        RECT 275.860 16.580 276.090 18.160 ;
        RECT 281.150 16.580 281.380 18.160 ;
        RECT 286.440 16.580 286.670 18.160 ;
        RECT 291.730 16.580 291.960 18.160 ;
        RECT 297.020 16.580 297.250 18.160 ;
        RECT 298.400 17.870 300.060 25.870 ;
        RECT 307.320 24.800 308.070 33.030 ;
        RECT 310.560 27.610 310.790 29.190 ;
        RECT 315.850 27.610 316.080 29.190 ;
        RECT 321.140 27.610 321.370 29.190 ;
        RECT 326.430 27.610 326.660 29.190 ;
        RECT 331.720 27.610 331.950 29.190 ;
        RECT 337.010 27.610 337.240 29.190 ;
        RECT 337.980 27.960 341.620 118.950 ;
        RECT 342.840 115.370 343.070 116.950 ;
        RECT 348.130 115.370 348.360 116.950 ;
        RECT 353.420 115.370 353.650 116.950 ;
        RECT 358.710 115.370 358.940 116.950 ;
        RECT 364.000 115.370 364.230 116.950 ;
        RECT 369.290 115.370 369.520 116.950 ;
        RECT 342.840 109.900 343.070 111.480 ;
        RECT 348.130 109.900 348.360 111.480 ;
        RECT 353.420 109.900 353.650 111.480 ;
        RECT 358.710 109.900 358.940 111.480 ;
        RECT 364.000 109.900 364.230 111.480 ;
        RECT 369.290 109.900 369.520 111.480 ;
        RECT 342.840 105.330 343.070 106.010 ;
        RECT 342.810 98.070 343.310 105.330 ;
        RECT 348.130 104.430 348.360 106.010 ;
        RECT 353.420 104.430 353.650 106.010 ;
        RECT 358.710 104.430 358.940 106.010 ;
        RECT 364.000 104.430 364.230 106.010 ;
        RECT 369.290 105.660 369.520 106.010 ;
        RECT 342.880 97.190 343.110 98.070 ;
        RECT 348.170 97.190 348.400 98.770 ;
        RECT 353.460 97.190 353.690 98.770 ;
        RECT 358.750 97.190 358.980 98.770 ;
        RECT 364.040 97.190 364.270 98.770 ;
        RECT 369.110 98.180 369.770 105.660 ;
        RECT 369.330 97.190 369.560 98.180 ;
        RECT 342.880 91.720 343.110 93.300 ;
        RECT 348.170 91.720 348.400 93.300 ;
        RECT 353.460 91.720 353.690 93.300 ;
        RECT 358.750 91.720 358.980 93.300 ;
        RECT 364.040 91.720 364.270 93.300 ;
        RECT 369.330 91.720 369.560 93.300 ;
        RECT 342.880 86.250 343.110 87.830 ;
        RECT 348.170 86.250 348.400 87.830 ;
        RECT 353.460 86.250 353.690 87.830 ;
        RECT 358.750 86.250 358.980 87.830 ;
        RECT 364.040 86.250 364.270 87.830 ;
        RECT 369.330 86.250 369.560 87.830 ;
        RECT 342.880 80.780 343.110 82.360 ;
        RECT 348.170 80.780 348.400 82.360 ;
        RECT 353.460 80.780 353.690 82.360 ;
        RECT 358.750 80.780 358.980 82.360 ;
        RECT 364.040 80.780 364.270 82.360 ;
        RECT 369.330 80.780 369.560 82.360 ;
        RECT 342.880 75.900 343.110 76.890 ;
        RECT 342.590 75.310 343.110 75.900 ;
        RECT 348.170 75.310 348.400 76.890 ;
        RECT 353.460 75.310 353.690 76.890 ;
        RECT 358.750 75.310 358.980 76.890 ;
        RECT 364.040 75.310 364.270 76.890 ;
        RECT 369.330 75.900 369.560 76.890 ;
        RECT 342.590 69.410 343.090 75.310 ;
        RECT 342.590 68.640 343.130 69.410 ;
        RECT 342.900 67.830 343.130 68.640 ;
        RECT 348.190 67.830 348.420 69.410 ;
        RECT 353.480 67.830 353.710 69.410 ;
        RECT 358.770 67.830 359.000 69.410 ;
        RECT 364.060 67.830 364.290 69.410 ;
        RECT 369.000 68.420 369.660 75.900 ;
        RECT 369.350 67.830 369.580 68.420 ;
        RECT 342.900 62.360 343.130 63.940 ;
        RECT 348.190 62.360 348.420 63.940 ;
        RECT 353.480 62.360 353.710 63.940 ;
        RECT 358.770 62.360 359.000 63.940 ;
        RECT 364.060 62.360 364.290 63.940 ;
        RECT 369.350 62.360 369.580 63.940 ;
        RECT 342.900 56.890 343.130 58.470 ;
        RECT 348.190 56.890 348.420 58.470 ;
        RECT 353.480 56.890 353.710 58.470 ;
        RECT 358.770 56.890 359.000 58.470 ;
        RECT 364.060 56.890 364.290 58.470 ;
        RECT 369.350 56.890 369.580 58.470 ;
        RECT 342.900 51.420 343.130 53.000 ;
        RECT 348.190 51.420 348.420 53.000 ;
        RECT 353.480 51.420 353.710 53.000 ;
        RECT 358.770 51.420 359.000 53.000 ;
        RECT 364.060 51.420 364.290 53.000 ;
        RECT 369.350 51.420 369.580 53.000 ;
        RECT 342.900 46.740 343.130 47.530 ;
        RECT 342.750 39.480 343.250 46.740 ;
        RECT 348.190 45.950 348.420 47.530 ;
        RECT 353.480 45.950 353.710 47.530 ;
        RECT 358.770 45.950 359.000 47.530 ;
        RECT 364.060 45.950 364.290 47.530 ;
        RECT 369.350 47.120 369.580 47.530 ;
        RECT 342.920 38.540 343.150 39.480 ;
        RECT 348.210 38.540 348.440 40.120 ;
        RECT 353.500 38.540 353.730 40.120 ;
        RECT 358.790 38.540 359.020 40.120 ;
        RECT 364.080 38.540 364.310 40.120 ;
        RECT 369.160 39.640 369.820 47.120 ;
        RECT 369.370 38.540 369.600 39.640 ;
        RECT 342.920 33.070 343.150 34.650 ;
        RECT 348.210 33.070 348.440 34.650 ;
        RECT 353.500 33.070 353.730 34.650 ;
        RECT 358.790 33.070 359.020 34.650 ;
        RECT 364.080 33.070 364.310 34.650 ;
        RECT 369.370 33.070 369.600 34.650 ;
        RECT 338.460 23.960 341.620 27.960 ;
        RECT 342.920 27.600 343.150 29.180 ;
        RECT 348.210 27.600 348.440 29.180 ;
        RECT 353.500 27.600 353.730 29.180 ;
        RECT 358.790 27.600 359.020 29.180 ;
        RECT 364.080 27.600 364.310 29.180 ;
        RECT 369.370 27.600 369.600 29.180 ;
        RECT 310.560 22.140 310.790 23.720 ;
        RECT 315.850 22.140 316.080 23.720 ;
        RECT 321.140 22.140 321.370 23.720 ;
        RECT 326.430 22.140 326.660 23.720 ;
        RECT 331.720 22.140 331.950 23.720 ;
        RECT 337.010 22.140 337.240 23.720 ;
        RECT 342.920 22.130 343.150 23.710 ;
        RECT 348.210 22.130 348.440 23.710 ;
        RECT 353.500 22.130 353.730 23.710 ;
        RECT 358.790 22.130 359.020 23.710 ;
        RECT 364.080 22.130 364.310 23.710 ;
        RECT 369.370 22.130 369.600 23.710 ;
        RECT 310.560 16.670 310.790 18.250 ;
        RECT 315.850 16.670 316.080 18.250 ;
        RECT 321.140 16.670 321.370 18.250 ;
        RECT 326.430 16.670 326.660 18.250 ;
        RECT 331.720 16.670 331.950 18.250 ;
        RECT 337.010 16.670 337.240 18.250 ;
        RECT 342.920 16.660 343.150 18.240 ;
        RECT 348.210 16.660 348.440 18.240 ;
        RECT 353.500 16.660 353.730 18.240 ;
        RECT 358.790 16.660 359.020 18.240 ;
        RECT 364.080 16.660 364.310 18.240 ;
        RECT 369.370 16.660 369.600 18.240 ;
        RECT 371.400 17.060 375.330 124.410 ;
        RECT 381.600 120.710 381.830 122.290 ;
        RECT 392.180 120.710 392.410 122.290 ;
        RECT 402.760 120.710 402.990 122.290 ;
        RECT 381.600 115.240 381.830 116.820 ;
        RECT 392.180 115.240 392.410 116.820 ;
        RECT 402.760 115.240 402.990 116.820 ;
        RECT 381.600 109.770 381.830 111.350 ;
        RECT 392.180 109.770 392.410 111.350 ;
        RECT 402.760 109.770 402.990 111.350 ;
        RECT 381.600 104.300 381.830 105.880 ;
        RECT 392.180 104.300 392.410 105.880 ;
        RECT 402.760 105.080 402.990 105.880 ;
        RECT 381.630 96.990 381.860 98.570 ;
        RECT 392.210 96.990 392.440 98.570 ;
        RECT 402.650 97.820 403.150 105.080 ;
        RECT 403.590 103.850 407.520 124.750 ;
        RECT 413.910 120.700 414.140 122.280 ;
        RECT 424.490 120.700 424.720 122.280 ;
        RECT 435.070 120.700 435.300 122.280 ;
        RECT 413.910 115.230 414.140 116.810 ;
        RECT 424.490 115.230 424.720 116.810 ;
        RECT 435.070 115.230 435.300 116.810 ;
        RECT 413.910 109.760 414.140 111.340 ;
        RECT 424.490 109.760 424.720 111.340 ;
        RECT 435.070 109.760 435.300 111.340 ;
        RECT 413.910 104.290 414.140 105.870 ;
        RECT 424.490 104.290 424.720 105.870 ;
        RECT 435.070 105.520 435.300 105.870 ;
        RECT 403.600 103.180 407.520 103.850 ;
        RECT 402.790 96.990 403.020 97.820 ;
        RECT 381.630 91.520 381.860 93.100 ;
        RECT 392.210 91.520 392.440 93.100 ;
        RECT 402.790 91.520 403.020 93.100 ;
        RECT 381.630 86.050 381.860 87.630 ;
        RECT 392.210 86.050 392.440 87.630 ;
        RECT 402.790 86.050 403.020 87.630 ;
        RECT 381.630 80.580 381.860 82.160 ;
        RECT 392.210 80.580 392.440 82.160 ;
        RECT 402.790 80.580 403.020 82.160 ;
        RECT 381.630 75.110 381.860 76.690 ;
        RECT 392.210 75.110 392.440 76.690 ;
        RECT 402.790 75.920 403.020 76.690 ;
        RECT 381.630 67.700 381.860 69.280 ;
        RECT 392.210 67.700 392.440 69.280 ;
        RECT 402.650 68.660 403.150 75.920 ;
        RECT 402.790 67.700 403.020 68.660 ;
        RECT 381.630 62.230 381.860 63.810 ;
        RECT 392.210 62.230 392.440 63.810 ;
        RECT 402.790 62.230 403.020 63.810 ;
        RECT 381.630 56.760 381.860 58.340 ;
        RECT 392.210 56.760 392.440 58.340 ;
        RECT 402.790 56.760 403.020 58.340 ;
        RECT 381.630 51.290 381.860 52.870 ;
        RECT 392.210 51.290 392.440 52.870 ;
        RECT 402.790 51.290 403.020 52.870 ;
        RECT 381.630 45.820 381.860 47.400 ;
        RECT 392.210 45.820 392.440 47.400 ;
        RECT 402.790 46.490 403.020 47.400 ;
        RECT 381.630 38.410 381.860 39.990 ;
        RECT 392.210 38.410 392.440 39.990 ;
        RECT 402.590 39.230 403.090 46.490 ;
        RECT 403.590 45.440 407.520 103.180 ;
        RECT 413.950 97.050 414.180 98.630 ;
        RECT 424.530 97.050 424.760 98.630 ;
        RECT 434.890 98.040 435.550 105.520 ;
        RECT 435.110 97.050 435.340 98.040 ;
        RECT 413.950 91.580 414.180 93.160 ;
        RECT 424.530 91.580 424.760 93.160 ;
        RECT 435.110 91.580 435.340 93.160 ;
        RECT 413.950 86.110 414.180 87.690 ;
        RECT 424.530 86.110 424.760 87.690 ;
        RECT 435.110 86.110 435.340 87.690 ;
        RECT 413.950 80.640 414.180 82.220 ;
        RECT 424.530 80.640 424.760 82.220 ;
        RECT 435.110 80.640 435.340 82.220 ;
        RECT 413.950 75.170 414.180 76.750 ;
        RECT 424.530 75.170 424.760 76.750 ;
        RECT 435.110 75.760 435.340 76.750 ;
        RECT 413.970 67.690 414.200 69.270 ;
        RECT 424.550 67.690 424.780 69.270 ;
        RECT 434.780 68.280 435.440 75.760 ;
        RECT 435.130 67.690 435.360 68.280 ;
        RECT 413.970 62.220 414.200 63.800 ;
        RECT 424.550 62.220 424.780 63.800 ;
        RECT 435.130 62.220 435.360 63.800 ;
        RECT 413.970 56.750 414.200 58.330 ;
        RECT 424.550 56.750 424.780 58.330 ;
        RECT 435.130 56.750 435.360 58.330 ;
        RECT 413.970 51.280 414.200 52.860 ;
        RECT 424.550 51.280 424.780 52.860 ;
        RECT 435.130 51.280 435.360 52.860 ;
        RECT 413.970 45.810 414.200 47.390 ;
        RECT 424.550 45.810 424.780 47.390 ;
        RECT 435.130 46.980 435.360 47.390 ;
        RECT 403.600 44.770 407.520 45.440 ;
        RECT 402.790 38.410 403.020 39.230 ;
        RECT 381.630 32.940 381.860 34.520 ;
        RECT 392.210 32.940 392.440 34.520 ;
        RECT 402.790 32.940 403.020 34.520 ;
        RECT 381.630 27.470 381.860 29.050 ;
        RECT 392.210 27.470 392.440 29.050 ;
        RECT 402.790 27.470 403.020 29.050 ;
        RECT 381.630 22.000 381.860 23.580 ;
        RECT 392.210 22.000 392.440 23.580 ;
        RECT 402.790 22.000 403.020 23.580 ;
        RECT 381.630 16.530 381.860 18.110 ;
        RECT 392.210 16.530 392.440 18.110 ;
        RECT 402.790 16.530 403.020 18.110 ;
        RECT 403.590 17.400 407.520 44.770 ;
        RECT 413.990 38.400 414.220 39.980 ;
        RECT 424.570 38.400 424.800 39.980 ;
        RECT 434.940 39.500 435.600 46.980 ;
        RECT 435.150 38.400 435.380 39.500 ;
        RECT 413.990 32.930 414.220 34.510 ;
        RECT 424.570 32.930 424.800 34.510 ;
        RECT 435.150 32.930 435.380 34.510 ;
        RECT 413.990 27.460 414.220 29.040 ;
        RECT 424.570 27.460 424.800 29.040 ;
        RECT 435.150 27.460 435.380 29.040 ;
        RECT 413.990 21.990 414.220 23.570 ;
        RECT 424.570 21.990 424.800 23.570 ;
        RECT 435.150 21.990 435.380 23.570 ;
        RECT 436.820 18.310 441.120 125.520 ;
        RECT 442.480 120.670 442.710 122.250 ;
        RECT 447.770 120.670 448.000 122.250 ;
        RECT 453.060 120.670 453.290 122.250 ;
        RECT 458.350 120.670 458.580 122.250 ;
        RECT 463.640 120.670 463.870 122.250 ;
        RECT 468.930 120.670 469.160 122.250 ;
        RECT 442.480 115.200 442.710 116.780 ;
        RECT 447.770 115.200 448.000 116.780 ;
        RECT 453.060 115.200 453.290 116.780 ;
        RECT 458.350 115.200 458.580 116.780 ;
        RECT 463.640 115.200 463.870 116.780 ;
        RECT 468.930 115.200 469.160 116.780 ;
        RECT 442.480 109.730 442.710 111.310 ;
        RECT 447.770 109.730 448.000 111.310 ;
        RECT 453.060 109.730 453.290 111.310 ;
        RECT 458.350 109.730 458.580 111.310 ;
        RECT 463.640 109.730 463.870 111.310 ;
        RECT 468.930 109.730 469.160 111.310 ;
        RECT 442.480 104.880 442.710 105.840 ;
        RECT 442.350 97.620 442.850 104.880 ;
        RECT 447.770 104.260 448.000 105.840 ;
        RECT 453.060 104.260 453.290 105.840 ;
        RECT 458.350 104.260 458.580 105.840 ;
        RECT 463.640 104.260 463.870 105.840 ;
        RECT 468.930 105.040 469.160 105.840 ;
        RECT 442.510 96.950 442.740 97.620 ;
        RECT 447.800 96.950 448.030 98.530 ;
        RECT 453.090 96.950 453.320 98.530 ;
        RECT 458.380 96.950 458.610 98.530 ;
        RECT 463.670 96.950 463.900 98.530 ;
        RECT 468.820 97.780 469.320 105.040 ;
        RECT 468.960 96.950 469.190 97.780 ;
        RECT 442.510 91.480 442.740 93.060 ;
        RECT 447.800 91.480 448.030 93.060 ;
        RECT 453.090 91.480 453.320 93.060 ;
        RECT 458.380 91.480 458.610 93.060 ;
        RECT 463.670 91.480 463.900 93.060 ;
        RECT 468.960 91.480 469.190 93.060 ;
        RECT 442.510 86.010 442.740 87.590 ;
        RECT 447.800 86.010 448.030 87.590 ;
        RECT 453.090 86.010 453.320 87.590 ;
        RECT 458.380 86.010 458.610 87.590 ;
        RECT 463.670 86.010 463.900 87.590 ;
        RECT 468.960 86.010 469.190 87.590 ;
        RECT 442.510 80.540 442.740 82.120 ;
        RECT 447.800 80.540 448.030 82.120 ;
        RECT 453.090 80.540 453.320 82.120 ;
        RECT 458.380 80.540 458.610 82.120 ;
        RECT 463.670 80.540 463.900 82.120 ;
        RECT 468.960 80.540 469.190 82.120 ;
        RECT 442.510 75.550 442.740 76.650 ;
        RECT 442.350 68.290 442.850 75.550 ;
        RECT 447.800 75.070 448.030 76.650 ;
        RECT 453.090 75.070 453.320 76.650 ;
        RECT 458.380 75.070 458.610 76.650 ;
        RECT 463.670 75.070 463.900 76.650 ;
        RECT 468.960 75.880 469.190 76.650 ;
        RECT 442.510 67.660 442.740 68.290 ;
        RECT 447.800 67.660 448.030 69.240 ;
        RECT 453.090 67.660 453.320 69.240 ;
        RECT 458.380 67.660 458.610 69.240 ;
        RECT 463.670 67.660 463.900 69.240 ;
        RECT 468.820 68.620 469.320 75.880 ;
        RECT 468.960 67.660 469.190 68.620 ;
        RECT 442.510 62.190 442.740 63.770 ;
        RECT 447.800 62.190 448.030 63.770 ;
        RECT 453.090 62.190 453.320 63.770 ;
        RECT 458.380 62.190 458.610 63.770 ;
        RECT 463.670 62.190 463.900 63.770 ;
        RECT 468.960 62.190 469.190 63.770 ;
        RECT 442.510 56.720 442.740 58.300 ;
        RECT 447.800 56.720 448.030 58.300 ;
        RECT 453.090 56.720 453.320 58.300 ;
        RECT 458.380 56.720 458.610 58.300 ;
        RECT 463.670 56.720 463.900 58.300 ;
        RECT 468.960 56.720 469.190 58.300 ;
        RECT 442.510 51.250 442.740 52.830 ;
        RECT 447.800 51.250 448.030 52.830 ;
        RECT 453.090 51.250 453.320 52.830 ;
        RECT 458.380 51.250 458.610 52.830 ;
        RECT 463.670 51.250 463.900 52.830 ;
        RECT 468.960 51.250 469.190 52.830 ;
        RECT 442.510 46.280 442.740 47.360 ;
        RECT 442.410 39.020 442.910 46.280 ;
        RECT 447.800 45.780 448.030 47.360 ;
        RECT 453.090 45.780 453.320 47.360 ;
        RECT 458.380 45.780 458.610 47.360 ;
        RECT 463.670 45.780 463.900 47.360 ;
        RECT 468.960 46.450 469.190 47.360 ;
        RECT 442.510 38.370 442.740 39.020 ;
        RECT 447.800 38.370 448.030 39.950 ;
        RECT 453.090 38.370 453.320 39.950 ;
        RECT 458.380 38.370 458.610 39.950 ;
        RECT 463.670 38.370 463.900 39.950 ;
        RECT 468.760 39.190 469.260 46.450 ;
        RECT 468.960 38.370 469.190 39.190 ;
        RECT 442.510 32.900 442.740 34.480 ;
        RECT 447.800 32.900 448.030 34.480 ;
        RECT 453.090 32.900 453.320 34.480 ;
        RECT 458.380 32.900 458.610 34.480 ;
        RECT 463.670 32.900 463.900 34.480 ;
        RECT 468.960 32.900 469.190 34.480 ;
        RECT 442.510 27.430 442.740 29.010 ;
        RECT 447.800 27.430 448.030 29.010 ;
        RECT 453.090 27.430 453.320 29.010 ;
        RECT 458.380 27.430 458.610 29.010 ;
        RECT 463.670 27.430 463.900 29.010 ;
        RECT 468.960 27.430 469.190 29.010 ;
        RECT 442.510 21.960 442.740 23.540 ;
        RECT 447.800 21.960 448.030 23.540 ;
        RECT 453.090 21.960 453.320 23.540 ;
        RECT 458.380 21.960 458.610 23.540 ;
        RECT 463.670 21.960 463.900 23.540 ;
        RECT 468.960 21.960 469.190 23.540 ;
        RECT 470.380 21.210 473.400 125.010 ;
        RECT 474.790 120.660 475.020 122.240 ;
        RECT 480.080 120.660 480.310 122.240 ;
        RECT 485.370 120.660 485.600 122.240 ;
        RECT 490.660 120.660 490.890 122.240 ;
        RECT 495.950 120.660 496.180 122.240 ;
        RECT 501.240 121.750 501.470 122.240 ;
        RECT 503.380 121.750 506.600 127.830 ;
        RECT 501.160 121.120 506.600 121.750 ;
        RECT 501.240 120.660 501.470 121.120 ;
        RECT 474.790 115.190 475.020 116.770 ;
        RECT 480.080 115.190 480.310 116.770 ;
        RECT 485.370 115.190 485.600 116.770 ;
        RECT 490.660 115.190 490.890 116.770 ;
        RECT 495.950 115.190 496.180 116.770 ;
        RECT 501.240 115.190 501.470 116.770 ;
        RECT 503.380 113.430 506.600 121.120 ;
        RECT 474.790 109.720 475.020 111.300 ;
        RECT 480.080 109.720 480.310 111.300 ;
        RECT 485.370 109.720 485.600 111.300 ;
        RECT 490.660 109.720 490.890 111.300 ;
        RECT 495.950 109.720 496.180 111.300 ;
        RECT 501.240 109.720 501.470 111.300 ;
        RECT 474.790 105.150 475.020 105.830 ;
        RECT 474.760 97.890 475.260 105.150 ;
        RECT 480.080 104.250 480.310 105.830 ;
        RECT 485.370 104.250 485.600 105.830 ;
        RECT 490.660 104.250 490.890 105.830 ;
        RECT 495.950 104.250 496.180 105.830 ;
        RECT 501.240 105.480 501.470 105.830 ;
        RECT 474.830 97.010 475.060 97.890 ;
        RECT 480.120 97.010 480.350 98.590 ;
        RECT 485.410 97.010 485.640 98.590 ;
        RECT 490.700 97.010 490.930 98.590 ;
        RECT 495.990 97.010 496.220 98.590 ;
        RECT 501.060 98.000 501.720 105.480 ;
        RECT 503.380 105.230 506.880 113.430 ;
        RECT 501.280 97.010 501.510 98.000 ;
        RECT 503.940 96.330 506.880 105.230 ;
        RECT 474.830 91.540 475.060 93.120 ;
        RECT 480.120 91.540 480.350 93.120 ;
        RECT 485.410 91.540 485.640 93.120 ;
        RECT 490.700 91.540 490.930 93.120 ;
        RECT 495.990 91.540 496.220 93.120 ;
        RECT 501.280 91.540 501.510 93.120 ;
        RECT 474.830 86.070 475.060 87.650 ;
        RECT 480.120 86.070 480.350 87.650 ;
        RECT 485.410 86.070 485.640 87.650 ;
        RECT 490.700 86.070 490.930 87.650 ;
        RECT 495.990 86.070 496.220 87.650 ;
        RECT 501.280 86.070 501.510 87.650 ;
        RECT 474.830 80.600 475.060 82.180 ;
        RECT 480.120 80.600 480.350 82.180 ;
        RECT 485.410 80.600 485.640 82.180 ;
        RECT 490.700 80.600 490.930 82.180 ;
        RECT 495.990 80.600 496.220 82.180 ;
        RECT 501.280 80.600 501.510 82.180 ;
        RECT 474.830 75.720 475.060 76.710 ;
        RECT 474.540 75.130 475.060 75.720 ;
        RECT 480.120 75.130 480.350 76.710 ;
        RECT 485.410 75.130 485.640 76.710 ;
        RECT 490.700 75.130 490.930 76.710 ;
        RECT 495.990 75.130 496.220 76.710 ;
        RECT 501.280 75.720 501.510 76.710 ;
        RECT 474.540 69.230 475.040 75.130 ;
        RECT 474.540 68.460 475.080 69.230 ;
        RECT 474.850 67.650 475.080 68.460 ;
        RECT 480.140 67.650 480.370 69.230 ;
        RECT 485.430 67.650 485.660 69.230 ;
        RECT 490.720 67.650 490.950 69.230 ;
        RECT 496.010 67.650 496.240 69.230 ;
        RECT 500.950 68.240 501.610 75.720 ;
        RECT 503.150 74.400 506.880 96.330 ;
        RECT 503.940 69.510 506.880 74.400 ;
        RECT 501.300 67.650 501.530 68.240 ;
        RECT 474.850 62.180 475.080 63.760 ;
        RECT 480.140 62.180 480.370 63.760 ;
        RECT 485.430 62.180 485.660 63.760 ;
        RECT 490.720 62.180 490.950 63.760 ;
        RECT 496.010 62.180 496.240 63.760 ;
        RECT 501.300 62.180 501.530 63.760 ;
        RECT 474.850 56.710 475.080 58.290 ;
        RECT 480.140 56.710 480.370 58.290 ;
        RECT 485.430 56.710 485.660 58.290 ;
        RECT 490.720 56.710 490.950 58.290 ;
        RECT 496.010 56.710 496.240 58.290 ;
        RECT 501.300 56.710 501.530 58.290 ;
        RECT 474.850 51.240 475.080 52.820 ;
        RECT 480.140 51.240 480.370 52.820 ;
        RECT 485.430 51.240 485.660 52.820 ;
        RECT 490.720 51.240 490.950 52.820 ;
        RECT 496.010 51.240 496.240 52.820 ;
        RECT 501.300 51.240 501.530 52.820 ;
        RECT 474.850 46.560 475.080 47.350 ;
        RECT 474.700 39.300 475.200 46.560 ;
        RECT 480.140 45.770 480.370 47.350 ;
        RECT 485.430 45.770 485.660 47.350 ;
        RECT 490.720 45.770 490.950 47.350 ;
        RECT 496.010 45.770 496.240 47.350 ;
        RECT 501.300 46.940 501.530 47.350 ;
        RECT 474.870 38.360 475.100 39.300 ;
        RECT 480.160 38.360 480.390 39.940 ;
        RECT 485.450 38.360 485.680 39.940 ;
        RECT 490.740 38.360 490.970 39.940 ;
        RECT 496.030 38.360 496.260 39.940 ;
        RECT 501.110 39.460 501.770 46.940 ;
        RECT 503.150 46.470 506.880 69.510 ;
        RECT 501.320 38.360 501.550 39.460 ;
        RECT 503.940 38.560 506.880 46.470 ;
        RECT 474.870 32.890 475.100 34.470 ;
        RECT 480.160 32.890 480.390 34.470 ;
        RECT 485.450 32.890 485.680 34.470 ;
        RECT 490.740 32.890 490.970 34.470 ;
        RECT 496.030 32.890 496.260 34.470 ;
        RECT 501.320 32.890 501.550 34.470 ;
        RECT 474.870 27.420 475.100 29.000 ;
        RECT 480.160 27.420 480.390 29.000 ;
        RECT 485.450 27.420 485.680 29.000 ;
        RECT 490.740 27.420 490.970 29.000 ;
        RECT 496.030 27.420 496.260 29.000 ;
        RECT 501.320 27.420 501.550 29.000 ;
        RECT 474.870 21.950 475.100 23.530 ;
        RECT 480.160 21.950 480.390 23.530 ;
        RECT 485.450 21.950 485.680 23.530 ;
        RECT 490.740 21.950 490.970 23.530 ;
        RECT 496.030 21.950 496.260 23.530 ;
        RECT 501.320 21.950 501.550 23.530 ;
        RECT 435.180 18.100 441.120 18.310 ;
        RECT 199.120 -6.260 207.850 -2.450 ;
        RECT 297.540 -3.440 303.030 -0.890 ;
        RECT 335.340 -0.990 346.330 4.230 ;
        RECT 201.420 -15.670 203.290 -6.260 ;
        RECT 299.050 -15.670 300.710 -3.440 ;
        RECT 338.160 -15.670 342.400 -0.990 ;
        RECT 368.310 -1.170 379.300 4.050 ;
        RECT 370.770 -15.670 376.290 -1.170 ;
        RECT 404.100 -15.670 406.860 17.400 ;
        RECT 413.990 16.520 414.220 18.100 ;
        RECT 424.570 16.520 424.800 18.100 ;
        RECT 435.150 17.950 441.120 18.100 ;
        RECT 435.030 16.700 441.120 17.950 ;
        RECT 435.150 16.560 441.120 16.700 ;
        RECT 435.150 16.520 435.380 16.560 ;
        RECT 438.380 16.280 441.120 16.560 ;
        RECT 442.510 16.490 442.740 18.070 ;
        RECT 447.800 16.490 448.030 18.070 ;
        RECT 453.090 16.490 453.320 18.070 ;
        RECT 458.380 16.490 458.610 18.070 ;
        RECT 463.670 16.490 463.900 18.070 ;
        RECT 468.960 16.490 469.190 18.070 ;
        RECT 438.360 -15.670 441.120 16.280 ;
        RECT 470.600 -15.670 473.360 21.210 ;
        RECT 474.870 16.480 475.100 18.060 ;
        RECT 480.160 16.480 480.390 18.060 ;
        RECT 485.450 16.480 485.680 18.060 ;
        RECT 490.740 16.480 490.970 18.060 ;
        RECT 496.030 16.480 496.260 18.060 ;
        RECT 501.320 16.480 501.550 18.060 ;
        RECT 503.040 15.860 506.880 38.560 ;
        RECT 503.940 -15.670 506.880 15.860 ;
        RECT 937.040 -15.400 1093.980 -15.040 ;
        RECT 1142.020 -15.400 1172.890 -14.900 ;
        RECT 937.040 -15.670 1173.000 -15.400 ;
        RECT -106.870 -40.280 1173.000 -15.670 ;
        RECT -106.870 -40.400 1138.080 -40.280 ;
        RECT -106.870 -40.670 1093.980 -40.400 ;
        RECT -106.270 -41.090 -64.700 -40.670 ;
        RECT 937.040 -41.400 1093.980 -40.670 ;
      LAYER via ;
        RECT -90.935 349.760 -77.555 351.620 ;
        RECT 654.060 350.925 654.320 351.185 ;
        RECT 839.650 350.770 839.910 351.030 ;
        RECT 664.550 328.570 664.810 328.830 ;
        RECT 664.870 328.570 665.130 328.830 ;
        RECT 670.550 328.550 670.810 328.810 ;
        RECT 670.870 328.550 671.130 328.810 ;
        RECT 675.900 328.530 676.160 328.790 ;
        RECT 676.220 328.530 676.480 328.790 ;
        RECT 683.580 328.510 683.840 328.770 ;
        RECT 683.900 328.510 684.160 328.770 ;
        RECT 689.310 328.550 689.570 328.810 ;
        RECT 689.630 328.550 689.890 328.810 ;
        RECT 596.765 325.860 597.025 326.120 ;
        RECT 605.465 322.975 605.725 323.235 ;
        RECT 605.785 322.975 606.045 323.235 ;
        RECT 635.200 326.145 635.460 326.405 ;
        RECT 627.155 322.740 627.415 323.000 ;
        RECT 659.060 322.245 659.320 322.505 ;
        RECT 659.380 322.245 659.640 322.505 ;
        RECT 664.030 322.245 664.290 322.505 ;
        RECT 664.350 322.245 664.610 322.505 ;
        RECT 689.210 322.100 689.790 322.680 ;
        RECT 646.375 319.715 649.195 321.895 ;
        RECT 661.830 316.250 662.410 316.830 ;
        RECT 596.615 307.690 596.875 307.950 ;
        RECT 605.315 304.805 605.575 305.065 ;
        RECT 605.635 304.805 605.895 305.065 ;
        RECT 635.050 307.975 635.310 308.235 ;
        RECT 627.005 304.570 627.265 304.830 ;
        RECT 646.255 301.705 649.075 303.885 ;
        RECT 843.735 304.140 843.995 304.400 ;
        RECT 596.565 288.510 596.825 288.770 ;
        RECT 605.265 285.625 605.525 285.885 ;
        RECT 605.585 285.625 605.845 285.885 ;
        RECT 635.000 288.795 635.260 289.055 ;
        RECT 626.955 285.390 627.215 285.650 ;
        RECT 646.055 282.615 648.875 284.795 ;
        RECT 596.485 270.040 596.745 270.300 ;
        RECT 605.185 267.155 605.445 267.415 ;
        RECT 605.505 267.155 605.765 267.415 ;
        RECT 634.920 270.325 635.180 270.585 ;
        RECT 626.875 266.920 627.135 267.180 ;
        RECT 857.785 294.610 858.045 294.870 ;
        RECT 857.785 294.290 858.045 294.550 ;
        RECT 839.770 292.445 840.030 292.705 ;
        RECT 862.190 290.685 862.450 290.945 ;
        RECT 821.390 289.290 821.970 289.870 ;
        RECT 824.885 287.215 825.145 287.475 ;
        RECT 839.800 287.265 840.060 287.525 ;
        RECT 862.190 290.365 862.450 290.625 ;
        RECT 857.670 289.005 857.930 289.265 ;
        RECT 857.670 288.685 857.930 288.945 ;
        RECT 844.705 286.755 845.285 287.335 ;
        RECT 821.715 284.215 821.975 284.475 ;
        RECT 857.715 283.425 857.975 283.685 ;
        RECT 862.030 281.455 862.290 281.715 ;
        RECT 862.350 281.455 862.610 281.715 ;
        RECT 799.430 279.615 799.690 279.875 ;
        RECT 799.430 279.295 799.690 279.555 ;
        RECT 821.795 279.195 822.055 279.455 ;
        RECT 845.195 279.100 845.455 279.360 ;
        RECT 845.195 278.780 845.455 279.040 ;
        RECT 694.530 277.780 695.110 278.360 ;
        RECT 857.785 278.005 858.045 278.265 ;
        RECT 749.720 274.720 749.980 274.980 ;
        RECT 689.530 272.560 689.790 272.820 ;
        RECT 689.850 272.560 690.110 272.820 ;
        RECT 694.760 272.380 695.340 272.960 ;
        RECT 706.760 272.580 707.020 272.840 ;
        RECT 707.080 272.580 707.340 272.840 ;
        RECT 724.330 272.680 724.590 272.940 ;
        RECT 724.650 272.680 724.910 272.940 ;
        RECT 741.500 272.710 741.760 272.970 ;
        RECT 741.820 272.710 742.080 272.970 ;
        RECT 798.895 274.305 799.475 274.885 ;
        RECT 759.310 272.770 759.570 273.030 ;
        RECT 759.630 272.770 759.890 273.030 ;
        RECT 857.740 271.605 858.000 271.865 ;
        RECT 749.885 268.520 750.145 268.780 ;
        RECT 689.800 266.750 690.060 267.010 ;
        RECT 690.120 266.750 690.380 267.010 ;
        RECT 707.030 266.770 707.290 267.030 ;
        RECT 707.350 266.770 707.610 267.030 ;
        RECT 724.600 266.870 724.860 267.130 ;
        RECT 724.920 266.870 725.180 267.130 ;
        RECT 741.770 266.900 742.030 267.160 ;
        RECT 742.090 266.900 742.350 267.160 ;
        RECT 759.580 266.960 759.840 267.220 ;
        RECT 759.900 266.960 760.160 267.220 ;
        RECT 763.790 267.195 764.050 267.455 ;
        RECT 646.095 263.925 648.915 266.105 ;
        RECT 780.765 263.755 781.345 264.335 ;
        RECT 857.740 271.285 858.000 271.545 ;
        RECT 862.030 268.110 862.290 268.370 ;
        RECT 862.350 268.110 862.610 268.370 ;
        RECT 845.240 265.230 846.140 266.130 ;
        RECT 857.720 264.955 857.980 265.215 ;
        RECT 857.720 264.635 857.980 264.895 ;
        RECT 756.530 258.755 756.790 259.015 ;
        RECT 756.530 258.435 756.790 258.695 ;
        RECT 694.510 256.250 695.090 256.830 ;
        RECT 857.690 255.625 857.950 255.885 ;
        RECT 857.690 255.305 857.950 255.565 ;
        RECT 596.335 252.310 596.595 252.570 ;
        RECT 605.035 249.425 605.295 249.685 ;
        RECT 605.355 249.425 605.615 249.685 ;
        RECT 679.920 252.980 680.180 253.240 ;
        RECT 634.770 252.595 635.030 252.855 ;
        RECT 749.700 253.190 749.960 253.450 ;
        RECT 689.510 251.030 689.770 251.290 ;
        RECT 689.830 251.030 690.090 251.290 ;
        RECT 694.740 250.850 695.320 251.430 ;
        RECT 706.740 251.050 707.000 251.310 ;
        RECT 707.060 251.050 707.320 251.310 ;
        RECT 724.310 251.150 724.570 251.410 ;
        RECT 724.630 251.150 724.890 251.410 ;
        RECT 741.480 251.180 741.740 251.440 ;
        RECT 741.800 251.180 742.060 251.440 ;
        RECT 756.445 252.560 756.705 252.820 ;
        RECT 862.015 252.815 862.595 253.395 ;
        RECT 756.445 252.240 756.705 252.500 ;
        RECT 759.290 251.240 759.550 251.500 ;
        RECT 759.610 251.240 759.870 251.500 ;
        RECT 626.725 249.190 626.985 249.450 ;
        RECT 601.805 248.470 602.065 248.730 ;
        RECT 602.125 248.470 602.385 248.730 ;
        RECT 857.685 249.880 857.945 250.140 ;
        RECT 857.685 249.560 857.945 249.820 ;
        RECT 591.305 244.750 592.205 245.970 ;
        RECT 646.175 246.195 648.995 248.375 ;
        RECT 680.085 246.780 680.345 247.040 ;
        RECT 749.865 246.990 750.125 247.250 ;
        RECT 756.490 246.850 756.750 247.110 ;
        RECT 756.490 246.530 756.750 246.790 ;
        RECT 601.845 245.125 603.065 245.705 ;
        RECT 676.580 244.490 678.120 246.350 ;
        RECT 689.780 245.220 690.040 245.480 ;
        RECT 690.100 245.220 690.360 245.480 ;
        RECT 707.010 245.240 707.270 245.500 ;
        RECT 707.330 245.240 707.590 245.500 ;
        RECT 724.580 245.340 724.840 245.600 ;
        RECT 724.900 245.340 725.160 245.600 ;
        RECT 741.750 245.370 742.010 245.630 ;
        RECT 742.070 245.370 742.330 245.630 ;
        RECT 759.560 245.430 759.820 245.690 ;
        RECT 759.880 245.430 760.140 245.690 ;
        RECT 192.120 239.295 198.780 243.715 ;
        RECT -91.555 227.910 -78.175 230.410 ;
        RECT 341.135 237.160 344.275 239.020 ;
        RECT -90.925 215.790 -77.545 218.290 ;
        RECT -91.385 127.950 -78.005 130.450 ;
        RECT -90.645 8.740 -77.265 11.240 ;
        RECT -106.095 -41.070 -64.875 -15.530 ;
        RECT 442.880 213.345 448.900 218.405 ;
        RECT 610.345 -25.410 624.045 -17.150 ;
        RECT 703.215 -26.215 715.955 -17.635 ;
        RECT 790.550 -23.430 802.330 -17.090 ;
        RECT 860.960 -22.690 872.740 -16.350 ;
        RECT 928.940 -23.060 940.720 -16.720 ;
        RECT 1142.125 -39.300 1172.785 -15.040 ;
      LAYER met2 ;
        RECT -90.980 349.580 -77.510 351.800 ;
        RECT 653.960 351.300 654.420 351.390 ;
        RECT 647.140 350.850 654.420 351.300 ;
        RECT 647.140 350.320 648.090 350.850 ;
        RECT 653.960 350.720 654.420 350.850 ;
        RECT 839.580 351.130 839.980 351.160 ;
        RECT 839.580 351.110 848.180 351.130 ;
        RECT 839.580 350.770 849.220 351.110 ;
        RECT 839.580 350.640 839.980 350.770 ;
        RECT 596.610 325.790 597.180 326.190 ;
        RECT 635.130 326.050 635.530 326.500 ;
        RECT 596.740 323.150 596.930 325.790 ;
        RECT 605.390 323.150 606.120 323.400 ;
        RECT 596.740 323.000 606.120 323.150 ;
        RECT 605.390 322.810 606.120 323.000 ;
        RECT 627.060 322.990 627.510 323.190 ;
        RECT 635.200 322.990 635.420 326.050 ;
        RECT 627.060 322.780 635.420 322.990 ;
        RECT 627.060 322.550 627.510 322.780 ;
        RECT 635.200 322.760 635.420 322.780 ;
        RECT 647.180 322.050 648.070 350.320 ;
        RECT 664.510 328.840 665.170 329.000 ;
        RECT 670.510 328.840 671.170 328.980 ;
        RECT 675.860 328.840 676.520 328.960 ;
        RECT 683.540 328.840 684.200 328.940 ;
        RECT 689.270 328.840 689.930 328.980 ;
        RECT 664.510 328.490 689.930 328.840 ;
        RECT 664.510 328.400 665.170 328.490 ;
        RECT 670.510 328.380 671.170 328.490 ;
        RECT 675.860 328.360 676.520 328.490 ;
        RECT 683.540 328.340 684.200 328.490 ;
        RECT 689.270 328.380 689.930 328.490 ;
        RECT 659.010 322.690 659.650 322.900 ;
        RECT 689.350 322.740 689.660 328.380 ;
        RECT 659.010 322.520 659.670 322.690 ;
        RECT 664.000 322.520 664.640 322.690 ;
        RECT 659.010 322.280 664.640 322.520 ;
        RECT 659.010 322.060 659.670 322.280 ;
        RECT 664.000 322.060 664.640 322.280 ;
        RECT 646.230 319.560 649.340 322.050 ;
        RECT 659.010 322.000 659.650 322.060 ;
        RECT 689.120 322.040 689.880 322.740 ;
        RECT 647.060 317.390 648.140 319.560 ;
        RECT 649.560 317.390 653.640 317.410 ;
        RECT 656.230 317.390 657.580 317.990 ;
        RECT 647.060 316.840 657.580 317.390 ;
        RECT 596.460 307.620 597.030 308.020 ;
        RECT 634.980 307.880 635.380 308.330 ;
        RECT 596.590 304.980 596.780 307.620 ;
        RECT 605.240 304.980 605.970 305.230 ;
        RECT 596.590 304.830 605.970 304.980 ;
        RECT 605.240 304.640 605.970 304.830 ;
        RECT 626.910 304.820 627.360 305.020 ;
        RECT 635.050 304.820 635.270 307.880 ;
        RECT 626.910 304.610 635.270 304.820 ;
        RECT 626.910 304.380 627.360 304.610 ;
        RECT 635.050 304.590 635.270 304.610 ;
        RECT 647.060 304.040 648.140 316.840 ;
        RECT 649.560 316.760 653.640 316.840 ;
        RECT 656.230 316.480 657.580 316.840 ;
        RECT 661.740 316.160 662.500 316.920 ;
        RECT 843.670 304.270 844.060 304.570 ;
        RECT 848.330 304.270 849.220 350.770 ;
        RECT 843.670 304.060 849.220 304.270 ;
        RECT 843.670 304.050 849.040 304.060 ;
        RECT 646.110 301.550 649.220 304.040 ;
        RECT 843.670 303.970 844.060 304.050 ;
        RECT 596.410 288.440 596.980 288.840 ;
        RECT 634.930 288.700 635.330 289.150 ;
        RECT 596.540 285.800 596.730 288.440 ;
        RECT 605.190 285.800 605.920 286.050 ;
        RECT 596.540 285.650 605.920 285.800 ;
        RECT 605.190 285.460 605.920 285.650 ;
        RECT 626.860 285.640 627.310 285.840 ;
        RECT 635.000 285.640 635.220 288.700 ;
        RECT 626.860 285.430 635.220 285.640 ;
        RECT 626.860 285.200 627.310 285.430 ;
        RECT 635.000 285.410 635.220 285.430 ;
        RECT 647.060 284.950 648.140 301.550 ;
        RECT 857.700 294.220 858.130 294.940 ;
        RECT 839.620 292.250 840.180 292.900 ;
        RECT 821.390 289.240 821.970 289.920 ;
        RECT 839.810 287.720 840.070 292.250 ;
        RECT 857.700 289.330 857.980 294.220 ;
        RECT 862.040 290.290 862.600 291.020 ;
        RECT 857.640 289.150 857.980 289.330 ;
        RECT 857.640 288.800 857.960 289.150 ;
        RECT 857.640 288.620 857.980 288.800 ;
        RECT 824.750 287.020 825.280 287.670 ;
        RECT 839.650 287.070 840.210 287.720 ;
        RECT 844.660 286.600 845.330 287.490 ;
        RECT 845.010 286.240 845.270 286.600 ;
        RECT 844.920 285.750 845.750 286.240 ;
        RECT 645.910 282.460 649.020 284.950 ;
        RECT 821.610 284.010 822.080 284.680 ;
        RECT 857.700 283.890 857.980 288.620 ;
        RECT 845.070 283.220 845.660 283.730 ;
        RECT 857.610 283.220 858.080 283.890 ;
        RECT 596.330 269.970 596.900 270.370 ;
        RECT 634.850 270.230 635.250 270.680 ;
        RECT 596.460 267.330 596.650 269.970 ;
        RECT 605.110 267.330 605.840 267.580 ;
        RECT 596.460 267.180 605.840 267.330 ;
        RECT 605.110 266.990 605.840 267.180 ;
        RECT 626.780 267.170 627.230 267.370 ;
        RECT 634.920 267.170 635.140 270.230 ;
        RECT 626.780 266.960 635.140 267.170 ;
        RECT 626.780 266.730 627.230 266.960 ;
        RECT 634.920 266.940 635.140 266.960 ;
        RECT 647.060 266.260 648.140 282.460 ;
        RECT 799.300 279.190 799.820 279.980 ;
        RECT 694.530 277.630 695.110 278.510 ;
        RECT 694.830 273.110 695.100 277.630 ;
        RECT 749.620 274.550 750.080 275.150 ;
        RECT 799.310 274.990 799.650 279.190 ;
        RECT 821.690 278.990 822.160 279.660 ;
        RECT 845.220 279.440 845.410 283.220 ;
        RECT 845.090 278.700 845.560 279.440 ;
        RECT 857.770 278.470 857.980 283.220 ;
        RECT 862.210 281.900 862.410 290.290 ;
        RECT 861.970 281.270 862.670 281.900 ;
        RECT 857.680 277.800 858.150 278.470 ;
        RECT 798.850 274.680 799.650 274.990 ;
        RECT 689.530 272.370 690.110 273.010 ;
        RECT 689.880 267.200 690.060 272.370 ;
        RECT 694.760 272.230 695.340 273.110 ;
        RECT 706.760 272.390 707.340 273.030 ;
        RECT 724.330 272.490 724.910 273.130 ;
        RECT 741.500 272.520 742.080 273.160 ;
        RECT 707.110 267.220 707.290 272.390 ;
        RECT 724.680 267.320 724.860 272.490 ;
        RECT 741.850 267.350 742.030 272.520 ;
        RECT 749.870 268.920 750.050 274.550 ;
        RECT 798.850 274.200 799.520 274.680 ;
        RECT 759.310 272.580 759.890 273.220 ;
        RECT 749.810 268.380 750.220 268.920 ;
        RECT 759.660 267.410 759.840 272.580 ;
        RECT 857.730 271.920 857.980 277.800 ;
        RECT 857.630 271.230 858.110 271.920 ;
        RECT 689.800 266.560 690.380 267.200 ;
        RECT 707.030 266.580 707.610 267.220 ;
        RECT 724.600 266.680 725.180 267.320 ;
        RECT 741.770 266.710 742.350 267.350 ;
        RECT 759.580 266.770 760.160 267.410 ;
        RECT 763.670 267.340 764.170 267.650 ;
        RECT 763.670 267.000 764.410 267.340 ;
        RECT 645.950 263.770 649.060 266.260 ;
        RECT 763.940 264.350 764.410 267.000 ;
        RECT 845.190 265.110 846.190 266.250 ;
        RECT 857.730 265.270 857.960 271.230 ;
        RECT 862.190 268.550 862.380 281.270 ;
        RECT 861.950 267.930 862.690 268.550 ;
        RECT 845.600 264.550 845.950 265.110 ;
        RECT 857.610 264.580 858.090 265.270 ;
        RECT 845.600 264.440 857.470 264.550 ;
        RECT 857.630 264.440 857.910 264.580 ;
        RECT 780.730 264.350 781.380 264.440 ;
        RECT 763.940 264.130 781.380 264.350 ;
        RECT 845.600 264.260 857.910 264.440 ;
        RECT 193.050 249.330 194.820 252.410 ;
        RECT 596.180 252.240 596.750 252.640 ;
        RECT 634.700 252.500 635.100 252.950 ;
        RECT 192.670 248.210 195.590 249.330 ;
        RECT 192.700 243.870 195.590 248.210 ;
        RECT 340.850 247.330 344.510 250.110 ;
        RECT 596.310 249.600 596.500 252.240 ;
        RECT 604.960 249.600 605.690 249.850 ;
        RECT 596.310 249.450 605.690 249.600 ;
        RECT 604.960 249.260 605.690 249.450 ;
        RECT 626.630 249.440 627.080 249.640 ;
        RECT 634.770 249.440 634.990 252.500 ;
        RECT 626.630 249.230 634.990 249.440 ;
        RECT 626.630 249.000 627.080 249.230 ;
        RECT 634.770 249.210 634.990 249.230 ;
        RECT 601.680 248.390 602.510 248.810 ;
        RECT 647.060 248.530 648.140 263.770 ;
        RECT 780.730 263.650 781.380 264.130 ;
        RECT 756.380 258.370 756.940 259.080 ;
        RECT 756.450 258.240 756.690 258.370 ;
        RECT 694.510 256.100 695.090 256.980 ;
        RECT 679.820 252.810 680.280 253.410 ;
        RECT 192.120 239.140 198.780 243.870 ;
        RECT 341.560 239.110 343.100 247.330 ;
        RECT 646.030 246.690 649.140 248.530 ;
        RECT 680.070 247.180 680.250 252.810 ;
        RECT 694.810 251.580 695.080 256.100 ;
        RECT 749.600 253.020 750.060 253.620 ;
        RECT 689.510 250.840 690.090 251.480 ;
        RECT 646.030 246.500 677.100 246.690 ;
        RECT 680.010 246.640 680.420 247.180 ;
        RECT 591.180 244.610 592.330 246.110 ;
        RECT 646.030 246.040 678.200 246.500 ;
        RECT 647.840 245.910 678.200 246.040 ;
        RECT 601.720 245.050 603.190 245.780 ;
        RECT 676.500 244.340 678.200 245.910 ;
        RECT 689.860 245.670 690.040 250.840 ;
        RECT 694.740 250.700 695.320 251.580 ;
        RECT 706.740 250.860 707.320 251.500 ;
        RECT 724.310 250.960 724.890 251.600 ;
        RECT 741.480 250.990 742.060 251.630 ;
        RECT 707.090 245.690 707.270 250.860 ;
        RECT 724.660 245.790 724.840 250.960 ;
        RECT 741.830 245.820 742.010 250.990 ;
        RECT 749.850 247.390 750.030 253.020 ;
        RECT 756.450 252.990 756.670 258.240 ;
        RECT 857.630 255.940 857.910 264.260 ;
        RECT 857.570 255.250 858.070 255.940 ;
        RECT 756.330 252.070 756.820 252.990 ;
        RECT 749.790 246.850 750.200 247.390 ;
        RECT 756.490 247.160 756.660 252.070 ;
        RECT 759.290 251.050 759.870 251.690 ;
        RECT 756.440 246.480 756.800 247.160 ;
        RECT 759.640 245.880 759.820 251.050 ;
        RECT 857.750 250.190 857.910 255.250 ;
        RECT 862.170 253.450 862.410 267.930 ;
        RECT 861.990 252.760 862.620 253.450 ;
        RECT 857.540 249.510 858.090 250.190 ;
        RECT 689.780 245.030 690.360 245.670 ;
        RECT 707.010 245.050 707.590 245.690 ;
        RECT 724.580 245.150 725.160 245.790 ;
        RECT 741.750 245.180 742.330 245.820 ;
        RECT 759.560 245.240 760.140 245.880 ;
        RECT 340.990 237.070 344.420 239.110 ;
        RECT -91.610 227.800 -78.120 230.520 ;
        RECT 443.540 226.200 448.930 229.140 ;
        RECT 444.910 218.470 447.070 226.200 ;
        RECT -90.980 215.680 -77.490 218.400 ;
        RECT 442.760 213.280 449.020 218.470 ;
        RECT -91.440 127.840 -77.950 130.560 ;
        RECT -90.700 8.630 -77.210 11.350 ;
        RECT -106.220 -41.140 -64.750 -15.460 ;
        RECT 610.340 -25.590 624.050 -16.970 ;
        RECT 703.100 -26.330 716.070 -17.520 ;
        RECT 790.400 -23.560 802.480 -16.960 ;
        RECT 860.810 -22.820 872.890 -16.220 ;
        RECT 928.790 -23.190 940.870 -16.590 ;
        RECT 1142.070 -39.490 1172.840 -14.850 ;
      LAYER via2 ;
        RECT -90.785 349.750 -77.705 351.630 ;
        RECT 659.190 322.510 659.470 322.790 ;
        RECT 659.190 322.110 659.470 322.390 ;
        RECT 656.365 316.695 657.445 317.775 ;
        RECT 661.780 316.400 662.060 316.680 ;
        RECT 662.180 316.400 662.460 316.680 ;
        RECT 821.540 289.440 821.820 289.720 ;
        RECT 824.875 287.205 825.155 287.485 ;
        RECT 844.995 285.855 845.275 286.135 ;
        RECT 845.395 285.855 845.675 286.135 ;
        RECT 821.705 284.205 821.985 284.485 ;
        RECT 845.225 283.335 845.505 283.615 ;
        RECT 821.785 279.185 822.065 279.465 ;
        RECT 193.195 249.210 194.675 252.290 ;
        RECT 340.940 247.380 344.420 250.060 ;
        RECT 601.755 248.460 602.035 248.740 ;
        RECT 602.155 248.460 602.435 248.740 ;
        RECT 591.215 244.820 592.295 245.900 ;
        RECT 601.915 245.275 602.195 245.555 ;
        RECT 602.315 245.275 602.595 245.555 ;
        RECT 602.715 245.275 602.995 245.555 ;
        RECT -91.605 228.020 -78.125 230.300 ;
        RECT 443.695 226.330 448.775 229.010 ;
        RECT -90.975 215.900 -77.495 218.180 ;
        RECT -91.435 128.060 -77.955 130.340 ;
        RECT -90.695 8.850 -77.215 11.130 ;
        RECT -106.025 -41.040 -64.945 -15.560 ;
        RECT 610.455 -25.420 623.935 -17.140 ;
        RECT 703.245 -26.265 715.925 -17.585 ;
        RECT 790.500 -23.400 802.380 -17.120 ;
        RECT 860.910 -22.660 872.790 -16.380 ;
        RECT 928.890 -23.030 940.770 -16.750 ;
        RECT 1142.115 -39.310 1172.795 -15.030 ;
      LAYER met3 ;
        RECT 1067.150 465.190 1172.740 466.100 ;
        RECT 1067.150 464.850 1172.790 465.190 ;
        RECT 935.630 463.770 1172.790 464.850 ;
        RECT 935.630 463.500 1173.090 463.770 ;
        RECT -107.100 462.100 1173.090 463.500 ;
        RECT -108.550 429.310 1173.090 462.100 ;
        RECT -108.550 429.040 1172.740 429.310 ;
        RECT -108.550 428.340 -4.380 429.040 ;
        RECT 935.630 428.890 1172.740 429.040 ;
        RECT 1067.150 428.850 1172.740 428.890 ;
        RECT -91.030 349.605 -77.460 351.775 ;
        RECT 164.400 339.390 190.600 343.470 ;
        RECT 164.220 323.170 190.660 339.390 ;
        RECT 164.220 322.920 193.150 323.170 ;
        RECT 164.220 320.610 194.420 322.920 ;
        RECT 164.220 301.770 190.660 320.610 ;
        RECT 192.540 301.770 194.420 320.610 ;
        RECT 164.220 299.210 194.420 301.770 ;
        RECT 164.220 280.450 190.660 299.210 ;
        RECT 192.540 280.450 194.420 299.210 ;
        RECT 312.180 308.100 338.620 325.840 ;
        RECT 658.960 322.025 659.700 322.875 ;
        RECT 656.180 317.410 657.630 317.965 ;
        RECT 659.200 317.410 659.630 322.025 ;
        RECT 656.180 316.860 659.650 317.410 ;
        RECT 656.180 316.505 657.630 316.860 ;
        RECT 659.200 316.710 659.650 316.860 ;
        RECT 661.690 316.710 662.550 316.895 ;
        RECT 659.200 316.340 662.550 316.710 ;
        RECT 661.690 316.185 662.550 316.340 ;
        RECT 312.180 305.460 338.850 308.100 ;
        RECT 312.180 300.240 338.620 305.460 ;
        RECT 312.180 297.540 343.290 300.240 ;
        RECT 312.180 286.690 338.620 297.540 ;
        RECT 312.180 284.050 338.850 286.690 ;
        RECT 164.220 277.810 194.480 280.450 ;
        RECT 312.180 278.200 338.620 284.050 ;
        RECT 340.690 278.200 343.270 297.540 ;
        RECT 821.340 289.265 822.020 289.895 ;
        RECT 821.550 287.530 821.850 289.265 ;
        RECT 824.700 287.530 825.330 287.645 ;
        RECT 821.550 287.220 825.330 287.530 ;
        RECT 821.550 284.655 821.850 287.220 ;
        RECT 824.700 287.045 825.330 287.220 ;
        RECT 844.870 285.775 845.800 286.215 ;
        RECT 821.550 284.420 822.130 284.655 ;
        RECT 821.560 284.035 822.130 284.420 ;
        RECT 821.790 279.635 822.130 284.035 ;
        RECT 845.180 283.705 845.500 285.775 ;
        RECT 845.020 283.245 845.710 283.705 ;
        RECT 821.640 279.015 822.210 279.635 ;
        RECT 164.220 259.040 190.660 277.810 ;
        RECT 192.540 259.040 194.420 277.810 ;
        RECT 312.180 276.350 343.270 278.200 ;
        RECT 312.180 276.080 342.750 276.350 ;
        RECT 312.360 276.020 342.750 276.080 ;
        RECT 164.220 256.400 194.730 259.040 ;
        RECT 312.360 258.240 338.560 276.020 ;
        RECT 341.600 266.160 342.750 276.020 ;
        RECT 164.220 248.430 190.660 256.400 ;
        RECT 192.540 256.370 194.730 256.400 ;
        RECT 192.990 252.385 194.730 256.370 ;
        RECT 192.990 252.160 194.870 252.385 ;
        RECT 193.000 249.115 194.870 252.160 ;
        RECT 341.600 250.085 342.880 266.160 ;
        RECT 415.620 260.070 442.060 262.670 ;
        RECT 415.620 257.370 443.010 260.070 ;
        RECT 164.400 230.590 190.600 248.430 ;
        RECT 340.800 247.355 344.560 250.085 ;
        RECT 415.620 246.520 442.060 257.370 ;
        RECT 601.630 248.415 602.560 248.785 ;
        RECT 415.620 243.880 442.290 246.520 ;
        RECT 591.130 245.570 592.380 246.085 ;
        RECT 599.280 245.570 600.320 245.830 ;
        RECT 601.770 245.755 602.330 248.415 ;
        RECT 601.670 245.570 603.240 245.755 ;
        RECT 591.130 245.075 603.240 245.570 ;
        RECT 591.130 245.060 602.210 245.075 ;
        RECT 591.130 244.635 592.380 245.060 ;
        RECT 415.620 238.700 442.060 243.880 ;
        RECT 599.240 240.570 600.320 245.060 ;
        RECT 415.620 238.210 447.320 238.700 ;
        RECT 415.620 235.910 447.360 238.210 ;
        RECT 415.800 235.470 447.360 235.910 ;
        RECT -91.660 227.825 -78.070 230.495 ;
        RECT -91.030 215.705 -77.440 218.375 ;
        RECT 415.800 218.070 442.000 235.470 ;
        RECT 444.520 229.115 447.360 235.470 ;
        RECT 443.490 226.225 448.980 229.115 ;
        RECT 599.240 221.970 600.240 240.570 ;
        RECT -91.490 127.865 -77.900 130.535 ;
        RECT 555.690 81.850 1017.970 221.970 ;
        RECT 586.130 80.780 596.190 81.850 ;
        RECT 612.950 45.590 617.530 81.850 ;
        RECT 706.970 54.420 711.770 81.850 ;
        RECT 793.150 54.420 797.950 81.850 ;
        RECT 863.830 54.420 868.630 81.850 ;
        RECT 931.680 54.420 936.480 81.850 ;
        RECT -90.750 8.655 -77.160 11.325 ;
        RECT -106.270 -41.115 -64.700 -15.485 ;
        RECT 613.410 -16.995 617.110 45.590 ;
        RECT 706.340 41.660 711.770 54.420 ;
        RECT 610.290 -25.565 624.100 -16.995 ;
        RECT 706.340 -17.545 711.530 41.660 ;
        RECT 793.100 -16.985 798.290 54.420 ;
        RECT 863.410 46.900 868.630 54.420 ;
        RECT 863.410 -16.245 868.600 46.900 ;
        RECT 703.050 -26.305 716.120 -17.545 ;
        RECT 790.350 -23.535 802.530 -16.985 ;
        RECT 860.760 -22.795 872.940 -16.245 ;
        RECT 931.400 -16.615 936.590 54.420 ;
        RECT 928.740 -23.165 940.920 -16.615 ;
        RECT 1142.020 -39.465 1172.890 -14.875 ;
      LAYER via3 ;
        RECT -108.425 428.460 -4.505 461.980 ;
        RECT 1072.700 431.550 1172.620 465.070 ;
        RECT -90.805 349.730 -77.685 351.650 ;
        RECT -91.425 228.000 -78.305 230.320 ;
        RECT -90.795 215.880 -77.675 218.200 ;
        RECT -91.255 128.040 -78.135 130.360 ;
        RECT -90.515 8.830 -77.395 11.150 ;
        RECT -106.045 -41.060 -64.925 -15.540 ;
        RECT 1142.095 -39.330 1172.815 -15.010 ;
      LAYER met4 ;
        RECT -22.640 462.105 -11.970 489.770 ;
        RECT 1067.150 465.195 1172.740 466.100 ;
        RECT -108.505 428.335 -4.425 462.105 ;
        RECT 1067.150 431.425 1172.745 465.195 ;
        RECT 1067.150 428.850 1172.740 431.425 ;
        RECT -105.550 -15.505 -68.700 428.335 ;
        RECT 1145.400 -14.895 1172.570 428.850 ;
        RECT -106.225 -16.260 -64.745 -15.505 ;
        RECT -106.225 -41.010 -64.550 -16.260 ;
        RECT 1142.065 -28.590 1172.845 -14.895 ;
        RECT 1141.160 -39.445 1172.845 -28.590 ;
        RECT 1141.160 -40.280 1172.620 -39.445 ;
        RECT -106.225 -41.095 -64.745 -41.010 ;
    END
  END vssa2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 352.710 376.120 411.040 377.760 ;
        RECT 352.710 375.150 411.110 376.120 ;
        RECT 352.860 371.270 411.110 375.150 ;
        RECT -53.480 351.095 -25.390 358.715 ;
        RECT 0.310 300.440 106.070 331.780 ;
        RECT 208.370 326.960 291.730 370.320 ;
        RECT 352.970 368.120 411.110 371.270 ;
        RECT 352.970 367.890 411.130 368.120 ;
        RECT 0.170 297.450 106.070 300.440 ;
        RECT 208.270 322.310 291.730 326.960 ;
        RECT -53.470 229.715 -25.380 237.335 ;
        RECT 0.170 234.280 105.930 297.450 ;
        RECT 208.270 284.020 291.630 322.310 ;
        RECT 207.990 278.950 291.630 284.020 ;
        RECT 207.990 236.010 291.350 278.950 ;
        RECT 352.980 254.470 411.130 367.890 ;
        RECT 653.640 355.340 655.740 355.345 ;
        RECT 653.640 355.335 657.550 355.340 ;
        RECT 653.640 355.310 673.240 355.335 ;
        RECT 690.870 355.315 693.280 355.320 ;
        RECT 708.710 355.315 710.910 355.320 ;
        RECT 726.550 355.315 729.260 355.330 ;
        RECT 653.640 355.295 675.610 355.310 ;
        RECT 690.870 355.295 744.990 355.315 ;
        RECT 653.640 355.290 744.990 355.295 ;
        RECT 653.640 355.285 747.000 355.290 ;
        RECT 653.640 355.130 762.760 355.285 ;
        RECT 782.940 355.240 798.960 355.245 ;
        RECT 801.320 355.240 817.340 355.255 ;
        RECT 782.940 355.235 820.290 355.240 ;
        RECT 782.940 355.230 836.140 355.235 ;
        RECT 782.940 355.215 838.930 355.230 ;
        RECT 782.940 355.210 840.690 355.215 ;
        RECT 780.590 355.205 840.690 355.210 ;
        RECT 764.780 355.130 840.690 355.205 ;
        RECT 653.640 352.750 840.690 355.130 ;
        RECT 653.640 352.745 673.240 352.750 ;
        RECT 655.490 352.735 673.240 352.745 ;
        RECT 655.490 352.720 657.550 352.735 ;
        RECT 675.270 352.720 840.690 352.750 ;
        RECT 675.270 352.715 726.730 352.720 ;
        RECT 728.970 352.715 840.690 352.720 ;
        RECT 675.270 352.695 693.280 352.715 ;
        RECT 708.710 352.700 710.910 352.715 ;
        RECT 744.720 352.710 840.690 352.715 ;
        RECT 690.870 352.690 693.280 352.695 ;
        RECT 746.740 352.690 840.690 352.710 ;
        RECT 746.740 352.685 762.760 352.690 ;
        RECT 764.780 352.670 840.690 352.690 ;
        RECT 764.780 352.655 817.340 352.670 ;
        RECT 764.780 352.645 801.590 352.655 ;
        RECT 764.780 352.605 783.170 352.645 ;
        RECT 798.730 352.640 801.590 352.645 ;
        RECT 820.120 352.635 840.690 352.670 ;
        RECT 780.590 352.580 783.170 352.605 ;
        RECT 835.880 352.615 840.690 352.635 ;
        RECT 835.880 352.590 838.930 352.615 ;
        RECT 791.530 347.165 794.160 347.180 ;
        RECT 791.530 347.110 809.540 347.165 ;
        RECT 791.530 347.105 813.160 347.110 ;
        RECT 790.060 347.075 813.160 347.105 ;
        RECT 828.740 347.075 830.460 347.120 ;
        RECT 783.500 347.070 787.520 347.075 ;
        RECT 790.060 347.070 830.460 347.075 ;
        RECT 783.500 344.580 830.460 347.070 ;
        RECT 783.500 344.565 809.540 344.580 ;
        RECT 783.500 344.530 794.160 344.565 ;
        RECT 783.500 344.505 792.160 344.530 ;
        RECT 783.500 344.475 790.340 344.505 ;
        RECT 812.880 344.475 830.460 344.580 ;
        RECT 787.370 344.470 790.340 344.475 ;
        RECT 828.740 344.440 830.460 344.475 ;
        RECT 595.040 328.595 597.140 331.195 ;
        RECT 600.430 328.610 631.350 334.660 ;
        RECT 666.620 332.985 668.720 333.000 ;
        RECT 662.860 332.980 672.510 332.985 ;
        RECT 662.860 332.885 674.600 332.980 ;
        RECT 678.080 332.925 681.690 332.970 ;
        RECT 685.110 332.935 687.790 332.940 ;
        RECT 685.110 332.925 691.160 332.935 ;
        RECT 678.080 332.885 691.160 332.925 ;
        RECT 634.930 329.045 637.030 331.645 ;
        RECT 639.120 329.135 641.220 331.735 ;
        RECT 645.080 331.715 646.440 331.720 ;
        RECT 643.220 329.120 646.440 331.715 ;
        RECT 662.860 330.385 691.160 332.885 ;
        RECT 856.270 331.170 868.120 332.150 ;
        RECT 856.220 330.950 868.120 331.170 ;
        RECT 856.220 330.490 868.100 330.950 ;
        RECT 666.620 330.320 667.720 330.385 ;
        RECT 672.160 330.350 691.160 330.385 ;
        RECT 674.250 330.335 691.160 330.350 ;
        RECT 674.250 330.325 687.790 330.335 ;
        RECT 674.250 330.285 681.690 330.325 ;
        RECT 685.110 330.320 687.790 330.325 ;
        RECT 678.080 330.220 681.690 330.285 ;
        RECT 856.200 330.130 868.100 330.490 ;
        RECT 643.220 329.115 645.320 329.120 ;
        RECT 600.410 327.640 631.350 328.610 ;
        RECT 600.410 322.360 604.880 327.640 ;
        RECT 626.890 326.230 631.350 327.640 ;
        RECT 690.400 326.685 693.130 326.690 ;
        RECT 626.890 322.980 631.460 326.230 ;
        RECT 658.430 324.085 660.530 326.685 ;
        RECT 663.330 324.045 665.430 326.645 ;
        RECT 667.920 326.620 670.020 326.675 ;
        RECT 673.870 326.665 676.560 326.670 ;
        RECT 679.660 326.665 682.390 326.670 ;
        RECT 685.100 326.665 687.700 326.670 ;
        RECT 690.400 326.665 696.440 326.685 ;
        RECT 673.870 326.655 696.440 326.665 ;
        RECT 672.460 326.620 696.440 326.655 ;
        RECT 667.920 324.360 696.440 326.620 ;
        RECT 667.920 324.075 670.020 324.360 ;
        RECT 672.460 324.085 696.440 324.360 ;
        RECT 672.460 324.065 693.130 324.085 ;
        RECT 672.460 324.055 676.560 324.065 ;
        RECT 673.870 324.050 676.560 324.055 ;
        RECT 679.660 324.050 682.390 324.065 ;
        RECT 685.100 324.060 687.700 324.065 ;
        RECT 690.400 324.050 693.130 324.065 ;
        RECT 856.150 323.280 868.100 330.130 ;
        RECT 626.890 322.410 631.350 322.980 ;
        RECT 675.630 320.825 678.350 320.830 ;
        RECT 680.990 320.825 683.680 320.830 ;
        RECT 686.780 320.825 689.040 320.830 ;
        RECT 672.330 320.820 689.040 320.825 ;
        RECT 664.890 320.815 667.600 320.820 ;
        RECT 670.320 320.815 689.040 320.820 ;
        RECT 664.890 320.805 689.040 320.815 ;
        RECT 691.220 320.805 693.900 320.810 ;
        RECT 661.070 318.225 696.280 320.805 ;
        RECT 661.070 318.215 672.920 318.225 ;
        RECT 675.630 318.220 678.350 318.225 ;
        RECT 680.990 318.220 683.680 318.225 ;
        RECT 686.780 318.220 696.280 318.225 ;
        RECT 661.070 318.205 667.600 318.215 ;
        RECT 670.320 318.210 672.920 318.215 ;
        RECT 688.820 318.205 696.280 318.220 ;
        RECT 664.890 318.200 667.600 318.205 ;
        RECT 691.220 318.200 693.900 318.205 ;
        RECT 594.890 310.425 596.990 313.025 ;
        RECT 600.280 310.440 631.200 316.490 ;
        RECT 856.150 313.600 872.700 323.280 ;
        RECT 634.780 310.875 636.880 313.475 ;
        RECT 638.970 310.965 641.070 313.565 ;
        RECT 645.050 313.545 646.410 313.570 ;
        RECT 643.070 310.970 646.410 313.545 ;
        RECT 856.150 313.270 864.130 313.600 ;
        RECT 643.070 310.945 645.170 310.970 ;
        RECT 600.260 309.470 631.200 310.440 ;
        RECT 600.260 304.190 604.730 309.470 ;
        RECT 626.740 308.060 631.200 309.470 ;
        RECT 833.100 308.545 835.550 308.560 ;
        RECT 840.800 308.545 842.810 308.560 ;
        RECT 833.100 308.530 844.460 308.545 ;
        RECT 811.900 308.515 814.190 308.520 ;
        RECT 829.450 308.515 844.460 308.530 ;
        RECT 626.740 304.810 631.310 308.060 ;
        RECT 796.150 305.945 844.460 308.515 ;
        RECT 796.150 305.915 835.550 305.945 ;
        RECT 811.900 305.910 814.190 305.915 ;
        RECT 829.450 305.910 835.550 305.915 ;
        RECT 831.450 305.900 835.550 305.910 ;
        RECT 840.800 305.900 842.810 305.945 ;
        RECT 831.450 305.885 833.550 305.900 ;
        RECT 626.740 304.240 631.200 304.810 ;
        RECT 679.730 299.420 695.750 299.455 ;
        RECT 714.830 299.440 730.850 299.475 ;
        RECT 712.840 299.430 730.850 299.440 ;
        RECT 712.840 299.425 732.870 299.430 ;
        RECT 748.270 299.425 750.570 299.430 ;
        RECT 679.730 299.415 697.750 299.420 ;
        RECT 712.840 299.415 750.570 299.425 ;
        RECT 594.840 291.245 596.940 293.845 ;
        RECT 600.230 291.260 631.150 297.310 ;
        RECT 679.730 296.875 766.290 299.415 ;
        RECT 859.300 298.775 861.710 298.820 ;
        RECT 679.730 296.855 715.270 296.875 ;
        RECT 730.520 296.870 766.290 296.875 ;
        RECT 695.210 296.850 715.270 296.855 ;
        RECT 697.220 296.815 715.270 296.850 ;
        RECT 732.530 296.830 766.290 296.870 ;
        RECT 732.530 296.825 748.550 296.830 ;
        RECT 750.270 296.815 766.290 296.830 ;
        RECT 712.840 296.800 715.270 296.815 ;
        RECT 842.940 296.795 845.410 296.810 ;
        RECT 839.060 295.145 845.410 296.795 ;
        RECT 855.470 296.175 861.710 298.775 ;
        RECT 634.730 291.695 636.830 294.295 ;
        RECT 638.920 291.785 641.020 294.385 ;
        RECT 645.030 294.365 646.390 294.380 ;
        RECT 643.020 291.780 646.390 294.365 ;
        RECT 839.060 294.195 848.780 295.145 ;
        RECT 842.760 294.190 848.780 294.195 ;
        RECT 822.340 293.785 824.550 293.800 ;
        RECT 818.610 292.090 824.550 293.785 ;
        RECT 843.460 292.545 848.780 294.190 ;
        RECT 860.440 294.875 861.710 296.175 ;
        RECT 860.440 293.510 864.870 294.875 ;
        RECT 859.330 293.245 864.870 293.510 ;
        RECT 843.460 292.540 845.310 292.545 ;
        RECT 643.020 291.765 645.120 291.780 ;
        RECT 600.210 290.290 631.150 291.260 ;
        RECT 818.610 291.615 824.890 292.090 ;
        RECT 843.460 291.680 844.810 292.540 ;
        RECT 842.970 291.675 844.810 291.680 ;
        RECT 827.590 291.635 830.080 291.640 ;
        RECT 827.590 291.615 835.540 291.635 ;
        RECT 818.610 291.185 835.540 291.615 ;
        RECT 822.570 291.180 835.540 291.185 ;
        RECT 600.210 285.010 604.680 290.290 ;
        RECT 626.690 288.880 631.150 290.290 ;
        RECT 823.350 289.035 835.540 291.180 ;
        RECT 839.070 290.540 844.810 291.675 ;
        RECT 855.510 292.275 864.870 293.245 ;
        RECT 855.510 292.270 860.990 292.275 ;
        RECT 855.510 290.645 859.530 292.270 ;
        RECT 839.070 289.075 843.090 290.540 ;
        RECT 823.350 289.020 830.080 289.035 ;
        RECT 823.350 289.015 828.080 289.020 ;
        RECT 626.690 285.630 631.260 288.880 ;
        RECT 823.350 288.630 824.230 289.015 ;
        RECT 822.550 288.625 824.230 288.630 ;
        RECT 818.580 288.320 824.230 288.625 ;
        RECT 818.580 288.180 824.210 288.320 ;
        RECT 818.580 287.750 824.200 288.180 ;
        RECT 818.580 287.680 823.490 287.750 ;
        RECT 818.580 286.025 822.600 287.680 ;
        RECT 855.580 287.140 859.600 287.845 ;
        RECT 855.580 285.825 861.790 287.140 ;
        RECT 626.690 285.060 631.150 285.630 ;
        RECT 855.580 285.245 864.950 285.825 ;
        RECT 859.300 285.220 864.950 285.245 ;
        RECT 684.660 282.715 686.360 282.740 ;
        RECT 702.000 282.725 705.300 282.790 ;
        RECT 719.830 282.725 722.400 282.760 ;
        RECT 737.050 282.725 739.310 282.790 ;
        RECT 679.060 282.710 686.360 282.715 ;
        RECT 679.060 280.115 687.310 282.710 ;
        RECT 696.340 280.125 705.300 282.725 ;
        RECT 714.110 280.125 722.400 282.725 ;
        RECT 731.350 280.125 739.310 282.725 ;
        RECT 748.830 282.730 754.770 282.735 ;
        RECT 748.830 280.140 756.030 282.730 ;
        RECT 799.200 281.335 801.300 283.935 ;
        RECT 819.020 280.995 824.960 283.595 ;
        RECT 830.910 283.505 833.660 283.510 ;
        RECT 838.120 283.505 840.870 283.510 ;
        RECT 843.970 283.505 846.630 283.510 ;
        RECT 827.630 283.500 851.910 283.505 ;
        RECT 827.630 280.905 852.840 283.500 ;
        RECT 859.610 283.225 864.950 285.220 ;
        RECT 859.610 283.220 861.190 283.225 ;
        RECT 859.610 282.390 860.810 283.220 ;
        RECT 859.500 282.385 860.810 282.390 ;
        RECT 830.910 280.900 833.660 280.905 ;
        RECT 838.120 280.900 840.870 280.905 ;
        RECT 843.970 280.900 846.630 280.905 ;
        RECT 851.650 280.870 852.840 280.905 ;
        RECT 855.600 281.220 860.810 282.385 ;
        RECT 748.830 280.135 754.770 280.140 ;
        RECT 684.660 280.100 687.310 280.115 ;
        RECT 685.020 280.080 687.310 280.100 ;
        RECT 702.000 280.070 705.300 280.125 ;
        RECT 719.830 280.050 722.400 280.125 ;
        RECT 737.050 280.090 739.310 280.125 ;
        RECT 855.600 279.785 859.620 281.220 ;
        RECT 594.760 272.775 596.860 275.375 ;
        RECT 600.150 272.790 631.070 278.840 ;
        RECT 749.250 277.230 755.190 277.265 ;
        RECT 749.250 277.225 757.210 277.230 ;
        RECT 714.270 277.140 720.210 277.175 ;
        RECT 731.440 277.170 737.380 277.205 ;
        RECT 731.440 277.165 739.400 277.170 ;
        RECT 714.270 277.135 722.220 277.140 ;
        RECT 679.470 277.020 685.410 277.055 ;
        RECT 696.700 277.040 702.640 277.075 ;
        RECT 696.700 277.035 704.660 277.040 ;
        RECT 679.470 277.015 687.410 277.020 ;
        RECT 634.650 273.225 636.750 275.825 ;
        RECT 638.840 273.315 640.940 275.915 ;
        RECT 644.960 275.895 646.320 275.900 ;
        RECT 642.940 273.300 646.320 275.895 ;
        RECT 679.470 274.455 692.650 277.015 ;
        RECT 696.700 274.475 709.880 277.035 ;
        RECT 714.270 274.575 727.450 277.135 ;
        RECT 731.440 274.605 744.620 277.165 ;
        RECT 749.250 274.665 762.430 277.225 ;
        RECT 789.030 275.895 792.990 277.530 ;
        RECT 796.420 275.895 799.870 275.900 ;
        RECT 754.480 274.650 762.430 274.665 ;
        RECT 756.490 274.625 762.430 274.650 ;
        RECT 780.630 275.885 799.870 275.895 ;
        RECT 780.630 275.860 815.540 275.885 ;
        RECT 780.630 275.855 818.690 275.860 ;
        RECT 780.630 275.850 834.390 275.855 ;
        RECT 838.090 275.850 842.590 275.895 ;
        RECT 736.660 274.600 744.620 274.605 ;
        RECT 719.510 274.570 727.450 274.575 ;
        RECT 721.510 274.535 727.450 274.570 ;
        RECT 738.680 274.565 744.620 274.600 ;
        RECT 780.630 274.540 842.590 275.850 ;
        RECT 701.930 274.460 709.880 274.475 ;
        RECT 684.710 274.450 692.650 274.455 ;
        RECT 686.710 274.415 692.650 274.450 ;
        RECT 703.940 274.435 709.880 274.460 ;
        RECT 780.630 274.530 844.600 274.540 ;
        RECT 780.630 273.635 845.230 274.530 ;
        RECT 855.600 274.510 859.620 275.845 ;
        RECT 855.600 274.480 862.520 274.510 ;
        RECT 847.750 273.645 850.370 273.650 ;
        RECT 847.750 273.635 851.850 273.645 ;
        RECT 642.940 273.295 645.040 273.300 ;
        RECT 780.630 273.295 851.850 273.635 ;
        RECT 796.420 273.285 838.450 273.295 ;
        RECT 842.350 273.290 851.850 273.295 ;
        RECT 796.420 273.260 799.870 273.285 ;
        RECT 815.300 273.260 838.450 273.285 ;
        RECT 815.300 273.255 834.390 273.260 ;
        RECT 815.300 273.240 818.690 273.255 ;
        RECT 600.130 271.820 631.070 272.790 ;
        RECT 600.130 266.540 604.600 271.820 ;
        RECT 626.610 270.410 631.070 271.820 ;
        RECT 758.360 271.615 761.060 271.620 ;
        RECT 758.360 271.595 764.400 271.615 ;
        RECT 755.030 271.590 764.400 271.595 ;
        RECT 753.010 271.585 764.400 271.590 ;
        RECT 740.560 271.555 743.250 271.560 ;
        RECT 740.560 271.535 746.590 271.555 ;
        RECT 737.220 271.530 746.590 271.535 ;
        RECT 735.200 271.525 746.590 271.530 ;
        RECT 725.400 271.520 729.420 271.525 ;
        RECT 718.030 271.505 720.420 271.510 ;
        RECT 723.370 271.505 729.420 271.520 ;
        RECT 718.030 271.495 729.420 271.505 ;
        RECT 707.830 271.420 711.850 271.425 ;
        RECT 700.470 271.405 702.850 271.410 ;
        RECT 705.800 271.405 711.850 271.420 ;
        RECT 690.600 271.400 694.620 271.405 ;
        RECT 683.250 271.385 685.620 271.390 ;
        RECT 688.580 271.385 694.620 271.400 ;
        RECT 700.470 271.395 711.850 271.405 ;
        RECT 683.250 271.375 694.620 271.385 ;
        RECT 626.610 267.160 631.180 270.410 ;
        RECT 679.590 268.805 694.620 271.375 ;
        RECT 696.820 268.825 711.850 271.395 ;
        RECT 714.390 268.925 729.420 271.495 ;
        RECT 731.560 268.955 746.590 271.525 ;
        RECT 749.370 269.015 764.400 271.585 ;
        RECT 844.340 271.045 851.850 273.290 ;
        RECT 855.600 273.245 862.530 274.480 ;
        RECT 859.640 272.455 862.530 273.245 ;
        RECT 844.340 271.035 850.370 271.045 ;
        RECT 847.750 271.020 850.370 271.035 ;
        RECT 749.370 268.995 761.060 269.015 ;
        RECT 749.370 268.990 755.420 268.995 ;
        RECT 749.370 268.985 753.390 268.990 ;
        RECT 758.360 268.980 761.060 268.995 ;
        RECT 731.560 268.940 743.250 268.955 ;
        RECT 731.560 268.935 741.240 268.940 ;
        RECT 731.560 268.925 737.580 268.935 ;
        RECT 714.390 268.905 726.110 268.925 ;
        RECT 735.200 268.920 737.580 268.925 ;
        RECT 714.390 268.895 720.420 268.905 ;
        RECT 723.370 268.900 726.110 268.905 ;
        RECT 718.030 268.880 720.420 268.895 ;
        RECT 696.820 268.805 708.530 268.825 ;
        RECT 679.590 268.785 691.280 268.805 ;
        RECT 696.820 268.795 702.850 268.805 ;
        RECT 705.800 268.800 708.530 268.805 ;
        RECT 700.470 268.790 702.850 268.795 ;
        RECT 679.590 268.775 685.620 268.785 ;
        RECT 688.580 268.780 691.280 268.785 ;
        RECT 683.250 268.770 685.620 268.775 ;
        RECT 799.170 268.390 815.190 268.395 ;
        RECT 780.640 268.320 796.660 268.335 ;
        RECT 799.170 268.320 816.160 268.390 ;
        RECT 626.610 266.590 631.070 267.160 ;
        RECT 780.640 265.795 816.160 268.320 ;
        RECT 838.100 267.735 842.120 270.335 ;
        RECT 859.640 269.855 864.940 272.455 ;
        RECT 859.640 269.850 861.240 269.855 ;
        RECT 859.640 269.175 860.570 269.850 ;
        RECT 855.680 267.980 860.570 269.175 ;
        RECT 855.680 266.575 859.700 267.980 ;
        RECT 780.640 265.740 798.380 265.795 ;
        RECT 815.010 265.760 816.160 265.795 ;
        RECT 780.640 265.735 796.660 265.740 ;
        RECT 684.860 261.185 686.370 261.200 ;
        RECT 702.050 261.195 703.430 261.220 ;
        RECT 719.760 261.195 721.190 261.200 ;
        RECT 737.090 261.195 738.410 261.200 ;
        RECT 594.610 255.045 596.710 257.645 ;
        RECT 600.000 255.060 630.920 261.110 ;
        RECT 679.040 258.585 686.370 261.185 ;
        RECT 696.320 258.595 703.430 261.195 ;
        RECT 714.090 258.595 721.190 261.195 ;
        RECT 731.330 258.595 738.410 261.195 ;
        RECT 748.810 261.180 754.750 261.205 ;
        RECT 748.810 258.605 756.310 261.180 ;
        RECT 684.860 258.570 686.370 258.585 ;
        RECT 702.050 258.560 703.430 258.595 ;
        RECT 719.760 258.570 721.190 258.595 ;
        RECT 737.090 258.570 738.410 258.595 ;
        RECT 754.480 258.580 756.310 258.605 ;
        RECT 855.550 259.500 859.570 259.865 ;
        RECT 855.550 259.490 861.590 259.500 ;
        RECT 634.500 255.495 636.600 258.095 ;
        RECT 638.690 255.585 640.790 258.185 ;
        RECT 644.780 258.165 646.140 258.200 ;
        RECT 642.790 255.600 646.140 258.165 ;
        RECT 855.550 257.375 861.720 259.490 ;
        RECT 855.550 257.265 864.880 257.375 ;
        RECT 749.230 255.700 755.170 255.735 ;
        RECT 749.230 255.695 757.190 255.700 ;
        RECT 731.420 255.670 737.360 255.675 ;
        RECT 714.250 255.610 720.190 255.645 ;
        RECT 731.420 255.635 739.370 255.670 ;
        RECT 714.250 255.605 722.190 255.610 ;
        RECT 642.790 255.565 644.890 255.600 ;
        RECT 679.450 255.500 685.390 255.525 ;
        RECT 696.680 255.510 702.620 255.545 ;
        RECT 696.680 255.505 704.630 255.510 ;
        RECT 352.790 254.120 411.130 254.470 ;
        RECT 352.790 248.420 411.110 254.120 ;
        RECT 599.980 254.090 630.920 255.060 ;
        RECT 599.980 248.810 604.450 254.090 ;
        RECT 626.460 252.680 630.920 254.090 ;
        RECT 679.450 255.485 687.400 255.500 ;
        RECT 679.450 252.925 692.630 255.485 ;
        RECT 696.680 252.945 709.860 255.505 ;
        RECT 714.250 253.045 727.430 255.605 ;
        RECT 731.420 253.075 744.600 255.635 ;
        RECT 749.230 253.135 762.410 255.695 ;
        RECT 860.000 254.775 864.880 257.265 ;
        RECT 860.000 254.760 860.990 254.775 ;
        RECT 860.000 254.100 860.850 254.760 ;
        RECT 859.520 254.095 860.850 254.100 ;
        RECT 754.470 253.130 762.410 253.135 ;
        RECT 756.470 253.095 762.410 253.130 ;
        RECT 855.610 253.250 860.850 254.095 ;
        RECT 736.650 253.070 744.600 253.075 ;
        RECT 719.480 253.030 727.430 253.045 ;
        RECT 738.660 253.035 744.600 253.070 ;
        RECT 721.490 253.005 727.430 253.030 ;
        RECT 701.920 252.940 709.860 252.945 ;
        RECT 684.700 252.920 692.630 252.925 ;
        RECT 686.690 252.885 692.630 252.920 ;
        RECT 703.920 252.905 709.860 252.940 ;
        RECT 626.460 249.430 631.030 252.680 ;
        RECT 855.610 251.495 859.630 253.250 ;
        RECT 758.340 250.085 761.040 250.100 ;
        RECT 752.980 250.065 755.370 250.070 ;
        RECT 758.340 250.065 764.380 250.085 ;
        RECT 752.980 250.055 764.380 250.065 ;
        RECT 740.530 250.025 743.240 250.040 ;
        RECT 723.360 249.995 726.040 250.010 ;
        RECT 735.200 250.005 737.590 250.010 ;
        RECT 740.530 250.005 746.570 250.025 ;
        RECT 735.200 249.995 746.570 250.005 ;
        RECT 723.360 249.975 729.400 249.995 ;
        RECT 720.030 249.970 729.400 249.975 ;
        RECT 718.000 249.965 729.400 249.970 ;
        RECT 705.790 249.895 708.490 249.900 ;
        RECT 688.550 249.875 691.270 249.890 ;
        RECT 700.440 249.875 702.850 249.880 ;
        RECT 705.790 249.875 711.830 249.895 ;
        RECT 688.550 249.855 694.600 249.875 ;
        RECT 700.440 249.865 711.830 249.875 ;
        RECT 685.230 249.850 694.600 249.855 ;
        RECT 683.200 249.845 694.600 249.850 ;
        RECT 626.460 248.860 630.920 249.430 ;
        RECT 679.570 247.275 694.600 249.845 ;
        RECT 696.800 247.295 711.830 249.865 ;
        RECT 714.370 247.395 729.400 249.965 ;
        RECT 731.540 247.425 746.570 249.995 ;
        RECT 749.350 247.485 764.380 250.055 ;
        RECT 749.350 247.465 761.040 247.485 ;
        RECT 749.350 247.455 755.370 247.465 ;
        RECT 752.980 247.450 755.370 247.455 ;
        RECT 758.340 247.450 761.040 247.465 ;
        RECT 731.540 247.405 743.240 247.425 ;
        RECT 731.540 247.395 737.590 247.405 ;
        RECT 740.530 247.400 743.240 247.405 ;
        RECT 714.370 247.380 726.040 247.395 ;
        RECT 735.200 247.390 737.590 247.395 ;
        RECT 714.370 247.375 724.050 247.380 ;
        RECT 714.370 247.365 720.430 247.375 ;
        RECT 718.000 247.360 720.430 247.365 ;
        RECT 696.800 247.275 708.490 247.295 ;
        RECT 679.570 247.260 691.270 247.275 ;
        RECT 696.800 247.265 702.850 247.275 ;
        RECT 700.440 247.260 702.850 247.265 ;
        RECT 705.790 247.260 708.490 247.275 ;
        RECT 679.570 247.255 689.250 247.260 ;
        RECT 679.570 247.245 685.620 247.255 ;
        RECT 683.200 247.240 685.620 247.245 ;
        RECT -53.360 217.565 -25.270 225.185 ;
        RECT -53.400 129.915 -25.310 137.535 ;
        RECT -53.280 10.475 -25.190 18.095 ;
      LAYER li1 ;
        RECT 362.820 371.640 364.540 372.690 ;
        RECT 401.570 371.830 404.570 373.040 ;
        RECT 363.140 371.050 363.770 371.640 ;
        RECT 369.770 371.050 370.150 371.070 ;
        RECT 356.640 371.030 370.150 371.050 ;
        RECT 356.620 370.540 370.150 371.030 ;
        RECT 401.730 371.020 402.220 371.060 ;
        RECT 402.570 371.020 403.240 371.830 ;
        RECT 408.340 371.020 408.720 371.040 ;
        RECT 395.210 371.000 408.720 371.020 ;
        RECT 382.480 370.950 382.970 370.990 ;
        RECT 389.090 370.950 389.470 370.970 ;
        RECT 375.960 370.930 389.470 370.950 ;
        RECT 356.620 369.350 356.890 370.540 ;
        RECT 363.140 370.530 363.770 370.540 ;
        RECT 359.980 369.630 360.150 370.280 ;
        RECT 363.160 369.950 363.650 370.530 ;
        RECT 366.380 369.970 367.000 370.540 ;
        RECT 213.770 366.830 227.000 368.840 ;
        RECT 233.810 366.820 247.040 368.830 ;
        RECT 253.870 366.820 267.100 368.830 ;
        RECT 273.920 366.820 287.150 368.830 ;
        RECT 356.480 366.370 356.940 369.350 ;
        RECT 359.840 368.950 360.230 369.630 ;
        RECT 363.270 369.260 363.440 369.950 ;
        RECT 366.560 369.580 366.730 369.970 ;
        RECT 369.770 369.820 370.150 370.540 ;
        RECT 375.940 370.440 389.470 370.930 ;
        RECT 366.430 369.480 366.820 369.580 ;
        RECT 366.310 369.410 366.820 369.480 ;
        RECT 366.310 368.960 366.840 369.410 ;
        RECT 369.850 369.260 370.020 369.820 ;
        RECT 375.940 369.250 376.210 370.440 ;
        RECT 382.480 369.850 382.970 370.440 ;
        RECT 365.740 368.950 366.840 368.960 ;
        RECT 359.840 368.570 366.840 368.950 ;
        RECT 359.840 368.560 365.820 368.570 ;
        RECT 359.900 368.550 365.820 368.560 ;
        RECT 366.440 368.530 366.840 368.570 ;
        RECT 369.660 366.410 370.550 366.460 ;
        RECT 369.620 366.370 370.550 366.410 ;
        RECT 226.430 366.220 227.750 366.290 ;
        RECT 246.470 366.220 247.790 366.280 ;
        RECT 266.530 366.220 267.850 366.280 ;
        RECT 286.580 366.220 287.900 366.280 ;
        RECT 212.340 366.140 287.900 366.220 ;
        RECT 356.460 366.160 370.550 366.370 ;
        RECT 375.800 366.270 376.260 369.250 ;
        RECT 382.590 369.160 382.760 369.850 ;
        RECT 389.090 369.720 389.470 370.440 ;
        RECT 395.190 370.510 408.720 371.000 ;
        RECT 389.170 369.160 389.340 369.720 ;
        RECT 395.190 369.320 395.460 370.510 ;
        RECT 398.550 369.600 398.720 370.250 ;
        RECT 401.730 369.920 402.220 370.510 ;
        RECT 402.570 370.480 403.240 370.510 ;
        RECT 388.980 366.310 389.870 366.360 ;
        RECT 395.050 366.340 395.510 369.320 ;
        RECT 398.410 368.920 398.800 369.600 ;
        RECT 401.840 369.230 402.010 369.920 ;
        RECT 404.980 369.880 405.450 370.510 ;
        RECT 405.130 369.550 405.300 369.880 ;
        RECT 408.340 369.790 408.720 370.510 ;
        RECT 405.000 369.450 405.390 369.550 ;
        RECT 404.880 369.380 405.390 369.450 ;
        RECT 404.880 368.930 405.410 369.380 ;
        RECT 408.420 369.230 408.590 369.790 ;
        RECT 404.310 368.920 405.410 368.930 ;
        RECT 398.410 368.540 405.410 368.920 ;
        RECT 398.410 368.530 404.390 368.540 ;
        RECT 398.470 368.520 404.390 368.530 ;
        RECT 405.010 368.500 405.410 368.540 ;
        RECT 408.230 366.380 409.120 366.430 ;
        RECT 408.190 366.340 409.120 366.380 ;
        RECT 388.940 366.270 389.870 366.310 ;
        RECT 211.970 365.970 287.900 366.140 ;
        RECT 212.340 365.960 287.900 365.970 ;
        RECT 212.420 365.930 227.750 365.960 ;
        RECT 226.430 365.910 227.750 365.930 ;
        RECT 232.460 365.920 247.790 365.960 ;
        RECT 252.520 365.920 267.850 365.960 ;
        RECT 272.570 365.920 287.900 365.960 ;
        RECT 211.160 362.910 212.590 362.980 ;
        RECT 211.160 362.850 226.840 362.910 ;
        RECT 211.160 362.680 226.870 362.850 ;
        RECT 211.160 362.640 226.840 362.680 ;
        RECT 211.160 362.600 212.590 362.640 ;
        RECT -44.590 358.325 -34.360 359.630 ;
        RECT -46.100 358.155 -32.770 358.325 ;
        RECT -44.590 357.990 -34.360 358.155 ;
        RECT -44.045 357.650 -43.865 357.990 ;
        RECT -51.735 357.630 -27.285 357.650 ;
        RECT -51.980 357.470 -26.890 357.630 ;
        RECT -51.980 357.460 -51.400 357.470 ;
        RECT -50.690 357.460 -50.110 357.470 ;
        RECT -49.400 357.460 -48.820 357.470 ;
        RECT -48.110 357.460 -47.530 357.470 ;
        RECT -46.820 357.460 -46.240 357.470 ;
        RECT -45.530 357.460 -44.950 357.470 ;
        RECT -44.240 357.460 -43.660 357.470 ;
        RECT -42.950 357.460 -42.370 357.470 ;
        RECT -41.660 357.460 -41.080 357.470 ;
        RECT -40.370 357.460 -39.790 357.470 ;
        RECT -39.080 357.460 -38.500 357.470 ;
        RECT -37.790 357.460 -37.210 357.470 ;
        RECT -36.500 357.460 -35.920 357.470 ;
        RECT -35.210 357.460 -34.630 357.470 ;
        RECT -33.920 357.460 -33.340 357.470 ;
        RECT -32.630 357.460 -32.050 357.470 ;
        RECT -31.340 357.460 -30.760 357.470 ;
        RECT -30.050 357.460 -29.470 357.470 ;
        RECT -28.760 357.460 -28.180 357.470 ;
        RECT -27.470 357.460 -26.890 357.470 ;
        RECT -53.090 353.355 -52.920 356.455 ;
        RECT -52.420 353.915 -52.250 355.535 ;
        RECT -49.840 353.915 -49.670 355.535 ;
        RECT -47.260 353.915 -47.090 355.535 ;
        RECT -44.680 353.915 -44.510 355.535 ;
        RECT -42.100 353.915 -41.930 355.535 ;
        RECT -39.520 353.915 -39.350 355.535 ;
        RECT -36.940 353.915 -36.770 355.535 ;
        RECT -34.360 353.915 -34.190 355.535 ;
        RECT -31.780 353.915 -31.610 355.535 ;
        RECT -29.200 353.915 -29.030 355.535 ;
        RECT -26.620 353.915 -26.450 355.535 ;
        RECT -25.950 353.355 -25.780 356.455 ;
        RECT 211.160 356.370 211.570 362.600 ;
        RECT 227.360 359.650 227.630 365.910 ;
        RECT 246.470 365.900 247.790 365.920 ;
        RECT 266.530 365.900 267.850 365.920 ;
        RECT 286.580 365.900 287.900 365.920 ;
        RECT 231.200 362.900 232.630 362.970 ;
        RECT 231.200 362.840 246.880 362.900 ;
        RECT 231.200 362.670 246.910 362.840 ;
        RECT 231.200 362.630 246.880 362.670 ;
        RECT 231.200 362.590 232.630 362.630 ;
        RECT 226.610 359.620 227.930 359.650 ;
        RECT 212.660 359.560 227.930 359.620 ;
        RECT 211.970 359.390 227.930 359.560 ;
        RECT 212.660 359.350 227.930 359.390 ;
        RECT 226.610 359.270 227.930 359.350 ;
        RECT 211.140 356.330 212.740 356.370 ;
        RECT 211.140 356.060 226.880 356.330 ;
        RECT 211.140 355.990 212.740 356.060 ;
        RECT -46.100 351.485 -32.770 351.655 ;
        RECT 211.160 349.870 211.570 355.990 ;
        RECT 227.360 353.080 227.630 359.270 ;
        RECT 231.200 356.360 231.610 362.590 ;
        RECT 247.400 359.640 247.670 365.900 ;
        RECT 251.260 362.900 252.690 362.970 ;
        RECT 251.260 362.840 266.940 362.900 ;
        RECT 251.260 362.670 266.970 362.840 ;
        RECT 251.260 362.630 266.940 362.670 ;
        RECT 251.260 362.590 252.690 362.630 ;
        RECT 246.650 359.610 247.970 359.640 ;
        RECT 232.700 359.550 247.970 359.610 ;
        RECT 232.010 359.380 247.970 359.550 ;
        RECT 232.700 359.340 247.970 359.380 ;
        RECT 246.650 359.260 247.970 359.340 ;
        RECT 231.180 356.320 232.780 356.360 ;
        RECT 231.180 356.050 246.920 356.320 ;
        RECT 231.180 355.980 232.780 356.050 ;
        RECT 226.460 353.010 227.780 353.080 ;
        RECT 212.650 352.980 227.780 353.010 ;
        RECT 211.970 352.810 227.780 352.980 ;
        RECT 212.650 352.740 227.780 352.810 ;
        RECT 226.460 352.700 227.780 352.740 ;
        RECT 227.360 352.690 227.630 352.700 ;
        RECT 211.070 349.840 211.570 349.870 ;
        RECT 211.070 349.790 212.640 349.840 ;
        RECT 231.200 349.830 231.610 355.980 ;
        RECT 247.400 353.070 247.670 359.260 ;
        RECT 251.260 356.360 251.670 362.590 ;
        RECT 267.460 359.640 267.730 365.900 ;
        RECT 271.310 362.900 272.740 362.970 ;
        RECT 271.310 362.840 286.990 362.900 ;
        RECT 271.310 362.670 287.020 362.840 ;
        RECT 271.310 362.630 286.990 362.670 ;
        RECT 271.310 362.590 272.740 362.630 ;
        RECT 266.710 359.610 268.030 359.640 ;
        RECT 252.760 359.550 268.030 359.610 ;
        RECT 252.070 359.380 268.030 359.550 ;
        RECT 252.760 359.340 268.030 359.380 ;
        RECT 266.710 359.260 268.030 359.340 ;
        RECT 251.240 356.320 252.840 356.360 ;
        RECT 251.240 356.050 266.980 356.320 ;
        RECT 251.240 355.980 252.840 356.050 ;
        RECT 246.500 353.000 247.820 353.070 ;
        RECT 232.690 352.970 247.820 353.000 ;
        RECT 232.010 352.800 247.820 352.970 ;
        RECT 232.690 352.730 247.820 352.800 ;
        RECT 246.500 352.690 247.820 352.730 ;
        RECT 247.400 352.680 247.670 352.690 ;
        RECT 251.260 349.830 251.670 355.980 ;
        RECT 267.460 353.070 267.730 359.260 ;
        RECT 271.310 356.360 271.720 362.590 ;
        RECT 287.510 359.640 287.780 365.900 ;
        RECT 355.060 363.620 356.140 365.630 ;
        RECT 356.480 363.620 356.760 366.160 ;
        RECT 359.840 365.550 360.010 365.710 ;
        RECT 355.060 363.150 356.760 363.620 ;
        RECT 286.760 359.610 288.080 359.640 ;
        RECT 272.810 359.550 288.080 359.610 ;
        RECT 272.120 359.380 288.080 359.550 ;
        RECT 272.810 359.340 288.080 359.380 ;
        RECT 286.760 359.260 288.080 359.340 ;
        RECT 271.290 356.320 272.890 356.360 ;
        RECT 271.290 356.050 287.030 356.320 ;
        RECT 271.290 355.980 272.890 356.050 ;
        RECT 266.560 353.000 267.880 353.070 ;
        RECT 252.750 352.970 267.880 353.000 ;
        RECT 252.070 352.800 267.880 352.970 ;
        RECT 252.750 352.730 267.880 352.800 ;
        RECT 266.560 352.690 267.880 352.730 ;
        RECT 267.460 352.680 267.730 352.690 ;
        RECT 271.310 349.830 271.720 355.980 ;
        RECT 287.510 353.070 287.780 359.260 ;
        RECT 286.610 353.000 287.930 353.070 ;
        RECT 272.800 352.970 287.930 353.000 ;
        RECT 272.120 352.800 287.930 352.970 ;
        RECT 272.800 352.730 287.930 352.800 ;
        RECT 286.610 352.690 287.930 352.730 ;
        RECT 231.180 349.790 232.680 349.830 ;
        RECT 251.240 349.790 252.740 349.830 ;
        RECT 271.290 349.790 272.790 349.830 ;
        RECT 211.070 349.730 286.370 349.790 ;
        RECT 211.070 349.680 287.000 349.730 ;
        RECT 211.070 349.530 287.020 349.680 ;
        RECT 211.070 349.520 226.870 349.530 ;
        RECT 211.070 349.470 226.850 349.520 ;
        RECT 231.180 349.510 246.910 349.530 ;
        RECT 251.240 349.510 266.970 349.530 ;
        RECT 271.290 349.510 287.020 349.530 ;
        RECT 211.070 349.460 212.550 349.470 ;
        RECT 231.180 349.460 246.890 349.510 ;
        RECT 251.240 349.460 266.950 349.510 ;
        RECT 271.290 349.460 287.000 349.510 ;
        RECT 211.070 349.450 211.570 349.460 ;
        RECT 231.180 349.450 232.590 349.460 ;
        RECT 251.240 349.450 252.650 349.460 ;
        RECT 271.290 349.450 272.700 349.460 ;
        RECT 211.070 341.990 211.480 349.450 ;
        RECT 231.200 349.440 231.610 349.450 ;
        RECT 251.260 349.440 251.670 349.450 ;
        RECT 271.310 349.440 271.720 349.450 ;
        RECT 287.490 348.240 287.920 352.690 ;
        RECT 355.060 351.330 356.140 363.150 ;
        RECT 356.480 351.510 356.760 363.150 ;
        RECT 359.790 351.550 360.070 365.550 ;
        RECT 363.070 365.530 363.350 366.160 ;
        RECT 369.620 366.110 370.550 366.160 ;
        RECT 356.420 351.390 356.760 351.510 ;
        RECT 288.460 348.240 289.350 348.760 ;
        RECT 213.730 345.840 226.960 347.850 ;
        RECT 233.700 345.840 246.930 347.850 ;
        RECT 253.810 345.840 267.040 347.850 ;
        RECT 273.920 345.840 287.150 347.850 ;
        RECT 287.490 347.570 289.350 348.240 ;
        RECT 287.490 345.300 287.920 347.570 ;
        RECT 288.460 347.040 289.350 347.570 ;
        RECT 356.420 347.490 356.750 351.390 ;
        RECT 359.740 351.330 360.070 351.550 ;
        RECT 363.060 365.370 363.350 365.530 ;
        RECT 359.740 350.340 360.040 351.330 ;
        RECT 363.060 351.310 363.340 365.370 ;
        RECT 366.420 365.320 366.590 365.710 ;
        RECT 366.360 351.540 366.640 365.320 ;
        RECT 369.620 365.220 370.000 366.110 ;
        RECT 375.780 366.060 389.870 366.270 ;
        RECT 395.030 366.130 409.120 366.340 ;
        RECT 363.130 350.810 363.300 351.310 ;
        RECT 366.360 351.100 366.680 351.540 ;
        RECT 369.630 351.120 369.910 365.220 ;
        RECT 374.380 351.230 375.460 365.530 ;
        RECT 375.800 351.410 376.080 366.060 ;
        RECT 382.390 365.430 382.670 366.060 ;
        RECT 375.740 351.290 376.080 351.410 ;
        RECT 382.380 365.270 382.670 365.430 ;
        RECT 388.940 366.010 389.870 366.060 ;
        RECT 366.380 350.360 366.680 351.100 ;
        RECT 369.710 350.810 369.880 351.120 ;
        RECT 366.380 350.340 367.170 350.360 ;
        RECT 359.740 350.030 367.170 350.340 ;
        RECT 359.740 350.000 360.040 350.030 ;
        RECT 366.290 350.010 366.680 350.030 ;
        RECT 366.380 349.990 366.680 350.010 ;
        RECT 369.640 347.530 370.530 347.580 ;
        RECT 369.600 347.490 370.530 347.530 ;
        RECT 356.420 347.280 370.530 347.490 ;
        RECT 356.420 347.200 356.750 347.280 ;
        RECT 226.390 345.210 227.710 345.300 ;
        RECT 246.360 345.210 247.680 345.300 ;
        RECT 266.470 345.210 267.790 345.300 ;
        RECT 286.580 345.210 287.920 345.300 ;
        RECT 212.380 345.150 287.920 345.210 ;
        RECT 211.930 344.980 287.920 345.150 ;
        RECT 212.380 344.960 287.920 344.980 ;
        RECT 212.380 344.950 287.900 344.960 ;
        RECT 212.380 344.940 227.710 344.950 ;
        RECT 232.350 344.940 247.680 344.950 ;
        RECT 252.460 344.940 267.790 344.950 ;
        RECT 272.570 344.940 287.900 344.950 ;
        RECT 226.390 344.920 227.710 344.940 ;
        RECT 246.360 344.920 247.680 344.940 ;
        RECT 266.470 344.920 267.790 344.940 ;
        RECT 286.580 344.920 287.900 344.940 ;
        RECT 211.070 341.920 212.550 341.990 ;
        RECT 211.070 341.860 226.800 341.920 ;
        RECT 211.070 341.690 226.830 341.860 ;
        RECT 211.070 341.650 226.800 341.690 ;
        RECT 211.070 341.610 212.550 341.650 ;
        RECT 211.070 341.110 211.530 341.610 ;
        RECT 211.120 335.380 211.530 341.110 ;
        RECT 227.320 338.660 227.590 344.920 ;
        RECT 231.090 341.920 232.520 341.990 ;
        RECT 231.090 341.860 246.770 341.920 ;
        RECT 231.090 341.690 246.800 341.860 ;
        RECT 231.090 341.650 246.770 341.690 ;
        RECT 231.090 341.610 232.520 341.650 ;
        RECT 226.570 338.630 227.890 338.660 ;
        RECT 212.620 338.570 227.890 338.630 ;
        RECT 211.930 338.400 227.890 338.570 ;
        RECT 212.620 338.360 227.890 338.400 ;
        RECT 226.570 338.280 227.890 338.360 ;
        RECT 211.100 335.340 212.700 335.380 ;
        RECT 211.100 335.070 226.840 335.340 ;
        RECT 211.100 335.000 212.700 335.070 ;
        RECT 4.860 328.790 13.020 329.810 ;
        RECT 18.200 328.770 26.360 329.790 ;
        RECT 31.570 328.800 39.730 329.820 ;
        RECT 44.800 328.800 52.960 329.820 ;
        RECT 58.070 328.770 66.230 329.790 ;
        RECT 71.340 328.800 79.500 329.820 ;
        RECT 84.470 328.820 92.630 329.840 ;
        RECT 96.960 328.620 103.140 329.970 ;
        RECT 211.120 328.850 211.530 335.000 ;
        RECT 227.320 332.090 227.590 338.280 ;
        RECT 231.090 335.380 231.500 341.610 ;
        RECT 247.290 338.660 247.560 344.920 ;
        RECT 251.200 341.920 252.630 341.990 ;
        RECT 251.200 341.860 266.880 341.920 ;
        RECT 251.200 341.690 266.910 341.860 ;
        RECT 251.200 341.650 266.880 341.690 ;
        RECT 251.200 341.610 252.630 341.650 ;
        RECT 246.540 338.630 247.860 338.660 ;
        RECT 232.590 338.570 247.860 338.630 ;
        RECT 231.900 338.400 247.860 338.570 ;
        RECT 232.590 338.360 247.860 338.400 ;
        RECT 246.540 338.280 247.860 338.360 ;
        RECT 231.070 335.340 232.670 335.380 ;
        RECT 231.070 335.070 246.810 335.340 ;
        RECT 231.070 335.000 232.670 335.070 ;
        RECT 226.420 332.020 227.740 332.090 ;
        RECT 212.610 331.990 227.740 332.020 ;
        RECT 211.930 331.820 227.740 331.990 ;
        RECT 212.610 331.750 227.740 331.820 ;
        RECT 226.420 331.710 227.740 331.750 ;
        RECT 227.320 331.700 227.590 331.710 ;
        RECT 231.090 328.850 231.500 335.000 ;
        RECT 247.290 332.090 247.560 338.280 ;
        RECT 251.200 335.380 251.610 341.610 ;
        RECT 267.400 338.660 267.670 344.920 ;
        RECT 287.310 344.210 287.780 344.920 ;
        RECT 271.310 341.920 272.740 341.990 ;
        RECT 271.310 341.860 286.990 341.920 ;
        RECT 271.310 341.690 287.020 341.860 ;
        RECT 271.310 341.650 286.990 341.690 ;
        RECT 271.310 341.610 272.740 341.650 ;
        RECT 266.650 338.630 267.970 338.660 ;
        RECT 252.700 338.570 267.970 338.630 ;
        RECT 252.010 338.400 267.970 338.570 ;
        RECT 252.700 338.360 267.970 338.400 ;
        RECT 266.650 338.280 267.970 338.360 ;
        RECT 251.180 335.340 252.780 335.380 ;
        RECT 251.180 335.070 266.920 335.340 ;
        RECT 251.180 335.000 252.780 335.070 ;
        RECT 246.390 332.020 247.710 332.090 ;
        RECT 232.580 331.990 247.710 332.020 ;
        RECT 231.900 331.820 247.710 331.990 ;
        RECT 232.580 331.750 247.710 331.820 ;
        RECT 246.390 331.710 247.710 331.750 ;
        RECT 247.290 331.700 247.560 331.710 ;
        RECT 251.200 328.850 251.610 335.000 ;
        RECT 267.400 332.090 267.670 338.280 ;
        RECT 271.310 335.380 271.720 341.610 ;
        RECT 287.510 338.660 287.780 344.210 ;
        RECT 286.760 338.630 288.080 338.660 ;
        RECT 272.810 338.570 288.080 338.630 ;
        RECT 272.120 338.400 288.080 338.570 ;
        RECT 272.810 338.360 288.080 338.400 ;
        RECT 286.760 338.280 288.080 338.360 ;
        RECT 271.290 335.340 272.890 335.380 ;
        RECT 271.290 335.070 287.030 335.340 ;
        RECT 271.290 335.000 272.890 335.070 ;
        RECT 266.500 332.020 267.820 332.090 ;
        RECT 252.690 331.990 267.820 332.020 ;
        RECT 252.010 331.820 267.820 331.990 ;
        RECT 252.690 331.750 267.820 331.820 ;
        RECT 266.500 331.710 267.820 331.750 ;
        RECT 267.400 331.700 267.670 331.710 ;
        RECT 271.310 328.850 271.720 335.000 ;
        RECT 287.510 332.090 287.780 338.280 ;
        RECT 355.040 332.450 356.120 346.750 ;
        RECT 356.460 332.810 356.740 347.200 ;
        RECT 359.820 346.670 359.990 346.830 ;
        RECT 286.610 332.040 287.930 332.090 ;
        RECT 286.610 332.020 288.020 332.040 ;
        RECT 272.800 331.990 288.020 332.020 ;
        RECT 272.120 331.820 288.020 331.990 ;
        RECT 272.800 331.750 288.020 331.820 ;
        RECT 286.610 331.710 288.020 331.750 ;
        RECT 211.100 328.790 212.600 328.850 ;
        RECT 231.070 328.790 232.570 328.850 ;
        RECT 251.180 328.790 252.680 328.850 ;
        RECT 271.290 328.790 272.790 328.850 ;
        RECT 287.250 328.830 288.020 331.710 ;
        RECT 285.800 328.790 288.280 328.830 ;
        RECT 102.000 328.410 102.610 328.620 ;
        RECT 211.100 328.530 288.280 328.790 ;
        RECT 211.100 328.480 226.810 328.530 ;
        RECT 231.070 328.480 246.780 328.530 ;
        RECT 251.180 328.480 266.890 328.530 ;
        RECT 271.290 328.480 288.280 328.530 ;
        RECT 356.380 328.640 356.790 332.810 ;
        RECT 359.770 332.670 360.050 346.670 ;
        RECT 363.050 346.650 363.330 347.280 ;
        RECT 369.600 347.230 370.530 347.280 ;
        RECT 375.740 347.390 376.070 351.290 ;
        RECT 382.380 351.210 382.660 365.270 ;
        RECT 388.940 365.120 389.320 366.010 ;
        RECT 382.450 350.710 382.620 351.210 ;
        RECT 388.950 351.020 389.230 365.120 ;
        RECT 393.630 364.280 394.710 365.600 ;
        RECT 395.050 364.280 395.330 366.130 ;
        RECT 398.410 365.520 398.580 365.680 ;
        RECT 393.630 363.900 395.330 364.280 ;
        RECT 393.630 351.300 394.710 363.900 ;
        RECT 395.050 351.480 395.330 363.900 ;
        RECT 398.360 351.520 398.640 365.520 ;
        RECT 401.640 365.500 401.920 366.130 ;
        RECT 408.190 366.080 409.120 366.130 ;
        RECT 394.990 351.360 395.330 351.480 ;
        RECT 389.030 350.710 389.200 351.020 ;
        RECT 388.960 347.430 389.850 347.480 ;
        RECT 388.920 347.390 389.850 347.430 ;
        RECT 359.720 332.450 360.050 332.670 ;
        RECT 363.040 346.490 363.330 346.650 ;
        RECT 359.720 331.460 360.020 332.450 ;
        RECT 363.040 332.430 363.320 346.490 ;
        RECT 366.400 346.440 366.570 346.830 ;
        RECT 366.340 332.660 366.620 346.440 ;
        RECT 369.600 346.340 369.980 347.230 ;
        RECT 375.740 347.180 389.850 347.390 ;
        RECT 375.740 347.100 376.070 347.180 ;
        RECT 363.110 331.930 363.280 332.430 ;
        RECT 366.340 332.220 366.660 332.660 ;
        RECT 369.610 332.240 369.890 346.340 ;
        RECT 374.360 332.350 375.440 346.650 ;
        RECT 375.780 332.710 376.060 347.100 ;
        RECT 382.370 346.550 382.650 347.180 ;
        RECT 382.360 346.390 382.650 346.550 ;
        RECT 388.920 347.130 389.850 347.180 ;
        RECT 394.990 347.460 395.320 351.360 ;
        RECT 398.310 351.300 398.640 351.520 ;
        RECT 401.630 365.340 401.920 365.500 ;
        RECT 398.310 350.310 398.610 351.300 ;
        RECT 401.630 351.280 401.910 365.340 ;
        RECT 404.990 365.290 405.160 365.680 ;
        RECT 404.930 351.510 405.210 365.290 ;
        RECT 408.190 365.190 408.570 366.080 ;
        RECT 401.700 350.780 401.870 351.280 ;
        RECT 404.930 351.070 405.250 351.510 ;
        RECT 408.200 351.090 408.480 365.190 ;
        RECT 653.970 354.845 655.410 355.015 ;
        RECT 654.730 353.035 655.320 354.615 ;
        RECT 655.990 354.130 656.950 354.940 ;
        RECT 657.550 354.835 672.910 355.005 ;
        RECT 658.190 353.045 659.135 354.585 ;
        RECT 659.745 353.735 660.640 354.555 ;
        RECT 661.475 353.525 662.425 354.555 ;
        RECT 664.170 354.305 665.120 354.605 ;
        RECT 666.510 354.075 667.460 354.555 ;
        RECT 669.560 354.220 669.890 354.555 ;
        RECT 671.690 353.575 672.280 354.555 ;
        RECT 673.870 354.120 674.700 354.850 ;
        RECT 675.600 354.795 690.960 354.965 ;
        RECT 676.240 353.005 677.185 354.545 ;
        RECT 677.795 353.695 678.690 354.515 ;
        RECT 679.525 353.485 680.475 354.515 ;
        RECT 682.220 354.265 683.170 354.565 ;
        RECT 684.560 354.035 685.510 354.515 ;
        RECT 687.610 354.180 687.940 354.515 ;
        RECT 689.740 353.535 690.330 354.515 ;
        RECT 691.530 354.150 692.780 354.920 ;
        RECT 693.190 354.815 708.550 354.985 ;
        RECT 693.830 353.025 694.775 354.565 ;
        RECT 695.385 353.715 696.280 354.535 ;
        RECT 697.115 353.505 698.065 354.535 ;
        RECT 699.810 354.285 700.760 354.585 ;
        RECT 702.150 354.055 703.100 354.535 ;
        RECT 705.200 354.200 705.530 354.535 ;
        RECT 707.330 353.555 707.920 354.535 ;
        RECT 709.230 354.020 710.310 354.830 ;
        RECT 711.040 354.815 726.400 354.985 ;
        RECT 711.680 353.025 712.625 354.565 ;
        RECT 713.235 353.715 714.130 354.535 ;
        RECT 714.965 353.505 715.915 354.535 ;
        RECT 717.660 354.285 718.610 354.585 ;
        RECT 720.000 354.055 720.950 354.535 ;
        RECT 723.050 354.200 723.380 354.535 ;
        RECT 725.180 353.555 725.770 354.535 ;
        RECT 727.330 353.910 728.290 354.840 ;
        RECT 729.300 354.815 744.660 354.985 ;
        RECT 729.940 353.025 730.885 354.565 ;
        RECT 731.495 353.715 732.390 354.535 ;
        RECT 733.225 353.505 734.175 354.535 ;
        RECT 735.920 354.285 736.870 354.585 ;
        RECT 738.260 354.055 739.210 354.535 ;
        RECT 741.310 354.200 741.640 354.535 ;
        RECT 743.440 353.555 744.030 354.535 ;
        RECT 745.210 354.140 746.480 354.940 ;
        RECT 747.070 354.785 762.430 354.955 ;
        RECT 747.710 352.995 748.655 354.535 ;
        RECT 749.265 353.685 750.160 354.505 ;
        RECT 750.995 353.475 751.945 354.505 ;
        RECT 753.690 354.255 754.640 354.555 ;
        RECT 756.030 354.025 756.980 354.505 ;
        RECT 759.080 354.170 759.410 354.505 ;
        RECT 761.210 353.525 761.800 354.505 ;
        RECT 763.250 354.070 764.080 354.730 ;
        RECT 765.110 354.705 780.470 354.875 ;
        RECT 765.750 352.915 766.695 354.455 ;
        RECT 767.305 353.605 768.200 354.425 ;
        RECT 769.035 353.395 769.985 354.425 ;
        RECT 771.730 354.175 772.680 354.475 ;
        RECT 774.070 353.945 775.020 354.425 ;
        RECT 777.120 354.090 777.450 354.425 ;
        RECT 779.250 353.445 779.840 354.425 ;
        RECT 781.260 354.020 782.430 354.820 ;
        RECT 783.270 354.745 798.630 354.915 ;
        RECT 783.910 352.955 784.855 354.495 ;
        RECT 785.465 353.645 786.360 354.465 ;
        RECT 787.195 353.435 788.145 354.465 ;
        RECT 789.890 354.215 790.840 354.515 ;
        RECT 792.230 353.985 793.180 354.465 ;
        RECT 795.280 354.130 795.610 354.465 ;
        RECT 797.410 353.485 798.000 354.465 ;
        RECT 799.490 353.740 800.420 354.780 ;
        RECT 801.650 354.755 817.010 354.925 ;
        RECT 802.290 352.965 803.235 354.505 ;
        RECT 803.845 353.655 804.740 354.475 ;
        RECT 805.575 353.445 806.525 354.475 ;
        RECT 808.270 354.225 809.220 354.525 ;
        RECT 810.610 353.995 811.560 354.475 ;
        RECT 813.660 354.140 813.990 354.475 ;
        RECT 815.790 353.495 816.380 354.475 ;
        RECT 817.790 354.110 819.140 354.880 ;
        RECT 820.450 354.735 835.810 354.905 ;
        RECT 821.090 352.945 822.035 354.485 ;
        RECT 822.645 353.635 823.540 354.455 ;
        RECT 824.375 353.425 825.325 354.455 ;
        RECT 827.070 354.205 828.020 354.505 ;
        RECT 829.410 353.975 830.360 354.455 ;
        RECT 832.460 354.120 832.790 354.455 ;
        RECT 834.590 353.475 835.180 354.455 ;
        RECT 836.990 353.750 837.920 354.840 ;
        RECT 838.920 354.715 840.360 354.885 ;
        RECT 839.680 352.905 840.270 354.485 ;
        RECT 832.065 351.560 832.395 352.855 ;
        RECT 404.950 350.330 405.250 351.070 ;
        RECT 408.280 350.780 408.450 351.090 ;
        RECT 404.950 350.310 405.740 350.330 ;
        RECT 398.310 350.000 405.740 350.310 ;
        RECT 398.310 349.970 398.610 350.000 ;
        RECT 404.860 349.980 405.250 350.000 ;
        RECT 404.950 349.960 405.250 349.980 ;
        RECT 408.210 347.500 409.100 347.550 ;
        RECT 408.170 347.460 409.100 347.500 ;
        RECT 394.990 347.250 409.100 347.460 ;
        RECT 394.990 347.170 395.320 347.250 ;
        RECT 366.360 331.480 366.660 332.220 ;
        RECT 369.690 331.930 369.860 332.240 ;
        RECT 366.360 331.460 367.150 331.480 ;
        RECT 359.720 331.150 367.150 331.460 ;
        RECT 359.720 331.120 360.020 331.150 ;
        RECT 366.360 331.110 366.660 331.150 ;
        RECT 369.640 328.680 370.530 328.730 ;
        RECT 369.600 328.640 370.530 328.680 ;
        RECT 356.380 328.480 370.530 328.640 ;
        RECT 211.100 328.470 212.510 328.480 ;
        RECT 231.070 328.470 232.480 328.480 ;
        RECT 251.180 328.470 252.590 328.480 ;
        RECT 271.290 328.470 272.700 328.480 ;
        RECT 211.120 328.460 211.530 328.470 ;
        RECT 231.090 328.460 231.500 328.470 ;
        RECT 251.200 328.460 251.610 328.470 ;
        RECT 271.310 328.460 271.720 328.470 ;
        RECT 11.940 328.200 102.780 328.410 ;
        RECT 285.800 328.210 288.280 328.480 ;
        RECT 356.440 328.430 370.530 328.480 ;
        RECT 11.940 328.160 102.900 328.200 ;
        RECT 11.940 327.940 102.940 328.160 ;
        RECT 4.680 327.620 102.940 327.940 ;
        RECT 11.940 327.560 102.940 327.620 ;
        RECT 3.870 324.620 5.470 324.730 ;
        RECT 3.870 324.610 12.510 324.620 ;
        RECT 3.780 324.560 12.510 324.610 ;
        RECT 3.780 324.390 12.710 324.560 ;
        RECT 3.780 324.360 12.510 324.390 ;
        RECT 3.780 324.120 5.470 324.360 ;
        RECT 3.780 318.120 4.240 324.120 ;
        RECT 13.190 321.310 13.530 327.560 ;
        RECT 17.210 324.600 18.810 324.710 ;
        RECT 17.210 324.590 25.850 324.600 ;
        RECT 4.920 321.270 13.530 321.310 ;
        RECT 4.750 321.100 13.530 321.270 ;
        RECT 4.920 321.050 13.530 321.100 ;
        RECT 12.090 321.040 13.530 321.050 ;
        RECT 3.780 318.010 5.400 318.120 ;
        RECT 3.780 317.980 12.530 318.010 ;
        RECT 3.780 317.810 12.710 317.980 ;
        RECT 3.780 317.750 12.530 317.810 ;
        RECT 3.780 317.510 5.400 317.750 ;
        RECT 3.780 311.550 4.240 317.510 ;
        RECT 13.190 314.750 13.530 321.040 ;
        RECT 12.150 314.740 13.530 314.750 ;
        RECT 4.990 314.690 13.530 314.740 ;
        RECT 4.750 314.520 13.530 314.690 ;
        RECT 4.990 314.480 13.530 314.520 ;
        RECT 3.750 311.440 5.350 311.550 ;
        RECT 3.750 311.400 12.580 311.440 ;
        RECT 3.750 311.230 12.710 311.400 ;
        RECT 3.750 311.180 12.580 311.230 ;
        RECT 3.750 310.940 5.350 311.180 ;
        RECT 3.780 305.110 4.240 310.940 ;
        RECT 13.190 308.160 13.530 314.480 ;
        RECT 17.120 324.540 25.850 324.590 ;
        RECT 17.120 324.370 26.050 324.540 ;
        RECT 17.120 324.340 25.850 324.370 ;
        RECT 17.120 324.100 18.810 324.340 ;
        RECT 17.120 318.100 17.580 324.100 ;
        RECT 26.530 321.290 26.870 327.560 ;
        RECT 30.580 324.630 32.180 324.740 ;
        RECT 30.580 324.620 39.220 324.630 ;
        RECT 18.260 321.250 26.870 321.290 ;
        RECT 18.090 321.080 26.870 321.250 ;
        RECT 18.260 321.030 26.870 321.080 ;
        RECT 25.430 321.020 26.870 321.030 ;
        RECT 17.120 317.990 18.740 318.100 ;
        RECT 17.120 317.960 25.870 317.990 ;
        RECT 17.120 317.790 26.050 317.960 ;
        RECT 17.120 317.730 25.870 317.790 ;
        RECT 17.120 317.490 18.740 317.730 ;
        RECT 17.120 311.530 17.580 317.490 ;
        RECT 26.530 314.730 26.870 321.020 ;
        RECT 25.490 314.720 26.870 314.730 ;
        RECT 18.330 314.670 26.870 314.720 ;
        RECT 18.090 314.500 26.870 314.670 ;
        RECT 18.330 314.460 26.870 314.500 ;
        RECT 17.090 311.420 18.690 311.530 ;
        RECT 17.090 311.380 25.920 311.420 ;
        RECT 17.090 311.210 26.050 311.380 ;
        RECT 17.090 311.160 25.920 311.210 ;
        RECT 17.090 310.920 18.690 311.160 ;
        RECT 12.100 308.150 13.530 308.160 ;
        RECT 5.110 308.110 13.530 308.150 ;
        RECT 4.750 307.940 13.530 308.110 ;
        RECT 5.110 307.890 13.530 307.940 ;
        RECT 3.700 304.870 5.300 305.110 ;
        RECT 3.700 304.610 12.820 304.870 ;
        RECT 13.190 304.730 13.530 307.890 ;
        RECT 3.700 304.500 5.300 304.610 ;
        RECT 13.140 304.520 13.530 304.730 ;
        RECT 15.430 305.050 16.520 305.350 ;
        RECT 17.120 305.090 17.580 310.920 ;
        RECT 26.530 308.140 26.870 314.460 ;
        RECT 30.490 324.570 39.220 324.620 ;
        RECT 30.490 324.400 39.420 324.570 ;
        RECT 30.490 324.370 39.220 324.400 ;
        RECT 30.490 324.130 32.180 324.370 ;
        RECT 30.490 318.130 30.950 324.130 ;
        RECT 39.900 321.320 40.240 327.560 ;
        RECT 43.810 324.630 45.410 324.740 ;
        RECT 43.810 324.620 52.450 324.630 ;
        RECT 31.630 321.280 40.240 321.320 ;
        RECT 31.460 321.110 40.240 321.280 ;
        RECT 31.630 321.060 40.240 321.110 ;
        RECT 38.800 321.050 40.240 321.060 ;
        RECT 30.490 318.020 32.110 318.130 ;
        RECT 30.490 317.990 39.240 318.020 ;
        RECT 30.490 317.820 39.420 317.990 ;
        RECT 30.490 317.760 39.240 317.820 ;
        RECT 30.490 317.520 32.110 317.760 ;
        RECT 30.490 311.560 30.950 317.520 ;
        RECT 39.900 314.760 40.240 321.050 ;
        RECT 38.860 314.750 40.240 314.760 ;
        RECT 31.700 314.700 40.240 314.750 ;
        RECT 31.460 314.530 40.240 314.700 ;
        RECT 31.700 314.490 40.240 314.530 ;
        RECT 30.460 311.450 32.060 311.560 ;
        RECT 30.460 311.410 39.290 311.450 ;
        RECT 30.460 311.240 39.420 311.410 ;
        RECT 30.460 311.190 39.290 311.240 ;
        RECT 30.460 310.950 32.060 311.190 ;
        RECT 25.440 308.130 26.870 308.140 ;
        RECT 18.450 308.090 26.870 308.130 ;
        RECT 18.090 307.920 26.870 308.090 ;
        RECT 18.450 307.870 26.870 307.920 ;
        RECT 17.040 305.050 18.640 305.090 ;
        RECT 15.430 304.850 18.640 305.050 ;
        RECT 15.430 304.590 26.160 304.850 ;
        RECT 26.530 304.710 26.870 307.870 ;
        RECT 13.140 301.600 13.510 304.520 ;
        RECT 15.430 304.480 18.640 304.590 ;
        RECT 26.480 304.500 26.870 304.710 ;
        RECT 28.600 305.100 29.780 305.520 ;
        RECT 30.490 305.120 30.950 310.950 ;
        RECT 39.900 308.170 40.240 314.490 ;
        RECT 43.720 324.570 52.450 324.620 ;
        RECT 43.720 324.400 52.650 324.570 ;
        RECT 43.720 324.370 52.450 324.400 ;
        RECT 43.720 324.130 45.410 324.370 ;
        RECT 43.720 318.130 44.180 324.130 ;
        RECT 53.130 321.320 53.470 327.560 ;
        RECT 57.080 324.600 58.680 324.710 ;
        RECT 57.080 324.590 65.720 324.600 ;
        RECT 44.860 321.280 53.470 321.320 ;
        RECT 44.690 321.110 53.470 321.280 ;
        RECT 44.860 321.060 53.470 321.110 ;
        RECT 52.030 321.050 53.470 321.060 ;
        RECT 43.720 318.020 45.340 318.130 ;
        RECT 43.720 317.990 52.470 318.020 ;
        RECT 43.720 317.820 52.650 317.990 ;
        RECT 43.720 317.760 52.470 317.820 ;
        RECT 43.720 317.520 45.340 317.760 ;
        RECT 43.720 311.560 44.180 317.520 ;
        RECT 53.130 314.760 53.470 321.050 ;
        RECT 52.090 314.750 53.470 314.760 ;
        RECT 44.930 314.700 53.470 314.750 ;
        RECT 44.690 314.530 53.470 314.700 ;
        RECT 44.930 314.490 53.470 314.530 ;
        RECT 43.690 311.450 45.290 311.560 ;
        RECT 43.690 311.410 52.520 311.450 ;
        RECT 43.690 311.240 52.650 311.410 ;
        RECT 43.690 311.190 52.520 311.240 ;
        RECT 43.690 310.950 45.290 311.190 ;
        RECT 38.810 308.160 40.240 308.170 ;
        RECT 31.820 308.120 40.240 308.160 ;
        RECT 31.460 307.950 40.240 308.120 ;
        RECT 31.820 307.900 40.240 307.950 ;
        RECT 30.410 305.100 32.010 305.120 ;
        RECT 28.600 304.880 32.010 305.100 ;
        RECT 28.600 304.620 39.530 304.880 ;
        RECT 39.900 304.740 40.240 307.900 ;
        RECT 28.600 304.550 32.010 304.620 ;
        RECT 15.430 304.340 17.660 304.480 ;
        RECT 15.430 303.580 16.520 304.340 ;
        RECT 12.420 301.570 13.530 301.600 ;
        RECT 26.480 301.580 26.850 304.500 ;
        RECT 28.600 303.710 29.780 304.550 ;
        RECT 30.410 304.510 32.010 304.550 ;
        RECT 39.850 304.530 40.240 304.740 ;
        RECT 41.900 305.180 42.910 305.900 ;
        RECT 43.720 305.180 44.180 310.950 ;
        RECT 53.130 308.170 53.470 314.490 ;
        RECT 56.990 324.540 65.720 324.590 ;
        RECT 56.990 324.370 65.920 324.540 ;
        RECT 56.990 324.340 65.720 324.370 ;
        RECT 56.990 324.100 58.680 324.340 ;
        RECT 56.990 318.100 57.450 324.100 ;
        RECT 66.400 321.290 66.740 327.560 ;
        RECT 70.350 324.630 71.950 324.740 ;
        RECT 70.350 324.620 78.990 324.630 ;
        RECT 58.130 321.250 66.740 321.290 ;
        RECT 57.960 321.080 66.740 321.250 ;
        RECT 58.130 321.030 66.740 321.080 ;
        RECT 65.300 321.020 66.740 321.030 ;
        RECT 56.990 317.990 58.610 318.100 ;
        RECT 56.990 317.960 65.740 317.990 ;
        RECT 56.990 317.790 65.920 317.960 ;
        RECT 56.990 317.730 65.740 317.790 ;
        RECT 56.990 317.490 58.610 317.730 ;
        RECT 56.990 311.530 57.450 317.490 ;
        RECT 66.400 314.730 66.740 321.020 ;
        RECT 65.360 314.720 66.740 314.730 ;
        RECT 58.200 314.670 66.740 314.720 ;
        RECT 57.960 314.500 66.740 314.670 ;
        RECT 58.200 314.460 66.740 314.500 ;
        RECT 56.960 311.420 58.560 311.530 ;
        RECT 56.960 311.380 65.790 311.420 ;
        RECT 56.960 311.210 65.920 311.380 ;
        RECT 56.960 311.160 65.790 311.210 ;
        RECT 56.960 310.920 58.560 311.160 ;
        RECT 52.040 308.160 53.470 308.170 ;
        RECT 45.050 308.120 53.470 308.160 ;
        RECT 44.690 307.950 53.470 308.120 ;
        RECT 45.050 307.900 53.470 307.950 ;
        RECT 41.900 305.120 44.250 305.180 ;
        RECT 41.900 304.880 45.240 305.120 ;
        RECT 41.900 304.620 52.760 304.880 ;
        RECT 53.130 304.740 53.470 307.900 ;
        RECT 41.900 304.550 45.240 304.620 ;
        RECT 39.850 301.610 40.220 304.530 ;
        RECT 41.900 303.460 42.910 304.550 ;
        RECT 43.640 304.510 45.240 304.550 ;
        RECT 53.080 304.530 53.470 304.740 ;
        RECT 55.280 305.140 56.370 305.480 ;
        RECT 56.990 305.140 57.450 310.920 ;
        RECT 66.400 308.140 66.740 314.460 ;
        RECT 70.260 324.570 78.990 324.620 ;
        RECT 70.260 324.400 79.190 324.570 ;
        RECT 70.260 324.370 78.990 324.400 ;
        RECT 70.260 324.130 71.950 324.370 ;
        RECT 70.260 318.130 70.720 324.130 ;
        RECT 79.670 321.320 80.010 327.560 ;
        RECT 83.480 324.650 85.080 324.760 ;
        RECT 83.480 324.640 92.120 324.650 ;
        RECT 71.400 321.280 80.010 321.320 ;
        RECT 71.230 321.110 80.010 321.280 ;
        RECT 71.400 321.060 80.010 321.110 ;
        RECT 78.570 321.050 80.010 321.060 ;
        RECT 70.260 318.020 71.880 318.130 ;
        RECT 70.260 317.990 79.010 318.020 ;
        RECT 70.260 317.820 79.190 317.990 ;
        RECT 70.260 317.760 79.010 317.820 ;
        RECT 70.260 317.520 71.880 317.760 ;
        RECT 70.260 311.560 70.720 317.520 ;
        RECT 79.670 314.760 80.010 321.050 ;
        RECT 78.630 314.750 80.010 314.760 ;
        RECT 71.470 314.700 80.010 314.750 ;
        RECT 71.230 314.530 80.010 314.700 ;
        RECT 71.470 314.490 80.010 314.530 ;
        RECT 70.230 311.450 71.830 311.560 ;
        RECT 70.230 311.410 79.060 311.450 ;
        RECT 70.230 311.240 79.190 311.410 ;
        RECT 70.230 311.190 79.060 311.240 ;
        RECT 70.230 310.950 71.830 311.190 ;
        RECT 65.310 308.130 66.740 308.140 ;
        RECT 58.320 308.090 66.740 308.130 ;
        RECT 57.960 307.920 66.740 308.090 ;
        RECT 58.320 307.870 66.740 307.920 ;
        RECT 55.280 304.850 59.740 305.140 ;
        RECT 55.280 304.590 66.030 304.850 ;
        RECT 66.400 304.710 66.740 307.870 ;
        RECT 55.280 304.550 59.740 304.590 ;
        RECT 53.080 301.610 53.450 304.530 ;
        RECT 55.280 303.290 56.370 304.550 ;
        RECT 56.910 304.480 58.510 304.550 ;
        RECT 66.350 304.500 66.740 304.710 ;
        RECT 68.530 305.010 69.370 305.640 ;
        RECT 70.260 305.120 70.720 310.950 ;
        RECT 79.670 308.170 80.010 314.490 ;
        RECT 83.390 324.590 92.120 324.640 ;
        RECT 83.390 324.420 92.320 324.590 ;
        RECT 83.390 324.390 92.120 324.420 ;
        RECT 83.390 324.150 85.080 324.390 ;
        RECT 83.390 318.150 83.850 324.150 ;
        RECT 92.800 321.340 93.140 327.560 ;
        RECT 96.820 324.890 98.230 324.940 ;
        RECT 96.820 324.830 102.210 324.890 ;
        RECT 102.530 324.830 102.940 327.560 ;
        RECT 96.820 324.600 103.230 324.830 ;
        RECT 96.820 324.460 98.230 324.600 ;
        RECT 101.980 324.580 103.230 324.600 ;
        RECT 84.530 321.300 93.140 321.340 ;
        RECT 84.360 321.130 93.140 321.300 ;
        RECT 84.530 321.080 93.140 321.130 ;
        RECT 91.700 321.070 93.140 321.080 ;
        RECT 83.390 318.040 85.010 318.150 ;
        RECT 83.390 318.010 92.140 318.040 ;
        RECT 83.390 317.840 92.320 318.010 ;
        RECT 83.390 317.780 92.140 317.840 ;
        RECT 83.390 317.540 85.010 317.780 ;
        RECT 83.390 311.580 83.850 317.540 ;
        RECT 92.800 314.780 93.140 321.070 ;
        RECT 91.760 314.770 93.140 314.780 ;
        RECT 84.600 314.720 93.140 314.770 ;
        RECT 84.360 314.550 93.140 314.720 ;
        RECT 84.600 314.510 93.140 314.550 ;
        RECT 83.360 311.470 84.960 311.580 ;
        RECT 83.360 311.430 92.190 311.470 ;
        RECT 83.360 311.260 92.320 311.430 ;
        RECT 83.360 311.210 92.190 311.260 ;
        RECT 83.360 310.970 84.960 311.210 ;
        RECT 78.580 308.160 80.010 308.170 ;
        RECT 71.590 308.120 80.010 308.160 ;
        RECT 71.230 307.950 80.010 308.120 ;
        RECT 71.590 307.900 80.010 307.950 ;
        RECT 70.180 305.010 71.780 305.120 ;
        RECT 68.530 304.880 72.440 305.010 ;
        RECT 68.530 304.620 79.300 304.880 ;
        RECT 79.670 304.740 80.010 307.900 ;
        RECT 39.130 301.580 40.240 301.610 ;
        RECT 52.360 301.580 53.470 301.610 ;
        RECT 66.350 301.580 66.720 304.500 ;
        RECT 68.530 304.420 72.440 304.620 ;
        RECT 79.620 304.530 80.010 304.740 ;
        RECT 81.610 305.180 82.880 305.350 ;
        RECT 83.390 305.180 83.850 310.970 ;
        RECT 92.800 308.190 93.140 314.510 ;
        RECT 96.900 318.360 97.240 324.460 ;
        RECT 98.200 321.540 102.210 321.570 ;
        RECT 102.530 321.540 102.940 324.580 ;
        RECT 213.670 323.470 226.900 325.480 ;
        RECT 265.770 325.470 268.720 325.670 ;
        RECT 285.800 325.470 286.630 328.210 ;
        RECT 233.710 323.460 246.940 325.470 ;
        RECT 253.770 323.550 268.720 325.470 ;
        RECT 253.770 323.460 267.000 323.550 ;
        RECT 273.820 323.460 287.050 325.470 ;
        RECT 226.330 322.860 227.650 322.930 ;
        RECT 246.370 322.860 247.690 322.920 ;
        RECT 266.430 322.860 267.750 322.920 ;
        RECT 284.260 322.860 284.830 323.460 ;
        RECT 286.480 322.880 287.800 322.920 ;
        RECT 286.480 322.860 289.780 322.880 ;
        RECT 212.240 322.780 289.780 322.860 ;
        RECT 211.870 322.610 289.780 322.780 ;
        RECT 212.240 322.600 289.780 322.610 ;
        RECT 212.320 322.570 227.650 322.600 ;
        RECT 226.330 322.550 227.650 322.570 ;
        RECT 232.360 322.560 247.690 322.600 ;
        RECT 252.420 322.560 267.750 322.600 ;
        RECT 272.470 322.560 289.780 322.600 ;
        RECT 98.200 321.520 102.940 321.540 ;
        RECT 97.780 321.350 102.940 321.520 ;
        RECT 98.200 321.280 102.940 321.350 ;
        RECT 101.660 321.190 102.940 321.280 ;
        RECT 102.530 320.600 102.940 321.190 ;
        RECT 103.460 320.600 104.050 320.720 ;
        RECT 102.530 320.350 104.050 320.600 ;
        RECT 96.900 318.310 98.330 318.360 ;
        RECT 96.900 318.230 102.250 318.310 ;
        RECT 96.900 318.060 102.270 318.230 ;
        RECT 96.900 318.020 102.250 318.060 ;
        RECT 96.900 317.880 98.330 318.020 ;
        RECT 96.900 311.720 97.240 317.880 ;
        RECT 98.260 314.950 102.270 314.970 ;
        RECT 102.530 314.950 102.940 320.350 ;
        RECT 103.460 320.160 104.050 320.350 ;
        RECT 227.260 316.290 227.530 322.550 ;
        RECT 246.370 322.540 247.690 322.560 ;
        RECT 266.430 322.540 267.750 322.560 ;
        RECT 226.510 316.260 227.830 316.290 ;
        RECT 247.300 316.280 247.570 322.540 ;
        RECT 267.360 316.280 267.630 322.540 ;
        RECT 284.260 322.520 284.830 322.560 ;
        RECT 286.480 322.540 289.780 322.560 ;
        RECT 287.040 322.100 289.780 322.540 ;
        RECT 287.410 316.280 287.680 322.100 ;
        RECT 212.560 316.200 227.830 316.260 ;
        RECT 246.550 316.250 247.870 316.280 ;
        RECT 266.610 316.250 267.930 316.280 ;
        RECT 286.660 316.250 287.980 316.280 ;
        RECT 211.870 316.030 227.830 316.200 ;
        RECT 232.600 316.190 247.870 316.250 ;
        RECT 252.660 316.190 267.930 316.250 ;
        RECT 272.710 316.190 287.980 316.250 ;
        RECT 212.560 315.990 227.830 316.030 ;
        RECT 231.910 316.020 247.870 316.190 ;
        RECT 251.970 316.020 267.930 316.190 ;
        RECT 272.020 316.020 287.980 316.190 ;
        RECT 226.510 315.910 227.830 315.990 ;
        RECT 232.600 315.980 247.870 316.020 ;
        RECT 252.660 315.980 267.930 316.020 ;
        RECT 272.710 315.980 287.980 316.020 ;
        RECT 98.260 314.940 103.030 314.950 ;
        RECT 97.780 314.770 103.030 314.940 ;
        RECT 98.260 314.680 103.030 314.770 ;
        RECT 101.810 314.600 103.030 314.680 ;
        RECT 96.880 311.650 102.190 311.720 ;
        RECT 96.880 311.480 102.270 311.650 ;
        RECT 96.880 311.430 102.190 311.480 ;
        RECT 96.880 311.240 98.290 311.430 ;
        RECT 91.710 308.180 93.140 308.190 ;
        RECT 84.720 308.140 93.140 308.180 ;
        RECT 84.360 307.970 93.140 308.140 ;
        RECT 84.720 307.920 93.140 307.970 ;
        RECT 81.610 304.900 85.310 305.180 ;
        RECT 81.610 304.640 92.430 304.900 ;
        RECT 92.800 304.760 93.140 307.920 ;
        RECT 68.530 303.500 69.370 304.420 ;
        RECT 79.620 301.610 79.990 304.530 ;
        RECT 81.610 304.390 85.310 304.640 ;
        RECT 92.750 304.550 93.140 304.760 ;
        RECT 94.360 305.560 95.410 305.810 ;
        RECT 96.900 305.560 97.240 311.240 ;
        RECT 102.530 308.430 102.940 314.600 ;
        RECT 227.260 309.720 227.530 315.910 ;
        RECT 246.550 315.900 247.870 315.980 ;
        RECT 266.610 315.900 267.930 315.980 ;
        RECT 286.660 315.900 287.980 315.980 ;
        RECT 226.360 309.650 227.680 309.720 ;
        RECT 247.300 309.710 247.570 315.900 ;
        RECT 267.360 309.710 267.630 315.900 ;
        RECT 287.410 309.710 287.680 315.900 ;
        RECT 355.040 313.600 356.120 327.900 ;
        RECT 356.460 314.190 356.740 328.430 ;
        RECT 359.820 327.820 359.990 327.980 ;
        RECT 356.440 309.820 356.740 314.190 ;
        RECT 359.770 313.820 360.050 327.820 ;
        RECT 363.050 327.800 363.330 328.430 ;
        RECT 369.600 328.380 370.530 328.430 ;
        RECT 375.700 328.540 376.110 332.710 ;
        RECT 382.360 332.330 382.640 346.390 ;
        RECT 388.920 346.240 389.300 347.130 ;
        RECT 382.430 331.830 382.600 332.330 ;
        RECT 388.930 332.140 389.210 346.240 ;
        RECT 393.610 332.420 394.690 346.720 ;
        RECT 395.030 332.780 395.310 347.170 ;
        RECT 398.390 346.640 398.560 346.800 ;
        RECT 389.010 331.830 389.180 332.140 ;
        RECT 388.960 328.580 389.850 328.630 ;
        RECT 388.920 328.540 389.850 328.580 ;
        RECT 375.700 328.380 389.850 328.540 ;
        RECT 394.950 328.610 395.360 332.780 ;
        RECT 398.340 332.640 398.620 346.640 ;
        RECT 401.620 346.620 401.900 347.250 ;
        RECT 408.170 347.200 409.100 347.250 ;
        RECT 398.290 332.420 398.620 332.640 ;
        RECT 401.610 346.460 401.900 346.620 ;
        RECT 398.290 331.430 398.590 332.420 ;
        RECT 401.610 332.400 401.890 346.460 ;
        RECT 404.970 346.410 405.140 346.800 ;
        RECT 404.910 332.630 405.190 346.410 ;
        RECT 408.170 346.310 408.550 347.200 ;
        RECT 783.830 346.575 787.190 346.745 ;
        RECT 401.680 331.900 401.850 332.400 ;
        RECT 404.910 332.190 405.230 332.630 ;
        RECT 408.180 332.210 408.460 346.310 ;
        RECT 784.390 344.845 785.640 346.345 ;
        RECT 786.170 344.845 787.100 346.295 ;
        RECT 788.280 346.140 789.060 346.710 ;
        RECT 790.390 346.605 791.830 346.775 ;
        RECT 791.150 344.795 791.740 346.375 ;
        RECT 792.440 346.080 793.190 346.700 ;
        RECT 793.850 346.665 809.210 346.835 ;
        RECT 794.490 344.875 795.435 346.415 ;
        RECT 796.045 345.565 796.940 346.385 ;
        RECT 797.775 345.355 798.725 346.385 ;
        RECT 800.470 346.135 801.420 346.435 ;
        RECT 802.810 345.905 803.760 346.385 ;
        RECT 805.860 346.050 806.190 346.385 ;
        RECT 807.990 345.405 808.580 346.385 ;
        RECT 810.590 346.010 811.400 346.720 ;
        RECT 813.210 346.575 828.570 346.745 ;
        RECT 813.850 344.785 814.795 346.325 ;
        RECT 815.405 345.475 816.300 346.295 ;
        RECT 817.135 345.265 818.085 346.295 ;
        RECT 819.830 346.045 820.780 346.345 ;
        RECT 822.170 345.815 823.120 346.295 ;
        RECT 825.220 345.960 825.550 346.295 ;
        RECT 827.350 345.315 827.940 346.295 ;
        RECT 829.180 345.820 829.950 346.670 ;
        RECT 404.930 331.450 405.230 332.190 ;
        RECT 408.260 331.900 408.430 332.210 ;
        RECT 404.930 331.430 405.720 331.450 ;
        RECT 398.290 331.120 405.720 331.430 ;
        RECT 398.290 331.090 398.590 331.120 ;
        RECT 404.930 331.080 405.230 331.120 ;
        RECT 595.370 330.695 596.810 330.865 ;
        RECT 596.130 328.885 596.720 330.465 ;
        RECT 601.180 330.000 601.920 332.860 ;
        RECT 602.630 332.050 602.800 332.470 ;
        RECT 604.210 332.050 604.380 332.470 ;
        RECT 605.790 332.050 605.960 332.470 ;
        RECT 607.150 332.060 607.320 332.480 ;
        RECT 608.730 332.060 608.900 332.480 ;
        RECT 610.310 332.060 610.480 332.480 ;
        RECT 611.670 332.060 611.840 332.480 ;
        RECT 613.250 332.060 613.420 332.480 ;
        RECT 614.830 332.060 615.000 332.480 ;
        RECT 616.100 332.040 616.270 332.460 ;
        RECT 617.680 332.040 617.850 332.460 ;
        RECT 619.260 332.040 619.430 332.460 ;
        RECT 620.480 332.050 620.650 332.470 ;
        RECT 622.060 332.050 622.230 332.470 ;
        RECT 623.640 332.050 623.810 332.470 ;
        RECT 624.800 332.040 624.970 332.460 ;
        RECT 626.380 332.040 626.550 332.460 ;
        RECT 627.960 332.040 628.130 332.460 ;
        RECT 602.630 330.580 602.800 331.000 ;
        RECT 604.210 330.580 604.380 331.000 ;
        RECT 605.790 330.580 605.960 331.000 ;
        RECT 607.150 330.590 607.320 331.010 ;
        RECT 608.730 330.590 608.900 331.010 ;
        RECT 610.310 330.590 610.480 331.010 ;
        RECT 611.670 330.590 611.840 331.010 ;
        RECT 613.250 330.590 613.420 331.010 ;
        RECT 614.830 330.590 615.000 331.010 ;
        RECT 616.100 330.570 616.270 330.990 ;
        RECT 617.680 330.570 617.850 330.990 ;
        RECT 619.260 330.570 619.430 330.990 ;
        RECT 620.480 330.580 620.650 331.000 ;
        RECT 622.060 330.580 622.230 331.000 ;
        RECT 623.640 330.580 623.810 331.000 ;
        RECT 624.800 330.570 624.970 330.990 ;
        RECT 626.380 330.570 626.550 330.990 ;
        RECT 627.960 330.570 628.130 330.990 ;
        RECT 628.880 329.830 629.750 333.150 ;
        RECT 663.190 332.485 666.550 332.655 ;
        RECT 668.820 332.485 672.180 332.655 ;
        RECT 674.580 332.385 677.940 332.555 ;
        RECT 681.610 332.425 685.450 332.595 ;
        RECT 687.470 332.435 690.830 332.605 ;
        RECT 635.260 331.145 636.700 331.315 ;
        RECT 639.450 331.235 640.890 331.405 ;
        RECT 643.550 331.215 644.990 331.385 ;
        RECT 635.350 329.335 635.940 330.915 ;
        RECT 639.540 329.425 640.130 331.005 ;
        RECT 643.640 329.405 644.230 330.985 ;
        RECT 645.340 329.590 645.980 330.900 ;
        RECT 663.280 330.755 664.210 332.205 ;
        RECT 664.740 330.755 665.990 332.255 ;
        RECT 668.910 330.755 669.840 332.205 ;
        RECT 670.370 330.755 671.620 332.255 ;
        RECT 675.410 330.655 677.380 332.155 ;
        RECT 678.370 330.930 679.130 331.840 ;
        RECT 682.170 331.110 683.120 332.145 ;
        RECT 683.810 330.615 684.760 332.195 ;
        RECT 687.560 330.705 688.490 332.155 ;
        RECT 689.020 330.705 690.270 332.205 ;
        RECT 862.390 329.040 863.760 331.120 ;
        RECT 408.210 328.650 409.100 328.700 ;
        RECT 408.170 328.610 409.100 328.650 ;
        RECT 394.950 328.450 409.100 328.610 ;
        RECT 395.010 328.400 409.100 328.450 ;
        RECT 359.720 313.600 360.050 313.820 ;
        RECT 363.040 327.640 363.330 327.800 ;
        RECT 359.720 312.610 360.020 313.600 ;
        RECT 363.040 313.580 363.320 327.640 ;
        RECT 366.400 327.590 366.570 327.980 ;
        RECT 366.340 313.810 366.620 327.590 ;
        RECT 369.600 327.490 369.980 328.380 ;
        RECT 375.760 328.330 389.850 328.380 ;
        RECT 363.110 313.080 363.280 313.580 ;
        RECT 366.340 313.370 366.660 313.810 ;
        RECT 369.610 313.390 369.890 327.490 ;
        RECT 374.360 313.500 375.440 327.800 ;
        RECT 375.780 314.090 376.060 328.330 ;
        RECT 382.370 327.700 382.650 328.330 ;
        RECT 366.360 312.630 366.660 313.370 ;
        RECT 369.690 313.080 369.860 313.390 ;
        RECT 366.360 312.610 367.150 312.630 ;
        RECT 359.720 312.300 367.150 312.610 ;
        RECT 359.720 312.270 360.020 312.300 ;
        RECT 366.360 312.260 366.660 312.300 ;
        RECT 369.640 309.860 370.530 309.910 ;
        RECT 369.600 309.820 370.530 309.860 ;
        RECT 212.550 309.620 227.680 309.650 ;
        RECT 246.400 309.640 247.720 309.710 ;
        RECT 266.460 309.640 267.780 309.710 ;
        RECT 286.510 309.640 287.830 309.710 ;
        RECT 211.870 309.450 227.680 309.620 ;
        RECT 232.590 309.610 247.720 309.640 ;
        RECT 252.650 309.610 267.780 309.640 ;
        RECT 272.700 309.610 287.830 309.640 ;
        RECT 356.440 309.610 370.530 309.820 ;
        RECT 212.550 309.380 227.680 309.450 ;
        RECT 231.910 309.440 247.720 309.610 ;
        RECT 251.970 309.440 267.780 309.610 ;
        RECT 272.020 309.440 287.830 309.610 ;
        RECT 226.360 309.340 227.680 309.380 ;
        RECT 232.590 309.370 247.720 309.440 ;
        RECT 252.650 309.370 267.780 309.440 ;
        RECT 272.700 309.370 287.830 309.440 ;
        RECT 227.260 309.330 227.530 309.340 ;
        RECT 246.400 309.330 247.720 309.370 ;
        RECT 266.460 309.330 267.780 309.370 ;
        RECT 286.510 309.330 287.830 309.370 ;
        RECT 247.300 309.320 247.570 309.330 ;
        RECT 267.360 309.320 267.630 309.330 ;
        RECT 101.720 308.370 102.940 308.430 ;
        RECT 98.180 308.360 102.940 308.370 ;
        RECT 97.780 308.190 102.940 308.360 ;
        RECT 98.180 308.080 102.940 308.190 ;
        RECT 94.360 305.170 97.240 305.560 ;
        RECT 94.360 305.120 98.310 305.170 ;
        RECT 94.360 305.070 102.110 305.120 ;
        RECT 94.360 304.900 102.270 305.070 ;
        RECT 94.360 304.830 102.110 304.900 ;
        RECT 94.360 304.720 98.310 304.830 ;
        RECT 81.610 304.000 82.880 304.390 ;
        RECT 92.750 301.630 93.120 304.550 ;
        RECT 94.360 304.080 95.410 304.720 ;
        RECT 96.900 304.690 98.310 304.720 ;
        RECT 102.530 301.900 102.940 308.080 ;
        RECT 213.630 302.480 226.860 304.490 ;
        RECT 233.600 302.480 246.830 304.490 ;
        RECT 253.710 302.480 266.940 304.490 ;
        RECT 273.820 302.480 287.050 304.490 ;
        RECT 287.390 301.940 287.820 309.330 ;
        RECT 101.720 301.840 102.940 301.900 ;
        RECT 226.290 301.850 227.610 301.940 ;
        RECT 246.260 301.850 247.580 301.940 ;
        RECT 266.370 301.850 267.690 301.940 ;
        RECT 286.480 301.850 287.820 301.940 ;
        RECT 98.100 301.780 102.940 301.840 ;
        RECT 212.280 301.790 287.820 301.850 ;
        RECT 78.900 301.580 80.010 301.610 ;
        RECT 92.030 301.600 93.140 301.630 ;
        RECT 97.780 301.610 102.940 301.780 ;
        RECT 211.830 301.620 287.820 301.790 ;
        RECT 5.290 301.530 13.530 301.570 ;
        RECT 25.760 301.550 26.870 301.580 ;
        RECT 4.750 301.360 13.530 301.530 ;
        RECT 18.630 301.510 26.870 301.550 ;
        RECT 32.000 301.540 40.240 301.580 ;
        RECT 45.230 301.540 53.470 301.580 ;
        RECT 65.630 301.550 66.740 301.580 ;
        RECT 5.290 301.310 13.530 301.360 ;
        RECT 18.090 301.340 26.870 301.510 ;
        RECT 31.460 301.370 40.240 301.540 ;
        RECT 44.690 301.370 53.470 301.540 ;
        RECT 58.500 301.510 66.740 301.550 ;
        RECT 71.770 301.540 80.010 301.580 ;
        RECT 84.900 301.560 93.140 301.600 ;
        RECT 12.420 301.250 13.530 301.310 ;
        RECT 18.630 301.290 26.870 301.340 ;
        RECT 32.000 301.320 40.240 301.370 ;
        RECT 45.230 301.320 53.470 301.370 ;
        RECT 57.960 301.340 66.740 301.510 ;
        RECT 71.230 301.370 80.010 301.540 ;
        RECT 84.360 301.390 93.140 301.560 ;
        RECT 98.100 301.550 102.940 301.610 ;
        RECT 212.280 301.600 287.820 301.620 ;
        RECT 212.280 301.590 287.800 301.600 ;
        RECT 212.280 301.580 227.610 301.590 ;
        RECT 232.250 301.580 247.580 301.590 ;
        RECT 252.360 301.580 267.690 301.590 ;
        RECT 272.470 301.580 287.800 301.590 ;
        RECT 226.290 301.560 227.610 301.580 ;
        RECT 246.260 301.560 247.580 301.580 ;
        RECT 266.370 301.560 267.690 301.580 ;
        RECT 286.480 301.560 287.800 301.580 ;
        RECT 102.530 301.520 102.940 301.550 ;
        RECT 25.760 301.230 26.870 301.290 ;
        RECT 39.130 301.260 40.240 301.320 ;
        RECT 52.360 301.260 53.470 301.320 ;
        RECT 58.500 301.290 66.740 301.340 ;
        RECT 71.770 301.320 80.010 301.370 ;
        RECT 84.900 301.340 93.140 301.390 ;
        RECT 65.630 301.230 66.740 301.290 ;
        RECT 78.900 301.260 80.010 301.320 ;
        RECT 92.030 301.280 93.140 301.340 ;
        RECT 91.200 298.500 93.400 299.010 ;
        RECT 4.720 297.450 12.880 298.470 ;
        RECT 18.060 297.430 26.220 298.450 ;
        RECT 31.430 297.460 39.590 298.480 ;
        RECT 44.660 297.460 52.820 298.480 ;
        RECT 57.930 297.430 66.090 298.450 ;
        RECT 71.200 297.460 79.360 298.480 ;
        RECT 84.330 297.710 93.400 298.500 ;
        RECT 84.330 297.480 92.490 297.710 ;
        RECT 96.820 297.280 103.000 298.630 ;
        RECT 227.220 295.300 227.490 301.560 ;
        RECT 247.190 295.300 247.460 301.560 ;
        RECT 267.300 295.300 267.570 301.560 ;
        RECT 287.210 300.850 287.680 301.560 ;
        RECT 287.410 295.300 287.680 300.850 ;
        RECT 226.470 295.270 227.790 295.300 ;
        RECT 246.440 295.270 247.760 295.300 ;
        RECT 266.550 295.270 267.870 295.300 ;
        RECT 286.660 295.270 287.980 295.300 ;
        RECT 212.520 295.210 227.790 295.270 ;
        RECT 232.490 295.210 247.760 295.270 ;
        RECT 252.600 295.210 267.870 295.270 ;
        RECT 272.710 295.210 287.980 295.270 ;
        RECT 211.830 295.040 227.790 295.210 ;
        RECT 231.800 295.040 247.760 295.210 ;
        RECT 251.910 295.040 267.870 295.210 ;
        RECT 272.020 295.040 287.980 295.210 ;
        RECT 212.520 295.000 227.790 295.040 ;
        RECT 232.490 295.000 247.760 295.040 ;
        RECT 252.600 295.000 267.870 295.040 ;
        RECT 272.710 295.000 287.980 295.040 ;
        RECT 226.470 294.920 227.790 295.000 ;
        RECT 246.440 294.920 247.760 295.000 ;
        RECT 266.550 294.920 267.870 295.000 ;
        RECT 286.660 294.920 287.980 295.000 ;
        RECT 96.680 293.550 98.090 293.600 ;
        RECT 96.680 293.470 102.070 293.550 ;
        RECT 3.730 293.280 5.330 293.390 ;
        RECT 3.730 293.270 12.370 293.280 ;
        RECT 3.640 293.220 12.370 293.270 ;
        RECT 17.070 293.260 18.670 293.370 ;
        RECT 30.440 293.290 32.040 293.400 ;
        RECT 43.670 293.290 45.270 293.400 ;
        RECT 30.440 293.280 39.080 293.290 ;
        RECT 43.670 293.280 52.310 293.290 ;
        RECT 17.070 293.250 25.710 293.260 ;
        RECT 3.640 293.050 12.570 293.220 ;
        RECT 16.980 293.200 25.710 293.250 ;
        RECT 30.350 293.230 39.080 293.280 ;
        RECT 43.580 293.230 52.310 293.280 ;
        RECT 56.940 293.260 58.540 293.370 ;
        RECT 70.210 293.290 71.810 293.400 ;
        RECT 83.340 293.310 84.940 293.420 ;
        RECT 83.340 293.300 91.980 293.310 ;
        RECT 70.210 293.280 78.850 293.290 ;
        RECT 56.940 293.250 65.580 293.260 ;
        RECT 3.640 293.020 12.370 293.050 ;
        RECT 16.980 293.030 25.910 293.200 ;
        RECT 30.350 293.060 39.280 293.230 ;
        RECT 43.580 293.060 52.510 293.230 ;
        RECT 56.850 293.200 65.580 293.250 ;
        RECT 70.120 293.230 78.850 293.280 ;
        RECT 83.250 293.250 91.980 293.300 ;
        RECT 96.680 293.300 102.130 293.470 ;
        RECT 96.680 293.260 102.070 293.300 ;
        RECT 30.350 293.030 39.080 293.060 ;
        RECT 43.580 293.030 52.310 293.060 ;
        RECT 56.850 293.030 65.780 293.200 ;
        RECT 70.120 293.060 79.050 293.230 ;
        RECT 83.250 293.080 92.180 293.250 ;
        RECT 96.680 293.120 98.090 293.260 ;
        RECT 70.120 293.030 78.850 293.060 ;
        RECT 83.250 293.050 91.980 293.080 ;
        RECT 3.640 292.780 5.330 293.020 ;
        RECT 16.980 293.000 25.710 293.030 ;
        RECT 1.110 286.490 2.770 289.370 ;
        RECT 3.640 286.780 4.100 292.780 ;
        RECT 16.980 292.760 18.670 293.000 ;
        RECT 30.350 292.790 32.040 293.030 ;
        RECT 43.580 292.790 45.270 293.030 ;
        RECT 56.850 293.000 65.580 293.030 ;
        RECT 3.640 286.670 5.260 286.780 ;
        RECT 16.980 286.760 17.440 292.760 ;
        RECT 30.350 286.790 30.810 292.790 ;
        RECT 43.580 286.790 44.040 292.790 ;
        RECT 56.850 292.760 58.540 293.000 ;
        RECT 70.120 292.790 71.810 293.030 ;
        RECT 83.250 292.810 84.940 293.050 ;
        RECT 3.640 286.640 12.390 286.670 ;
        RECT 16.980 286.650 18.600 286.760 ;
        RECT 30.350 286.680 31.970 286.790 ;
        RECT 43.580 286.680 45.200 286.790 ;
        RECT 56.850 286.760 57.310 292.760 ;
        RECT 70.120 286.790 70.580 292.790 ;
        RECT 83.250 286.810 83.710 292.810 ;
        RECT 96.760 287.020 97.100 293.120 ;
        RECT 227.220 288.730 227.490 294.920 ;
        RECT 247.190 288.730 247.460 294.920 ;
        RECT 267.300 288.730 267.570 294.920 ;
        RECT 287.410 288.730 287.680 294.920 ;
        RECT 355.040 294.780 356.120 309.080 ;
        RECT 356.460 295.780 356.740 309.610 ;
        RECT 359.820 309.000 359.990 309.160 ;
        RECT 356.440 290.940 356.820 295.780 ;
        RECT 359.770 295.000 360.050 309.000 ;
        RECT 363.050 308.980 363.330 309.610 ;
        RECT 369.600 309.560 370.530 309.610 ;
        RECT 375.760 309.720 376.060 314.090 ;
        RECT 382.360 327.540 382.650 327.700 ;
        RECT 388.920 328.280 389.850 328.330 ;
        RECT 382.360 313.480 382.640 327.540 ;
        RECT 388.920 327.390 389.300 328.280 ;
        RECT 382.430 312.980 382.600 313.480 ;
        RECT 388.930 313.290 389.210 327.390 ;
        RECT 393.610 313.570 394.690 327.870 ;
        RECT 395.030 314.160 395.310 328.400 ;
        RECT 398.390 327.790 398.560 327.950 ;
        RECT 389.010 312.980 389.180 313.290 ;
        RECT 388.960 309.760 389.850 309.810 ;
        RECT 388.920 309.720 389.850 309.760 ;
        RECT 359.720 294.780 360.050 295.000 ;
        RECT 363.040 308.820 363.330 308.980 ;
        RECT 359.720 293.790 360.020 294.780 ;
        RECT 363.040 294.760 363.320 308.820 ;
        RECT 366.400 308.770 366.570 309.160 ;
        RECT 366.340 294.990 366.620 308.770 ;
        RECT 369.600 308.670 369.980 309.560 ;
        RECT 375.760 309.510 389.850 309.720 ;
        RECT 395.010 309.790 395.310 314.160 ;
        RECT 398.340 313.790 398.620 327.790 ;
        RECT 401.620 327.770 401.900 328.400 ;
        RECT 408.170 328.350 409.100 328.400 ;
        RECT 398.290 313.570 398.620 313.790 ;
        RECT 401.610 327.610 401.900 327.770 ;
        RECT 398.290 312.580 398.590 313.570 ;
        RECT 401.610 313.550 401.890 327.610 ;
        RECT 404.970 327.560 405.140 327.950 ;
        RECT 404.910 313.780 405.190 327.560 ;
        RECT 408.170 327.460 408.550 328.350 ;
        RECT 401.680 313.050 401.850 313.550 ;
        RECT 404.910 313.340 405.230 313.780 ;
        RECT 408.180 313.360 408.460 327.460 ;
        RECT 858.170 327.420 858.340 327.840 ;
        RECT 860.750 327.420 860.920 327.840 ;
        RECT 658.760 326.185 660.200 326.355 ;
        RECT 663.660 326.145 665.100 326.315 ;
        RECT 668.250 326.175 669.690 326.345 ;
        RECT 672.790 326.155 674.230 326.325 ;
        RECT 676.220 326.165 680.060 326.335 ;
        RECT 681.990 326.165 685.350 326.335 ;
        RECT 687.440 326.165 690.800 326.335 ;
        RECT 692.750 326.185 696.110 326.355 ;
        RECT 591.830 323.470 592.180 325.630 ;
        RECT 658.850 324.375 659.440 325.955 ;
        RECT 663.750 324.335 664.340 325.915 ;
        RECT 668.340 324.365 668.930 325.945 ;
        RECT 670.660 324.700 671.340 325.780 ;
        RECT 672.880 324.345 673.470 325.925 ;
        RECT 676.780 324.850 677.730 325.885 ;
        RECT 678.420 324.355 679.370 325.935 ;
        RECT 682.080 324.435 683.010 325.885 ;
        RECT 683.540 324.435 684.790 325.935 ;
        RECT 687.530 324.435 688.460 325.885 ;
        RECT 688.990 324.435 690.240 325.935 ;
        RECT 691.280 324.570 692.030 325.670 ;
        RECT 693.580 324.455 695.550 325.955 ;
        RECT 858.170 325.950 858.340 326.370 ;
        RECT 860.750 325.950 860.920 326.370 ;
        RECT 858.170 324.480 858.340 324.900 ;
        RECT 860.750 324.480 860.920 324.900 ;
        RECT 858.170 323.010 858.340 323.430 ;
        RECT 860.750 323.010 860.920 323.430 ;
        RECT 858.170 321.540 858.340 321.960 ;
        RECT 860.750 321.540 860.920 321.960 ;
        RECT 661.400 320.305 665.240 320.475 ;
        RECT 667.220 320.315 670.580 320.485 ;
        RECT 672.660 320.325 676.020 320.495 ;
        RECT 677.980 320.325 681.340 320.495 ;
        RECT 683.330 320.325 686.690 320.495 ;
        RECT 689.150 320.305 691.550 320.475 ;
        RECT 661.960 318.990 662.910 320.025 ;
        RECT 663.600 318.495 664.550 320.075 ;
        RECT 667.310 318.585 668.240 320.035 ;
        RECT 668.770 318.585 670.020 320.085 ;
        RECT 671.050 319.500 672.200 320.230 ;
        RECT 672.750 318.595 673.680 320.045 ;
        RECT 674.210 318.595 675.460 320.095 ;
        RECT 678.810 318.595 680.780 320.095 ;
        RECT 681.830 319.140 682.660 320.020 ;
        RECT 683.420 318.595 684.350 320.045 ;
        RECT 684.880 318.595 686.130 320.095 ;
        RECT 690.265 318.495 690.820 320.075 ;
        RECT 691.930 319.730 693.110 320.460 ;
        RECT 693.550 320.305 695.950 320.475 ;
        RECT 694.665 318.495 695.220 320.075 ;
        RECT 858.170 320.070 858.340 320.490 ;
        RECT 860.750 320.070 860.920 320.490 ;
        RECT 864.740 320.450 864.910 320.870 ;
        RECT 867.320 320.450 867.490 320.870 ;
        RECT 868.680 320.440 868.850 320.860 ;
        RECT 871.260 320.440 871.430 320.860 ;
        RECT 858.170 318.600 858.340 319.020 ;
        RECT 860.750 318.600 860.920 319.020 ;
        RECT 864.740 318.980 864.910 319.400 ;
        RECT 867.320 318.980 867.490 319.400 ;
        RECT 868.680 318.970 868.850 319.390 ;
        RECT 871.260 318.970 871.430 319.390 ;
        RECT 858.170 317.130 858.340 317.550 ;
        RECT 860.750 317.130 860.920 317.550 ;
        RECT 864.740 317.510 864.910 317.930 ;
        RECT 867.320 317.510 867.490 317.930 ;
        RECT 868.680 317.500 868.850 317.920 ;
        RECT 871.260 317.500 871.430 317.920 ;
        RECT 858.170 315.660 858.340 316.080 ;
        RECT 860.750 315.660 860.920 316.080 ;
        RECT 864.740 316.040 864.910 316.460 ;
        RECT 867.320 316.040 867.490 316.460 ;
        RECT 868.680 316.030 868.850 316.450 ;
        RECT 871.260 316.030 871.430 316.450 ;
        RECT 871.830 315.090 872.310 319.010 ;
        RECT 404.930 312.600 405.230 313.340 ;
        RECT 408.260 313.050 408.430 313.360 ;
        RECT 404.930 312.580 405.720 312.600 ;
        RECT 398.290 312.270 405.720 312.580 ;
        RECT 595.220 312.525 596.660 312.695 ;
        RECT 398.290 312.240 398.590 312.270 ;
        RECT 404.930 312.230 405.230 312.270 ;
        RECT 595.980 310.715 596.570 312.295 ;
        RECT 601.030 311.830 601.770 314.690 ;
        RECT 602.480 313.880 602.650 314.300 ;
        RECT 604.060 313.880 604.230 314.300 ;
        RECT 605.640 313.880 605.810 314.300 ;
        RECT 607.000 313.890 607.170 314.310 ;
        RECT 608.580 313.890 608.750 314.310 ;
        RECT 610.160 313.890 610.330 314.310 ;
        RECT 611.520 313.890 611.690 314.310 ;
        RECT 613.100 313.890 613.270 314.310 ;
        RECT 614.680 313.890 614.850 314.310 ;
        RECT 615.950 313.870 616.120 314.290 ;
        RECT 617.530 313.870 617.700 314.290 ;
        RECT 619.110 313.870 619.280 314.290 ;
        RECT 620.330 313.880 620.500 314.300 ;
        RECT 621.910 313.880 622.080 314.300 ;
        RECT 623.490 313.880 623.660 314.300 ;
        RECT 624.650 313.870 624.820 314.290 ;
        RECT 626.230 313.870 626.400 314.290 ;
        RECT 627.810 313.870 627.980 314.290 ;
        RECT 602.480 312.410 602.650 312.830 ;
        RECT 604.060 312.410 604.230 312.830 ;
        RECT 605.640 312.410 605.810 312.830 ;
        RECT 607.000 312.420 607.170 312.840 ;
        RECT 608.580 312.420 608.750 312.840 ;
        RECT 610.160 312.420 610.330 312.840 ;
        RECT 611.520 312.420 611.690 312.840 ;
        RECT 613.100 312.420 613.270 312.840 ;
        RECT 614.680 312.420 614.850 312.840 ;
        RECT 615.950 312.400 616.120 312.820 ;
        RECT 617.530 312.400 617.700 312.820 ;
        RECT 619.110 312.400 619.280 312.820 ;
        RECT 620.330 312.410 620.500 312.830 ;
        RECT 621.910 312.410 622.080 312.830 ;
        RECT 623.490 312.410 623.660 312.830 ;
        RECT 624.650 312.400 624.820 312.820 ;
        RECT 626.230 312.400 626.400 312.820 ;
        RECT 627.810 312.400 627.980 312.820 ;
        RECT 628.730 311.660 629.600 314.980 ;
        RECT 858.170 314.190 858.340 314.610 ;
        RECT 860.750 314.190 860.920 314.610 ;
        RECT 864.740 314.570 864.910 314.990 ;
        RECT 867.320 314.570 867.490 314.990 ;
        RECT 868.680 314.560 868.850 314.980 ;
        RECT 871.260 314.560 871.430 314.980 ;
        RECT 635.110 312.975 636.550 313.145 ;
        RECT 639.300 313.065 640.740 313.235 ;
        RECT 643.400 313.045 644.840 313.215 ;
        RECT 635.200 311.165 635.790 312.745 ;
        RECT 639.390 311.255 639.980 312.835 ;
        RECT 643.490 311.235 644.080 312.815 ;
        RECT 645.240 311.610 645.880 312.920 ;
        RECT 408.210 309.830 409.100 309.880 ;
        RECT 408.170 309.790 409.100 309.830 ;
        RECT 395.010 309.580 409.100 309.790 ;
        RECT 363.110 294.260 363.280 294.760 ;
        RECT 366.340 294.550 366.660 294.990 ;
        RECT 369.610 294.570 369.890 308.670 ;
        RECT 374.360 294.680 375.440 308.980 ;
        RECT 375.780 295.680 376.060 309.510 ;
        RECT 382.370 308.880 382.650 309.510 ;
        RECT 382.360 308.720 382.650 308.880 ;
        RECT 388.920 309.460 389.850 309.510 ;
        RECT 366.360 293.810 366.660 294.550 ;
        RECT 369.690 294.260 369.860 294.570 ;
        RECT 366.360 293.790 367.150 293.810 ;
        RECT 359.720 293.480 367.150 293.790 ;
        RECT 359.720 293.450 360.020 293.480 ;
        RECT 366.360 293.440 366.660 293.480 ;
        RECT 369.640 290.980 370.530 291.030 ;
        RECT 369.600 290.940 370.530 290.980 ;
        RECT 356.440 290.730 370.530 290.940 ;
        RECT 356.440 290.440 356.820 290.730 ;
        RECT 226.320 288.660 227.640 288.730 ;
        RECT 246.290 288.660 247.610 288.730 ;
        RECT 266.400 288.660 267.720 288.730 ;
        RECT 286.510 288.660 287.830 288.730 ;
        RECT 212.510 288.630 227.640 288.660 ;
        RECT 232.480 288.630 247.610 288.660 ;
        RECT 252.590 288.630 267.720 288.660 ;
        RECT 272.700 288.630 287.830 288.660 ;
        RECT 211.830 288.460 227.640 288.630 ;
        RECT 231.800 288.460 247.610 288.630 ;
        RECT 251.910 288.460 267.720 288.630 ;
        RECT 272.020 288.460 287.830 288.630 ;
        RECT 212.510 288.390 227.640 288.460 ;
        RECT 232.480 288.390 247.610 288.460 ;
        RECT 252.590 288.390 267.720 288.460 ;
        RECT 272.700 288.390 287.830 288.460 ;
        RECT 226.320 288.350 227.640 288.390 ;
        RECT 246.290 288.350 247.610 288.390 ;
        RECT 266.400 288.350 267.720 288.390 ;
        RECT 286.510 288.350 287.830 288.390 ;
        RECT 227.220 288.340 227.490 288.350 ;
        RECT 247.190 288.340 247.460 288.350 ;
        RECT 267.300 288.340 267.570 288.350 ;
        RECT 287.410 288.340 287.680 288.350 ;
        RECT 96.760 286.970 98.190 287.020 ;
        RECT 96.760 286.890 102.110 286.970 ;
        RECT 30.350 286.650 39.100 286.680 ;
        RECT 43.580 286.650 52.330 286.680 ;
        RECT 56.850 286.650 58.470 286.760 ;
        RECT 70.120 286.680 71.740 286.790 ;
        RECT 83.250 286.700 84.870 286.810 ;
        RECT 96.760 286.720 102.130 286.890 ;
        RECT 70.120 286.650 78.870 286.680 ;
        RECT 83.250 286.670 92.000 286.700 ;
        RECT 96.760 286.680 102.110 286.720 ;
        RECT 3.640 286.490 12.570 286.640 ;
        RECT 1.110 286.470 12.570 286.490 ;
        RECT 16.980 286.620 25.730 286.650 ;
        RECT 1.110 286.410 12.390 286.470 ;
        RECT 16.980 286.450 25.910 286.620 ;
        RECT 30.350 286.480 39.280 286.650 ;
        RECT 43.580 286.480 52.510 286.650 ;
        RECT 56.850 286.620 65.600 286.650 ;
        RECT 1.110 286.170 5.260 286.410 ;
        RECT 16.980 286.390 25.730 286.450 ;
        RECT 30.350 286.420 39.100 286.480 ;
        RECT 43.580 286.420 52.330 286.480 ;
        RECT 56.850 286.450 65.780 286.620 ;
        RECT 70.120 286.480 79.050 286.650 ;
        RECT 83.250 286.500 92.180 286.670 ;
        RECT 96.760 286.540 98.190 286.680 ;
        RECT 1.110 285.920 4.270 286.170 ;
        RECT 16.980 286.150 18.600 286.390 ;
        RECT 30.350 286.180 31.970 286.420 ;
        RECT 43.580 286.180 45.200 286.420 ;
        RECT 56.850 286.390 65.600 286.450 ;
        RECT 70.120 286.420 78.870 286.480 ;
        RECT 83.250 286.440 92.000 286.500 ;
        RECT 1.110 282.760 2.770 285.920 ;
        RECT 3.640 280.210 4.100 285.920 ;
        RECT 3.610 280.100 5.210 280.210 ;
        RECT 16.980 280.190 17.440 286.150 ;
        RECT 30.350 280.220 30.810 286.180 ;
        RECT 43.580 280.220 44.040 286.180 ;
        RECT 56.850 286.150 58.470 286.390 ;
        RECT 70.120 286.180 71.740 286.420 ;
        RECT 83.250 286.200 84.870 286.440 ;
        RECT 3.610 280.060 12.440 280.100 ;
        RECT 16.950 280.080 18.550 280.190 ;
        RECT 30.320 280.110 31.920 280.220 ;
        RECT 43.550 280.110 45.150 280.220 ;
        RECT 56.850 280.190 57.310 286.150 ;
        RECT 70.120 280.220 70.580 286.180 ;
        RECT 83.250 280.240 83.710 286.200 ;
        RECT 96.760 280.380 97.100 286.540 ;
        RECT 213.390 280.530 226.620 282.540 ;
        RECT 233.430 280.520 246.660 282.530 ;
        RECT 253.490 280.520 266.720 282.530 ;
        RECT 273.540 280.520 286.770 282.530 ;
        RECT 96.740 280.310 102.050 280.380 ;
        RECT 3.610 279.890 12.570 280.060 ;
        RECT 16.950 280.040 25.780 280.080 ;
        RECT 30.320 280.070 39.150 280.110 ;
        RECT 43.550 280.070 52.380 280.110 ;
        RECT 56.820 280.080 58.420 280.190 ;
        RECT 70.090 280.110 71.690 280.220 ;
        RECT 83.220 280.130 84.820 280.240 ;
        RECT 96.740 280.140 102.130 280.310 ;
        RECT 3.610 279.840 12.440 279.890 ;
        RECT 16.950 279.870 25.910 280.040 ;
        RECT 30.320 279.900 39.280 280.070 ;
        RECT 43.550 279.900 52.510 280.070 ;
        RECT 56.820 280.040 65.650 280.080 ;
        RECT 70.090 280.070 78.920 280.110 ;
        RECT 83.220 280.090 92.050 280.130 ;
        RECT 96.740 280.090 102.050 280.140 ;
        RECT 3.610 279.600 5.210 279.840 ;
        RECT 16.950 279.820 25.780 279.870 ;
        RECT 30.320 279.850 39.150 279.900 ;
        RECT 43.550 279.850 52.380 279.900 ;
        RECT 56.820 279.870 65.780 280.040 ;
        RECT 70.090 279.900 79.050 280.070 ;
        RECT 83.220 279.920 92.180 280.090 ;
        RECT 3.640 273.770 4.100 279.600 ;
        RECT 16.950 279.580 18.550 279.820 ;
        RECT 30.320 279.610 31.920 279.850 ;
        RECT 43.550 279.610 45.150 279.850 ;
        RECT 56.820 279.820 65.650 279.870 ;
        RECT 70.090 279.850 78.920 279.900 ;
        RECT 83.220 279.870 92.050 279.920 ;
        RECT 96.740 279.900 98.150 280.090 ;
        RECT 226.050 279.920 227.370 279.990 ;
        RECT 246.090 279.920 247.410 279.980 ;
        RECT 266.150 279.920 267.470 279.980 ;
        RECT 286.200 279.920 287.520 279.980 ;
        RECT 3.560 273.530 5.160 273.770 ;
        RECT 15.290 273.710 16.380 274.010 ;
        RECT 16.980 273.750 17.440 279.580 ;
        RECT 28.460 273.760 29.640 274.180 ;
        RECT 30.350 273.780 30.810 279.610 ;
        RECT 41.760 273.840 42.770 274.560 ;
        RECT 43.580 273.840 44.040 279.610 ;
        RECT 56.820 279.580 58.420 279.820 ;
        RECT 70.090 279.610 71.690 279.850 ;
        RECT 83.220 279.630 84.820 279.870 ;
        RECT 41.760 273.780 44.110 273.840 ;
        RECT 55.140 273.800 56.230 274.140 ;
        RECT 56.850 273.800 57.310 279.580 ;
        RECT 30.270 273.760 31.870 273.780 ;
        RECT 16.900 273.710 18.500 273.750 ;
        RECT 3.560 273.270 12.680 273.530 ;
        RECT 15.290 273.510 18.500 273.710 ;
        RECT 28.460 273.540 31.870 273.760 ;
        RECT 41.760 273.540 45.100 273.780 ;
        RECT 3.560 273.160 5.160 273.270 ;
        RECT 15.290 273.250 26.020 273.510 ;
        RECT 28.460 273.280 39.390 273.540 ;
        RECT 41.760 273.280 52.620 273.540 ;
        RECT 55.140 273.510 59.600 273.800 ;
        RECT 68.390 273.670 69.230 274.300 ;
        RECT 70.120 273.780 70.580 279.610 ;
        RECT 81.470 273.840 82.740 274.010 ;
        RECT 83.250 273.840 83.710 279.630 ;
        RECT 94.220 274.220 95.270 274.470 ;
        RECT 96.760 274.220 97.100 279.900 ;
        RECT 211.960 279.840 287.520 279.920 ;
        RECT 211.590 279.670 287.520 279.840 ;
        RECT 211.960 279.660 287.520 279.670 ;
        RECT 212.040 279.630 227.370 279.660 ;
        RECT 226.050 279.610 227.370 279.630 ;
        RECT 232.080 279.620 247.410 279.660 ;
        RECT 252.140 279.620 267.470 279.660 ;
        RECT 272.190 279.620 287.520 279.660 ;
        RECT 70.040 273.670 71.640 273.780 ;
        RECT 68.390 273.540 72.300 273.670 ;
        RECT 81.470 273.560 85.170 273.840 ;
        RECT 94.220 273.830 97.100 274.220 ;
        RECT 210.780 276.610 212.210 276.680 ;
        RECT 210.780 276.550 226.460 276.610 ;
        RECT 210.780 276.380 226.490 276.550 ;
        RECT 210.780 276.340 226.460 276.380 ;
        RECT 210.780 276.300 212.210 276.340 ;
        RECT 94.220 273.780 98.170 273.830 ;
        RECT 94.220 273.730 101.970 273.780 ;
        RECT 94.220 273.560 102.130 273.730 ;
        RECT 15.290 273.140 18.500 273.250 ;
        RECT 28.460 273.210 31.870 273.280 ;
        RECT 15.290 273.000 17.520 273.140 ;
        RECT 15.290 272.240 16.380 273.000 ;
        RECT 28.460 272.370 29.640 273.210 ;
        RECT 30.270 273.170 31.870 273.210 ;
        RECT 41.760 273.210 45.100 273.280 ;
        RECT 41.760 272.120 42.770 273.210 ;
        RECT 43.500 273.170 45.100 273.210 ;
        RECT 55.140 273.250 65.890 273.510 ;
        RECT 68.390 273.280 79.160 273.540 ;
        RECT 81.470 273.300 92.290 273.560 ;
        RECT 94.220 273.490 101.970 273.560 ;
        RECT 94.220 273.380 98.170 273.490 ;
        RECT 55.140 273.210 59.600 273.250 ;
        RECT 55.140 271.950 56.230 273.210 ;
        RECT 56.770 273.140 58.370 273.210 ;
        RECT 68.390 273.080 72.300 273.280 ;
        RECT 68.390 272.160 69.230 273.080 ;
        RECT 81.470 273.050 85.170 273.300 ;
        RECT 81.470 272.660 82.740 273.050 ;
        RECT 94.220 272.740 95.270 273.380 ;
        RECT 96.760 273.350 98.170 273.380 ;
        RECT 210.780 270.070 211.190 276.300 ;
        RECT 226.980 273.350 227.250 279.610 ;
        RECT 246.090 279.600 247.410 279.620 ;
        RECT 266.150 279.600 267.470 279.620 ;
        RECT 286.200 279.600 287.520 279.620 ;
        RECT 230.820 276.600 232.250 276.670 ;
        RECT 230.820 276.540 246.500 276.600 ;
        RECT 230.820 276.370 246.530 276.540 ;
        RECT 230.820 276.330 246.500 276.370 ;
        RECT 230.820 276.290 232.250 276.330 ;
        RECT 226.230 273.320 227.550 273.350 ;
        RECT 212.280 273.260 227.550 273.320 ;
        RECT 211.590 273.090 227.550 273.260 ;
        RECT 212.280 273.050 227.550 273.090 ;
        RECT 226.230 272.970 227.550 273.050 ;
        RECT 210.760 270.030 212.360 270.070 ;
        RECT 210.760 269.760 226.500 270.030 ;
        RECT 210.760 269.690 212.360 269.760 ;
        RECT 4.720 265.620 12.880 266.640 ;
        RECT 18.060 265.600 26.220 266.620 ;
        RECT 31.430 265.630 39.590 266.650 ;
        RECT 44.660 265.630 52.820 266.650 ;
        RECT 57.930 265.600 66.090 266.620 ;
        RECT 71.200 265.630 79.360 266.650 ;
        RECT 84.330 265.650 92.490 266.670 ;
        RECT 96.820 265.450 103.000 266.800 ;
        RECT 11.800 265.030 102.640 265.240 ;
        RECT 11.800 264.990 102.760 265.030 ;
        RECT 11.800 264.770 102.800 264.990 ;
        RECT 4.540 264.450 102.800 264.770 ;
        RECT 11.800 264.390 102.800 264.450 ;
        RECT 3.730 261.450 5.330 261.560 ;
        RECT 3.730 261.440 12.370 261.450 ;
        RECT 3.640 261.390 12.370 261.440 ;
        RECT 3.640 261.220 12.570 261.390 ;
        RECT 3.640 261.190 12.370 261.220 ;
        RECT 3.640 260.950 5.330 261.190 ;
        RECT 3.640 254.950 4.100 260.950 ;
        RECT 13.050 258.140 13.390 264.390 ;
        RECT 17.070 261.430 18.670 261.540 ;
        RECT 17.070 261.420 25.710 261.430 ;
        RECT 4.780 258.100 13.390 258.140 ;
        RECT 4.610 257.930 13.390 258.100 ;
        RECT 4.780 257.880 13.390 257.930 ;
        RECT 11.950 257.870 13.390 257.880 ;
        RECT 3.640 254.840 5.260 254.950 ;
        RECT 3.640 254.810 12.390 254.840 ;
        RECT 3.640 254.640 12.570 254.810 ;
        RECT 3.640 254.580 12.390 254.640 ;
        RECT 3.640 254.340 5.260 254.580 ;
        RECT 3.640 248.380 4.100 254.340 ;
        RECT 13.050 251.580 13.390 257.870 ;
        RECT 12.010 251.570 13.390 251.580 ;
        RECT 4.850 251.520 13.390 251.570 ;
        RECT 4.610 251.350 13.390 251.520 ;
        RECT 4.850 251.310 13.390 251.350 ;
        RECT 3.610 248.270 5.210 248.380 ;
        RECT 3.610 248.230 12.440 248.270 ;
        RECT 3.610 248.060 12.570 248.230 ;
        RECT 3.610 248.010 12.440 248.060 ;
        RECT 3.610 247.770 5.210 248.010 ;
        RECT 3.640 241.940 4.100 247.770 ;
        RECT 13.050 244.990 13.390 251.310 ;
        RECT 16.980 261.370 25.710 261.420 ;
        RECT 16.980 261.200 25.910 261.370 ;
        RECT 16.980 261.170 25.710 261.200 ;
        RECT 16.980 260.930 18.670 261.170 ;
        RECT 16.980 254.930 17.440 260.930 ;
        RECT 26.390 258.120 26.730 264.390 ;
        RECT 30.440 261.460 32.040 261.570 ;
        RECT 30.440 261.450 39.080 261.460 ;
        RECT 18.120 258.080 26.730 258.120 ;
        RECT 17.950 257.910 26.730 258.080 ;
        RECT 18.120 257.860 26.730 257.910 ;
        RECT 25.290 257.850 26.730 257.860 ;
        RECT 16.980 254.820 18.600 254.930 ;
        RECT 16.980 254.790 25.730 254.820 ;
        RECT 16.980 254.620 25.910 254.790 ;
        RECT 16.980 254.560 25.730 254.620 ;
        RECT 16.980 254.320 18.600 254.560 ;
        RECT 16.980 248.360 17.440 254.320 ;
        RECT 26.390 251.560 26.730 257.850 ;
        RECT 25.350 251.550 26.730 251.560 ;
        RECT 18.190 251.500 26.730 251.550 ;
        RECT 17.950 251.330 26.730 251.500 ;
        RECT 18.190 251.290 26.730 251.330 ;
        RECT 16.950 248.250 18.550 248.360 ;
        RECT 16.950 248.210 25.780 248.250 ;
        RECT 16.950 248.040 25.910 248.210 ;
        RECT 16.950 247.990 25.780 248.040 ;
        RECT 16.950 247.750 18.550 247.990 ;
        RECT 11.960 244.980 13.390 244.990 ;
        RECT 4.970 244.940 13.390 244.980 ;
        RECT 4.610 244.770 13.390 244.940 ;
        RECT 4.970 244.720 13.390 244.770 ;
        RECT 3.560 241.700 5.160 241.940 ;
        RECT 3.560 241.440 12.680 241.700 ;
        RECT 13.050 241.560 13.390 244.720 ;
        RECT 3.560 241.330 5.160 241.440 ;
        RECT 13.000 241.350 13.390 241.560 ;
        RECT 15.290 241.880 16.380 242.180 ;
        RECT 16.980 241.920 17.440 247.750 ;
        RECT 26.390 244.970 26.730 251.290 ;
        RECT 30.350 261.400 39.080 261.450 ;
        RECT 30.350 261.230 39.280 261.400 ;
        RECT 30.350 261.200 39.080 261.230 ;
        RECT 30.350 260.960 32.040 261.200 ;
        RECT 30.350 254.960 30.810 260.960 ;
        RECT 39.760 258.150 40.100 264.390 ;
        RECT 43.670 261.460 45.270 261.570 ;
        RECT 43.670 261.450 52.310 261.460 ;
        RECT 31.490 258.110 40.100 258.150 ;
        RECT 31.320 257.940 40.100 258.110 ;
        RECT 31.490 257.890 40.100 257.940 ;
        RECT 38.660 257.880 40.100 257.890 ;
        RECT 30.350 254.850 31.970 254.960 ;
        RECT 30.350 254.820 39.100 254.850 ;
        RECT 30.350 254.650 39.280 254.820 ;
        RECT 30.350 254.590 39.100 254.650 ;
        RECT 30.350 254.350 31.970 254.590 ;
        RECT 30.350 248.390 30.810 254.350 ;
        RECT 39.760 251.590 40.100 257.880 ;
        RECT 38.720 251.580 40.100 251.590 ;
        RECT 31.560 251.530 40.100 251.580 ;
        RECT 31.320 251.360 40.100 251.530 ;
        RECT 31.560 251.320 40.100 251.360 ;
        RECT 30.320 248.280 31.920 248.390 ;
        RECT 30.320 248.240 39.150 248.280 ;
        RECT 30.320 248.070 39.280 248.240 ;
        RECT 30.320 248.020 39.150 248.070 ;
        RECT 30.320 247.780 31.920 248.020 ;
        RECT 25.300 244.960 26.730 244.970 ;
        RECT 18.310 244.920 26.730 244.960 ;
        RECT 17.950 244.750 26.730 244.920 ;
        RECT 18.310 244.700 26.730 244.750 ;
        RECT 16.900 241.880 18.500 241.920 ;
        RECT 15.290 241.680 18.500 241.880 ;
        RECT 15.290 241.420 26.020 241.680 ;
        RECT 26.390 241.540 26.730 244.700 ;
        RECT -46.120 236.660 -32.630 239.280 ;
        RECT 13.000 238.430 13.370 241.350 ;
        RECT 15.290 241.310 18.500 241.420 ;
        RECT 26.340 241.330 26.730 241.540 ;
        RECT 28.460 241.930 29.640 242.350 ;
        RECT 30.350 241.950 30.810 247.780 ;
        RECT 39.760 245.000 40.100 251.320 ;
        RECT 43.580 261.400 52.310 261.450 ;
        RECT 43.580 261.230 52.510 261.400 ;
        RECT 43.580 261.200 52.310 261.230 ;
        RECT 43.580 260.960 45.270 261.200 ;
        RECT 43.580 254.960 44.040 260.960 ;
        RECT 52.990 258.150 53.330 264.390 ;
        RECT 56.940 261.430 58.540 261.540 ;
        RECT 56.940 261.420 65.580 261.430 ;
        RECT 44.720 258.110 53.330 258.150 ;
        RECT 44.550 257.940 53.330 258.110 ;
        RECT 44.720 257.890 53.330 257.940 ;
        RECT 51.890 257.880 53.330 257.890 ;
        RECT 43.580 254.850 45.200 254.960 ;
        RECT 43.580 254.820 52.330 254.850 ;
        RECT 43.580 254.650 52.510 254.820 ;
        RECT 43.580 254.590 52.330 254.650 ;
        RECT 43.580 254.350 45.200 254.590 ;
        RECT 43.580 248.390 44.040 254.350 ;
        RECT 52.990 251.590 53.330 257.880 ;
        RECT 51.950 251.580 53.330 251.590 ;
        RECT 44.790 251.530 53.330 251.580 ;
        RECT 44.550 251.360 53.330 251.530 ;
        RECT 44.790 251.320 53.330 251.360 ;
        RECT 43.550 248.280 45.150 248.390 ;
        RECT 43.550 248.240 52.380 248.280 ;
        RECT 43.550 248.070 52.510 248.240 ;
        RECT 43.550 248.020 52.380 248.070 ;
        RECT 43.550 247.780 45.150 248.020 ;
        RECT 38.670 244.990 40.100 245.000 ;
        RECT 31.680 244.950 40.100 244.990 ;
        RECT 31.320 244.780 40.100 244.950 ;
        RECT 31.680 244.730 40.100 244.780 ;
        RECT 30.270 241.930 31.870 241.950 ;
        RECT 28.460 241.710 31.870 241.930 ;
        RECT 28.460 241.450 39.390 241.710 ;
        RECT 39.760 241.570 40.100 244.730 ;
        RECT 28.460 241.380 31.870 241.450 ;
        RECT 15.290 241.170 17.520 241.310 ;
        RECT 15.290 240.410 16.380 241.170 ;
        RECT 12.280 238.400 13.390 238.430 ;
        RECT 26.340 238.410 26.710 241.330 ;
        RECT 28.460 240.540 29.640 241.380 ;
        RECT 30.270 241.340 31.870 241.380 ;
        RECT 39.710 241.360 40.100 241.570 ;
        RECT 41.760 242.010 42.770 242.730 ;
        RECT 43.580 242.010 44.040 247.780 ;
        RECT 52.990 245.000 53.330 251.320 ;
        RECT 56.850 261.370 65.580 261.420 ;
        RECT 56.850 261.200 65.780 261.370 ;
        RECT 56.850 261.170 65.580 261.200 ;
        RECT 56.850 260.930 58.540 261.170 ;
        RECT 56.850 254.930 57.310 260.930 ;
        RECT 66.260 258.120 66.600 264.390 ;
        RECT 70.210 261.460 71.810 261.570 ;
        RECT 70.210 261.450 78.850 261.460 ;
        RECT 57.990 258.080 66.600 258.120 ;
        RECT 57.820 257.910 66.600 258.080 ;
        RECT 57.990 257.860 66.600 257.910 ;
        RECT 65.160 257.850 66.600 257.860 ;
        RECT 56.850 254.820 58.470 254.930 ;
        RECT 56.850 254.790 65.600 254.820 ;
        RECT 56.850 254.620 65.780 254.790 ;
        RECT 56.850 254.560 65.600 254.620 ;
        RECT 56.850 254.320 58.470 254.560 ;
        RECT 56.850 248.360 57.310 254.320 ;
        RECT 66.260 251.560 66.600 257.850 ;
        RECT 65.220 251.550 66.600 251.560 ;
        RECT 58.060 251.500 66.600 251.550 ;
        RECT 57.820 251.330 66.600 251.500 ;
        RECT 58.060 251.290 66.600 251.330 ;
        RECT 56.820 248.250 58.420 248.360 ;
        RECT 56.820 248.210 65.650 248.250 ;
        RECT 56.820 248.040 65.780 248.210 ;
        RECT 56.820 247.990 65.650 248.040 ;
        RECT 56.820 247.750 58.420 247.990 ;
        RECT 51.900 244.990 53.330 245.000 ;
        RECT 44.910 244.950 53.330 244.990 ;
        RECT 44.550 244.780 53.330 244.950 ;
        RECT 44.910 244.730 53.330 244.780 ;
        RECT 41.760 241.950 44.110 242.010 ;
        RECT 41.760 241.710 45.100 241.950 ;
        RECT 41.760 241.450 52.620 241.710 ;
        RECT 52.990 241.570 53.330 244.730 ;
        RECT 41.760 241.380 45.100 241.450 ;
        RECT 39.710 238.440 40.080 241.360 ;
        RECT 41.760 240.290 42.770 241.380 ;
        RECT 43.500 241.340 45.100 241.380 ;
        RECT 52.940 241.360 53.330 241.570 ;
        RECT 55.140 241.970 56.230 242.310 ;
        RECT 56.850 241.970 57.310 247.750 ;
        RECT 66.260 244.970 66.600 251.290 ;
        RECT 70.120 261.400 78.850 261.450 ;
        RECT 70.120 261.230 79.050 261.400 ;
        RECT 70.120 261.200 78.850 261.230 ;
        RECT 70.120 260.960 71.810 261.200 ;
        RECT 70.120 254.960 70.580 260.960 ;
        RECT 79.530 258.150 79.870 264.390 ;
        RECT 83.340 261.480 84.940 261.590 ;
        RECT 83.340 261.470 91.980 261.480 ;
        RECT 71.260 258.110 79.870 258.150 ;
        RECT 71.090 257.940 79.870 258.110 ;
        RECT 71.260 257.890 79.870 257.940 ;
        RECT 78.430 257.880 79.870 257.890 ;
        RECT 70.120 254.850 71.740 254.960 ;
        RECT 70.120 254.820 78.870 254.850 ;
        RECT 70.120 254.650 79.050 254.820 ;
        RECT 70.120 254.590 78.870 254.650 ;
        RECT 70.120 254.350 71.740 254.590 ;
        RECT 70.120 248.390 70.580 254.350 ;
        RECT 79.530 251.590 79.870 257.880 ;
        RECT 78.490 251.580 79.870 251.590 ;
        RECT 71.330 251.530 79.870 251.580 ;
        RECT 71.090 251.360 79.870 251.530 ;
        RECT 71.330 251.320 79.870 251.360 ;
        RECT 70.090 248.280 71.690 248.390 ;
        RECT 70.090 248.240 78.920 248.280 ;
        RECT 70.090 248.070 79.050 248.240 ;
        RECT 70.090 248.020 78.920 248.070 ;
        RECT 70.090 247.780 71.690 248.020 ;
        RECT 65.170 244.960 66.600 244.970 ;
        RECT 58.180 244.920 66.600 244.960 ;
        RECT 57.820 244.750 66.600 244.920 ;
        RECT 58.180 244.700 66.600 244.750 ;
        RECT 55.140 241.680 59.600 241.970 ;
        RECT 55.140 241.420 65.890 241.680 ;
        RECT 66.260 241.540 66.600 244.700 ;
        RECT 55.140 241.380 59.600 241.420 ;
        RECT 52.940 238.440 53.310 241.360 ;
        RECT 55.140 240.120 56.230 241.380 ;
        RECT 56.770 241.310 58.370 241.380 ;
        RECT 66.210 241.330 66.600 241.540 ;
        RECT 68.390 241.840 69.230 242.470 ;
        RECT 70.120 241.950 70.580 247.780 ;
        RECT 79.530 245.000 79.870 251.320 ;
        RECT 83.250 261.420 91.980 261.470 ;
        RECT 83.250 261.250 92.180 261.420 ;
        RECT 83.250 261.220 91.980 261.250 ;
        RECT 83.250 260.980 84.940 261.220 ;
        RECT 83.250 254.980 83.710 260.980 ;
        RECT 92.660 258.170 93.000 264.390 ;
        RECT 96.680 261.720 98.090 261.770 ;
        RECT 96.680 261.640 102.070 261.720 ;
        RECT 96.680 261.470 102.130 261.640 ;
        RECT 96.680 261.430 102.070 261.470 ;
        RECT 96.680 261.290 98.090 261.430 ;
        RECT 84.390 258.130 93.000 258.170 ;
        RECT 84.220 257.960 93.000 258.130 ;
        RECT 84.390 257.910 93.000 257.960 ;
        RECT 91.560 257.900 93.000 257.910 ;
        RECT 83.250 254.870 84.870 254.980 ;
        RECT 83.250 254.840 92.000 254.870 ;
        RECT 83.250 254.670 92.180 254.840 ;
        RECT 83.250 254.610 92.000 254.670 ;
        RECT 83.250 254.370 84.870 254.610 ;
        RECT 83.250 248.410 83.710 254.370 ;
        RECT 92.660 251.610 93.000 257.900 ;
        RECT 91.620 251.600 93.000 251.610 ;
        RECT 84.460 251.550 93.000 251.600 ;
        RECT 84.220 251.380 93.000 251.550 ;
        RECT 84.460 251.340 93.000 251.380 ;
        RECT 83.220 248.300 84.820 248.410 ;
        RECT 83.220 248.260 92.050 248.300 ;
        RECT 83.220 248.090 92.180 248.260 ;
        RECT 83.220 248.040 92.050 248.090 ;
        RECT 83.220 247.800 84.820 248.040 ;
        RECT 78.440 244.990 79.870 245.000 ;
        RECT 71.450 244.950 79.870 244.990 ;
        RECT 71.090 244.780 79.870 244.950 ;
        RECT 71.450 244.730 79.870 244.780 ;
        RECT 70.040 241.840 71.640 241.950 ;
        RECT 68.390 241.710 72.300 241.840 ;
        RECT 68.390 241.450 79.160 241.710 ;
        RECT 79.530 241.570 79.870 244.730 ;
        RECT 38.990 238.410 40.100 238.440 ;
        RECT 52.220 238.410 53.330 238.440 ;
        RECT 66.210 238.410 66.580 241.330 ;
        RECT 68.390 241.250 72.300 241.450 ;
        RECT 79.480 241.360 79.870 241.570 ;
        RECT 81.470 242.010 82.740 242.180 ;
        RECT 83.250 242.010 83.710 247.800 ;
        RECT 92.660 245.020 93.000 251.340 ;
        RECT 96.760 255.190 97.100 261.290 ;
        RECT 98.060 258.370 102.070 258.400 ;
        RECT 102.390 258.370 102.800 264.390 ;
        RECT 210.780 263.570 211.190 269.690 ;
        RECT 226.980 266.780 227.250 272.970 ;
        RECT 230.820 270.060 231.230 276.290 ;
        RECT 247.020 273.340 247.290 279.600 ;
        RECT 250.880 276.600 252.310 276.670 ;
        RECT 250.880 276.540 266.560 276.600 ;
        RECT 250.880 276.370 266.590 276.540 ;
        RECT 250.880 276.330 266.560 276.370 ;
        RECT 250.880 276.290 252.310 276.330 ;
        RECT 246.270 273.310 247.590 273.340 ;
        RECT 232.320 273.250 247.590 273.310 ;
        RECT 231.630 273.080 247.590 273.250 ;
        RECT 232.320 273.040 247.590 273.080 ;
        RECT 246.270 272.960 247.590 273.040 ;
        RECT 230.800 270.020 232.400 270.060 ;
        RECT 230.800 269.750 246.540 270.020 ;
        RECT 230.800 269.680 232.400 269.750 ;
        RECT 226.080 266.710 227.400 266.780 ;
        RECT 212.270 266.680 227.400 266.710 ;
        RECT 211.590 266.510 227.400 266.680 ;
        RECT 212.270 266.440 227.400 266.510 ;
        RECT 226.080 266.400 227.400 266.440 ;
        RECT 226.980 266.390 227.250 266.400 ;
        RECT 98.060 258.350 102.800 258.370 ;
        RECT 97.640 258.180 102.800 258.350 ;
        RECT 98.060 258.110 102.800 258.180 ;
        RECT 101.520 258.020 102.800 258.110 ;
        RECT 96.760 255.140 98.190 255.190 ;
        RECT 96.760 255.060 102.110 255.140 ;
        RECT 96.760 254.890 102.130 255.060 ;
        RECT 96.760 254.850 102.110 254.890 ;
        RECT 96.760 254.710 98.190 254.850 ;
        RECT 96.760 248.550 97.100 254.710 ;
        RECT 98.120 251.780 102.130 251.800 ;
        RECT 102.390 251.780 102.800 258.020 ;
        RECT 210.690 263.540 211.190 263.570 ;
        RECT 210.690 263.490 212.260 263.540 ;
        RECT 230.820 263.530 231.230 269.680 ;
        RECT 247.020 266.770 247.290 272.960 ;
        RECT 250.880 270.060 251.290 276.290 ;
        RECT 267.080 273.340 267.350 279.600 ;
        RECT 270.930 276.600 272.360 276.670 ;
        RECT 270.930 276.540 286.610 276.600 ;
        RECT 270.930 276.370 286.640 276.540 ;
        RECT 270.930 276.330 286.610 276.370 ;
        RECT 270.930 276.290 272.360 276.330 ;
        RECT 266.330 273.310 267.650 273.340 ;
        RECT 252.380 273.250 267.650 273.310 ;
        RECT 251.690 273.080 267.650 273.250 ;
        RECT 252.380 273.040 267.650 273.080 ;
        RECT 266.330 272.960 267.650 273.040 ;
        RECT 250.860 270.020 252.460 270.060 ;
        RECT 250.860 269.750 266.600 270.020 ;
        RECT 250.860 269.680 252.460 269.750 ;
        RECT 246.120 266.700 247.440 266.770 ;
        RECT 232.310 266.670 247.440 266.700 ;
        RECT 231.630 266.500 247.440 266.670 ;
        RECT 232.310 266.430 247.440 266.500 ;
        RECT 246.120 266.390 247.440 266.430 ;
        RECT 247.020 266.380 247.290 266.390 ;
        RECT 250.880 263.530 251.290 269.680 ;
        RECT 267.080 266.770 267.350 272.960 ;
        RECT 270.930 270.060 271.340 276.290 ;
        RECT 287.130 273.340 287.400 279.600 ;
        RECT 355.040 275.900 356.120 290.200 ;
        RECT 356.460 276.840 356.740 290.440 ;
        RECT 359.820 290.120 359.990 290.280 ;
        RECT 356.460 275.960 356.860 276.840 ;
        RECT 359.770 276.120 360.050 290.120 ;
        RECT 363.050 290.100 363.330 290.730 ;
        RECT 369.600 290.680 370.530 290.730 ;
        RECT 375.760 290.840 376.140 295.680 ;
        RECT 382.360 294.660 382.640 308.720 ;
        RECT 388.920 308.570 389.300 309.460 ;
        RECT 382.430 294.160 382.600 294.660 ;
        RECT 388.930 294.470 389.210 308.570 ;
        RECT 393.610 294.750 394.690 309.050 ;
        RECT 395.030 295.750 395.310 309.580 ;
        RECT 398.390 308.970 398.560 309.130 ;
        RECT 389.010 294.160 389.180 294.470 ;
        RECT 388.960 290.880 389.850 290.930 ;
        RECT 388.920 290.840 389.850 290.880 ;
        RECT 286.380 273.310 287.700 273.340 ;
        RECT 272.430 273.250 287.700 273.310 ;
        RECT 271.740 273.080 287.700 273.250 ;
        RECT 272.430 273.040 287.700 273.080 ;
        RECT 286.380 272.960 287.700 273.040 ;
        RECT 270.910 270.020 272.510 270.060 ;
        RECT 270.910 269.750 286.650 270.020 ;
        RECT 270.910 269.680 272.510 269.750 ;
        RECT 266.180 266.700 267.500 266.770 ;
        RECT 252.370 266.670 267.500 266.700 ;
        RECT 251.690 266.500 267.500 266.670 ;
        RECT 252.370 266.430 267.500 266.500 ;
        RECT 266.180 266.390 267.500 266.430 ;
        RECT 267.080 266.380 267.350 266.390 ;
        RECT 270.930 263.530 271.340 269.680 ;
        RECT 287.130 266.770 287.400 272.960 ;
        RECT 356.480 272.080 356.860 275.960 ;
        RECT 359.720 275.900 360.050 276.120 ;
        RECT 363.040 289.940 363.330 290.100 ;
        RECT 359.720 274.910 360.020 275.900 ;
        RECT 363.040 275.880 363.320 289.940 ;
        RECT 366.400 289.890 366.570 290.280 ;
        RECT 366.340 276.110 366.620 289.890 ;
        RECT 369.600 289.790 369.980 290.680 ;
        RECT 375.760 290.630 389.850 290.840 ;
        RECT 375.760 290.340 376.140 290.630 ;
        RECT 363.110 275.380 363.280 275.880 ;
        RECT 366.340 275.670 366.660 276.110 ;
        RECT 369.610 275.690 369.890 289.790 ;
        RECT 374.360 275.800 375.440 290.100 ;
        RECT 375.780 276.740 376.060 290.340 ;
        RECT 382.370 290.000 382.650 290.630 ;
        RECT 382.360 289.840 382.650 290.000 ;
        RECT 388.920 290.580 389.850 290.630 ;
        RECT 395.010 290.910 395.390 295.750 ;
        RECT 398.340 294.970 398.620 308.970 ;
        RECT 401.620 308.950 401.900 309.580 ;
        RECT 408.170 309.530 409.100 309.580 ;
        RECT 398.290 294.750 398.620 294.970 ;
        RECT 401.610 308.790 401.900 308.950 ;
        RECT 398.290 293.760 398.590 294.750 ;
        RECT 401.610 294.730 401.890 308.790 ;
        RECT 404.970 308.740 405.140 309.130 ;
        RECT 404.910 294.960 405.190 308.740 ;
        RECT 408.170 308.640 408.550 309.530 ;
        RECT 401.680 294.230 401.850 294.730 ;
        RECT 404.910 294.520 405.230 294.960 ;
        RECT 408.180 294.540 408.460 308.640 ;
        RECT 796.480 308.015 811.840 308.185 ;
        RECT 797.110 306.755 797.700 307.735 ;
        RECT 799.500 307.400 799.830 307.735 ;
        RECT 801.930 307.255 802.880 307.735 ;
        RECT 804.270 307.485 805.220 307.785 ;
        RECT 806.965 306.705 807.915 307.735 ;
        RECT 808.750 306.915 809.645 307.735 ;
        RECT 810.255 306.225 811.200 307.765 ;
        RECT 812.180 307.320 813.390 308.140 ;
        RECT 814.240 308.015 829.600 308.185 ;
        RECT 814.870 306.755 815.460 307.735 ;
        RECT 817.260 307.400 817.590 307.735 ;
        RECT 819.690 307.255 820.640 307.735 ;
        RECT 822.030 307.485 822.980 307.785 ;
        RECT 824.725 306.705 825.675 307.735 ;
        RECT 826.510 306.915 827.405 307.735 ;
        RECT 828.015 306.225 828.960 307.765 ;
        RECT 830.070 307.320 831.280 308.170 ;
        RECT 831.780 307.985 833.220 308.155 ;
        RECT 835.420 308.045 840.700 308.215 ;
        RECT 831.870 306.175 832.460 307.755 ;
        RECT 835.980 306.845 837.950 307.815 ;
        RECT 838.480 307.365 840.140 307.815 ;
        RECT 841.170 307.300 842.380 308.150 ;
        RECT 842.690 308.045 844.130 308.215 ;
        RECT 842.780 306.235 843.370 307.815 ;
        RECT 680.060 298.955 695.420 299.125 ;
        RECT 680.690 297.695 681.280 298.675 ;
        RECT 683.080 298.340 683.410 298.675 ;
        RECT 685.510 298.195 686.460 298.675 ;
        RECT 687.850 298.425 688.800 298.725 ;
        RECT 690.545 297.645 691.495 298.675 ;
        RECT 692.330 297.855 693.225 298.675 ;
        RECT 693.835 297.165 694.780 298.705 ;
        RECT 695.850 297.880 696.860 299.030 ;
        RECT 697.550 298.915 712.910 299.085 ;
        RECT 698.180 297.655 698.770 298.635 ;
        RECT 700.570 298.300 700.900 298.635 ;
        RECT 703.000 298.155 703.950 298.635 ;
        RECT 705.340 298.385 706.290 298.685 ;
        RECT 708.035 297.605 708.985 298.635 ;
        RECT 709.820 297.815 710.715 298.635 ;
        RECT 711.325 297.125 712.270 298.665 ;
        RECT 713.500 298.240 714.440 299.110 ;
        RECT 715.160 298.975 730.520 299.145 ;
        RECT 715.790 297.715 716.380 298.695 ;
        RECT 718.180 298.360 718.510 298.695 ;
        RECT 720.610 298.215 721.560 298.695 ;
        RECT 722.950 298.445 723.900 298.745 ;
        RECT 725.645 297.665 726.595 298.695 ;
        RECT 727.430 297.875 728.325 298.695 ;
        RECT 728.935 297.185 729.880 298.725 ;
        RECT 731.130 298.080 732.050 299.060 ;
        RECT 732.860 298.925 748.220 299.095 ;
        RECT 733.490 297.665 734.080 298.645 ;
        RECT 735.880 298.310 736.210 298.645 ;
        RECT 738.310 298.165 739.260 298.645 ;
        RECT 740.650 298.395 741.600 298.695 ;
        RECT 743.345 297.615 744.295 298.645 ;
        RECT 745.130 297.825 746.025 298.645 ;
        RECT 746.635 297.135 747.580 298.675 ;
        RECT 748.900 298.060 749.740 299.080 ;
        RECT 750.600 298.915 765.960 299.085 ;
        RECT 751.230 297.655 751.820 298.635 ;
        RECT 753.620 298.300 753.950 298.635 ;
        RECT 756.050 298.155 757.000 298.635 ;
        RECT 758.390 298.385 759.340 298.685 ;
        RECT 761.085 297.605 762.035 298.635 ;
        RECT 762.870 297.815 763.765 298.635 ;
        RECT 764.375 297.125 765.320 298.665 ;
        RECT 855.800 298.275 859.160 298.445 ;
        RECT 855.890 296.545 856.820 297.995 ;
        RECT 857.350 296.545 858.600 298.045 ;
        RECT 859.720 297.680 860.310 298.420 ;
        RECT 839.390 296.295 842.750 296.465 ;
        RECT 404.930 293.780 405.230 294.520 ;
        RECT 408.260 294.230 408.430 294.540 ;
        RECT 404.930 293.760 405.720 293.780 ;
        RECT 398.290 293.450 405.720 293.760 ;
        RECT 398.290 293.420 398.590 293.450 ;
        RECT 404.930 293.410 405.230 293.450 ;
        RECT 595.170 293.345 596.610 293.515 ;
        RECT 595.930 291.535 596.520 293.115 ;
        RECT 600.980 292.650 601.720 295.510 ;
        RECT 602.430 294.700 602.600 295.120 ;
        RECT 604.010 294.700 604.180 295.120 ;
        RECT 605.590 294.700 605.760 295.120 ;
        RECT 606.950 294.710 607.120 295.130 ;
        RECT 608.530 294.710 608.700 295.130 ;
        RECT 610.110 294.710 610.280 295.130 ;
        RECT 611.470 294.710 611.640 295.130 ;
        RECT 613.050 294.710 613.220 295.130 ;
        RECT 614.630 294.710 614.800 295.130 ;
        RECT 615.900 294.690 616.070 295.110 ;
        RECT 617.480 294.690 617.650 295.110 ;
        RECT 619.060 294.690 619.230 295.110 ;
        RECT 620.280 294.700 620.450 295.120 ;
        RECT 621.860 294.700 622.030 295.120 ;
        RECT 623.440 294.700 623.610 295.120 ;
        RECT 624.600 294.690 624.770 295.110 ;
        RECT 626.180 294.690 626.350 295.110 ;
        RECT 627.760 294.690 627.930 295.110 ;
        RECT 602.430 293.230 602.600 293.650 ;
        RECT 604.010 293.230 604.180 293.650 ;
        RECT 605.590 293.230 605.760 293.650 ;
        RECT 606.950 293.240 607.120 293.660 ;
        RECT 608.530 293.240 608.700 293.660 ;
        RECT 610.110 293.240 610.280 293.660 ;
        RECT 611.470 293.240 611.640 293.660 ;
        RECT 613.050 293.240 613.220 293.660 ;
        RECT 614.630 293.240 614.800 293.660 ;
        RECT 615.900 293.220 616.070 293.640 ;
        RECT 617.480 293.220 617.650 293.640 ;
        RECT 619.060 293.220 619.230 293.640 ;
        RECT 620.280 293.230 620.450 293.650 ;
        RECT 621.860 293.230 622.030 293.650 ;
        RECT 623.440 293.230 623.610 293.650 ;
        RECT 624.600 293.220 624.770 293.640 ;
        RECT 626.180 293.220 626.350 293.640 ;
        RECT 627.760 293.220 627.930 293.640 ;
        RECT 628.680 292.480 629.550 295.800 ;
        RECT 839.480 294.565 840.410 296.015 ;
        RECT 840.940 294.565 842.190 296.065 ;
        RECT 843.310 295.390 844.180 296.430 ;
        RECT 845.090 294.645 848.450 294.815 ;
        RECT 635.060 293.795 636.500 293.965 ;
        RECT 639.250 293.885 640.690 294.055 ;
        RECT 643.350 293.865 644.790 294.035 ;
        RECT 635.150 291.985 635.740 293.565 ;
        RECT 639.340 292.075 639.930 293.655 ;
        RECT 643.440 292.055 644.030 293.635 ;
        RECT 645.310 292.340 645.950 293.650 ;
        RECT 818.940 293.285 822.300 293.455 ;
        RECT 819.030 291.555 819.960 293.005 ;
        RECT 820.490 291.555 821.740 293.055 ;
        RECT 845.920 292.915 847.890 294.415 ;
        RECT 861.180 294.375 864.540 294.545 ;
        RECT 822.770 292.210 823.750 292.830 ;
        RECT 855.840 292.745 859.200 292.915 ;
        RECT 862.010 292.645 863.980 294.145 ;
        RECT 824.390 291.115 827.750 291.285 ;
        RECT 408.210 290.950 409.100 291.000 ;
        RECT 408.170 290.910 409.100 290.950 ;
        RECT 395.010 290.700 409.100 290.910 ;
        RECT 375.780 275.860 376.180 276.740 ;
        RECT 366.360 274.930 366.660 275.670 ;
        RECT 369.690 275.380 369.860 275.690 ;
        RECT 366.360 274.910 367.150 274.930 ;
        RECT 359.720 274.600 367.150 274.910 ;
        RECT 359.720 274.570 360.020 274.600 ;
        RECT 366.360 274.560 366.660 274.600 ;
        RECT 369.660 272.120 370.550 272.170 ;
        RECT 369.620 272.080 370.550 272.120 ;
        RECT 356.460 271.870 370.550 272.080 ;
        RECT 375.800 271.980 376.180 275.860 ;
        RECT 382.360 275.780 382.640 289.840 ;
        RECT 388.920 289.690 389.300 290.580 ;
        RECT 395.010 290.410 395.390 290.700 ;
        RECT 382.430 275.280 382.600 275.780 ;
        RECT 388.930 275.590 389.210 289.690 ;
        RECT 393.610 275.870 394.690 290.170 ;
        RECT 395.030 276.810 395.310 290.410 ;
        RECT 398.390 290.090 398.560 290.250 ;
        RECT 395.030 275.930 395.430 276.810 ;
        RECT 398.340 276.090 398.620 290.090 ;
        RECT 401.620 290.070 401.900 290.700 ;
        RECT 408.170 290.650 409.100 290.700 ;
        RECT 389.010 275.280 389.180 275.590 ;
        RECT 388.980 272.020 389.870 272.070 ;
        RECT 395.050 272.050 395.430 275.930 ;
        RECT 398.290 275.870 398.620 276.090 ;
        RECT 401.610 289.910 401.900 290.070 ;
        RECT 398.290 274.880 398.590 275.870 ;
        RECT 401.610 275.850 401.890 289.910 ;
        RECT 404.970 289.860 405.140 290.250 ;
        RECT 404.910 276.080 405.190 289.860 ;
        RECT 408.170 289.760 408.550 290.650 ;
        RECT 401.680 275.350 401.850 275.850 ;
        RECT 404.910 275.640 405.230 276.080 ;
        RECT 408.180 275.660 408.460 289.760 ;
        RECT 824.480 289.385 825.410 290.835 ;
        RECT 825.940 289.385 827.190 290.885 ;
        RECT 828.220 290.410 828.930 291.270 ;
        RECT 829.930 291.135 835.210 291.305 ;
        RECT 839.400 291.175 842.760 291.345 ;
        RECT 855.930 291.015 856.860 292.465 ;
        RECT 857.390 291.015 858.640 292.515 ;
        RECT 830.490 289.935 832.460 290.905 ;
        RECT 832.990 290.455 834.650 290.905 ;
        RECT 839.490 289.445 840.420 290.895 ;
        RECT 840.950 289.445 842.200 290.945 ;
        RECT 818.910 288.125 822.270 288.295 ;
        RECT 819.000 286.395 819.930 287.845 ;
        RECT 820.460 286.395 821.710 287.895 ;
        RECT 855.910 287.345 859.270 287.515 ;
        RECT 856.000 285.615 856.930 287.065 ;
        RECT 857.460 285.615 858.710 287.115 ;
        RECT 860.060 285.200 860.940 286.160 ;
        RECT 861.260 285.325 864.620 285.495 ;
        RECT 799.530 283.435 800.970 283.605 ;
        RECT 862.090 283.595 864.060 285.095 ;
        RECT 679.390 282.215 684.670 282.385 ;
        RECT 679.950 281.015 681.920 281.985 ;
        RECT 682.450 281.535 684.110 281.985 ;
        RECT 685.190 281.630 685.940 282.340 ;
        RECT 696.670 282.225 701.950 282.395 ;
        RECT 697.230 281.025 699.200 281.995 ;
        RECT 699.730 281.545 701.390 281.995 ;
        RECT 702.800 281.400 703.490 282.380 ;
        RECT 714.440 282.225 719.720 282.395 ;
        RECT 715.000 281.025 716.970 281.995 ;
        RECT 717.500 281.545 719.160 281.995 ;
        RECT 720.220 281.450 721.180 282.330 ;
        RECT 731.680 282.225 736.960 282.395 ;
        RECT 732.240 281.025 734.210 281.995 ;
        RECT 734.740 281.545 736.400 281.995 ;
        RECT 737.630 281.300 738.670 282.440 ;
        RECT 749.160 282.235 754.440 282.405 ;
        RECT 749.720 281.035 751.690 282.005 ;
        RECT 752.220 281.555 753.880 282.005 ;
        RECT 754.830 281.640 755.580 282.390 ;
        RECT 799.620 281.625 800.210 283.205 ;
        RECT 819.350 283.095 824.630 283.265 ;
        RECT 841.640 283.175 841.990 283.290 ;
        RECT 827.960 283.005 831.320 283.175 ;
        RECT 819.910 281.895 821.880 282.865 ;
        RECT 822.410 282.415 824.070 282.865 ;
        RECT 828.050 281.275 828.980 282.725 ;
        RECT 829.510 281.275 830.760 282.775 ;
        RECT 831.640 282.250 832.740 283.090 ;
        RECT 833.250 283.005 838.530 283.175 ;
        RECT 833.810 281.805 835.780 282.775 ;
        RECT 836.310 282.325 837.970 282.775 ;
        RECT 838.950 282.390 839.860 283.110 ;
        RECT 840.460 283.005 844.300 283.175 ;
        RECT 846.300 283.005 851.580 283.175 ;
        RECT 841.640 282.725 841.990 283.005 ;
        RECT 841.020 282.400 841.990 282.725 ;
        RECT 841.020 281.690 841.970 282.400 ;
        RECT 842.660 281.195 843.610 282.775 ;
        RECT 846.860 281.805 848.830 282.775 ;
        RECT 849.360 282.325 851.020 282.775 ;
        RECT 851.880 282.530 852.500 283.150 ;
        RECT 855.930 281.885 859.290 282.055 ;
        RECT 699.550 280.390 699.880 280.400 ;
        RECT 717.340 280.390 717.670 280.440 ;
        RECT 734.600 280.390 734.930 280.470 ;
        RECT 752.070 280.400 752.400 280.460 ;
        RECT 681.435 280.005 682.625 280.380 ;
        RECT 698.715 280.015 699.905 280.390 ;
        RECT 716.485 280.015 717.675 280.390 ;
        RECT 733.725 280.190 734.930 280.390 ;
        RECT 733.725 280.015 734.915 280.190 ;
        RECT 751.205 280.180 752.400 280.400 ;
        RECT 751.205 280.025 752.395 280.180 ;
        RECT 856.020 280.155 856.950 281.605 ;
        RECT 857.480 280.155 858.730 281.655 ;
        RECT 404.930 274.900 405.230 275.640 ;
        RECT 408.260 275.350 408.430 275.660 ;
        RECT 404.930 274.880 405.720 274.900 ;
        RECT 398.290 274.570 405.720 274.880 ;
        RECT 595.090 274.875 596.530 275.045 ;
        RECT 409.470 274.730 409.640 274.770 ;
        RECT 409.470 274.590 410.640 274.730 ;
        RECT 398.290 274.540 398.590 274.570 ;
        RECT 404.930 274.530 405.230 274.570 ;
        RECT 408.230 272.090 409.120 272.140 ;
        RECT 408.190 272.050 409.120 272.090 ;
        RECT 388.940 271.980 389.870 272.020 ;
        RECT 356.480 271.500 356.860 271.870 ;
        RECT 286.230 266.700 287.550 266.770 ;
        RECT 272.420 266.670 287.550 266.700 ;
        RECT 271.740 266.500 287.550 266.670 ;
        RECT 272.420 266.430 287.550 266.500 ;
        RECT 286.230 266.390 287.550 266.430 ;
        RECT 230.800 263.490 232.300 263.530 ;
        RECT 250.860 263.490 252.360 263.530 ;
        RECT 270.910 263.490 272.410 263.530 ;
        RECT 210.690 263.430 285.990 263.490 ;
        RECT 210.690 263.380 286.620 263.430 ;
        RECT 210.690 263.230 286.640 263.380 ;
        RECT 210.690 263.220 226.490 263.230 ;
        RECT 210.690 263.170 226.470 263.220 ;
        RECT 230.800 263.210 246.530 263.230 ;
        RECT 250.860 263.210 266.590 263.230 ;
        RECT 270.910 263.210 286.640 263.230 ;
        RECT 210.690 263.160 212.170 263.170 ;
        RECT 230.800 263.160 246.510 263.210 ;
        RECT 250.860 263.160 266.570 263.210 ;
        RECT 270.910 263.160 286.620 263.210 ;
        RECT 210.690 263.150 211.190 263.160 ;
        RECT 230.800 263.150 232.210 263.160 ;
        RECT 250.860 263.150 252.270 263.160 ;
        RECT 270.910 263.150 272.320 263.160 ;
        RECT 210.690 255.690 211.100 263.150 ;
        RECT 230.820 263.140 231.230 263.150 ;
        RECT 250.880 263.140 251.290 263.150 ;
        RECT 270.930 263.140 271.340 263.150 ;
        RECT 213.350 259.540 226.580 261.550 ;
        RECT 233.320 259.540 246.550 261.550 ;
        RECT 253.430 259.540 266.660 261.550 ;
        RECT 273.540 259.540 286.770 261.550 ;
        RECT 287.110 261.520 287.540 266.390 ;
        RECT 288.050 261.520 289.000 262.250 ;
        RECT 287.110 260.270 289.000 261.520 ;
        RECT 287.110 259.000 287.540 260.270 ;
        RECT 288.050 259.540 289.000 260.270 ;
        RECT 226.010 258.910 227.330 259.000 ;
        RECT 245.980 258.910 247.300 259.000 ;
        RECT 266.090 258.910 267.410 259.000 ;
        RECT 286.200 258.910 287.540 259.000 ;
        RECT 212.000 258.850 287.540 258.910 ;
        RECT 211.550 258.680 287.540 258.850 ;
        RECT 212.000 258.660 287.540 258.680 ;
        RECT 212.000 258.650 287.520 258.660 ;
        RECT 212.000 258.640 227.330 258.650 ;
        RECT 231.970 258.640 247.300 258.650 ;
        RECT 252.080 258.640 267.410 258.650 ;
        RECT 272.190 258.640 287.520 258.650 ;
        RECT 226.010 258.620 227.330 258.640 ;
        RECT 245.980 258.620 247.300 258.640 ;
        RECT 266.090 258.620 267.410 258.640 ;
        RECT 286.200 258.620 287.520 258.640 ;
        RECT 210.690 255.620 212.170 255.690 ;
        RECT 210.690 255.560 226.420 255.620 ;
        RECT 210.690 255.390 226.450 255.560 ;
        RECT 210.690 255.350 226.420 255.390 ;
        RECT 210.690 255.310 212.170 255.350 ;
        RECT 210.690 254.810 211.150 255.310 ;
        RECT 98.120 251.770 102.890 251.780 ;
        RECT 97.640 251.600 102.890 251.770 ;
        RECT 98.120 251.510 102.890 251.600 ;
        RECT 101.670 251.430 102.890 251.510 ;
        RECT 96.740 248.480 102.050 248.550 ;
        RECT 96.740 248.310 102.130 248.480 ;
        RECT 96.740 248.260 102.050 248.310 ;
        RECT 96.740 248.070 98.150 248.260 ;
        RECT 91.570 245.010 93.000 245.020 ;
        RECT 84.580 244.970 93.000 245.010 ;
        RECT 84.220 244.800 93.000 244.970 ;
        RECT 84.580 244.750 93.000 244.800 ;
        RECT 81.470 241.730 85.170 242.010 ;
        RECT 81.470 241.470 92.290 241.730 ;
        RECT 92.660 241.590 93.000 244.750 ;
        RECT 68.390 240.330 69.230 241.250 ;
        RECT 79.480 238.440 79.850 241.360 ;
        RECT 81.470 241.220 85.170 241.470 ;
        RECT 92.610 241.380 93.000 241.590 ;
        RECT 94.220 242.390 95.270 242.640 ;
        RECT 96.760 242.390 97.100 248.070 ;
        RECT 102.390 245.260 102.800 251.430 ;
        RECT 210.740 249.080 211.150 254.810 ;
        RECT 226.940 252.360 227.210 258.620 ;
        RECT 230.710 255.620 232.140 255.690 ;
        RECT 230.710 255.560 246.390 255.620 ;
        RECT 230.710 255.390 246.420 255.560 ;
        RECT 230.710 255.350 246.390 255.390 ;
        RECT 230.710 255.310 232.140 255.350 ;
        RECT 226.190 252.330 227.510 252.360 ;
        RECT 212.240 252.270 227.510 252.330 ;
        RECT 211.550 252.100 227.510 252.270 ;
        RECT 212.240 252.060 227.510 252.100 ;
        RECT 226.190 251.980 227.510 252.060 ;
        RECT 210.720 249.040 212.320 249.080 ;
        RECT 210.720 248.770 226.460 249.040 ;
        RECT 210.720 248.700 212.320 248.770 ;
        RECT 101.580 245.200 102.800 245.260 ;
        RECT 98.040 245.190 102.800 245.200 ;
        RECT 97.640 245.020 102.800 245.190 ;
        RECT 98.040 244.910 102.800 245.020 ;
        RECT 94.220 242.000 97.100 242.390 ;
        RECT 102.390 243.690 102.800 244.910 ;
        RECT 103.270 243.690 103.830 243.790 ;
        RECT 102.390 243.490 103.830 243.690 ;
        RECT 94.220 241.950 98.170 242.000 ;
        RECT 94.220 241.930 101.970 241.950 ;
        RECT 102.390 241.930 102.800 243.490 ;
        RECT 103.270 243.330 103.830 243.490 ;
        RECT 210.740 242.550 211.150 248.700 ;
        RECT 226.940 245.790 227.210 251.980 ;
        RECT 230.710 249.080 231.120 255.310 ;
        RECT 246.910 252.360 247.180 258.620 ;
        RECT 250.820 255.620 252.250 255.690 ;
        RECT 250.820 255.560 266.500 255.620 ;
        RECT 250.820 255.390 266.530 255.560 ;
        RECT 250.820 255.350 266.500 255.390 ;
        RECT 250.820 255.310 252.250 255.350 ;
        RECT 246.160 252.330 247.480 252.360 ;
        RECT 232.210 252.270 247.480 252.330 ;
        RECT 231.520 252.100 247.480 252.270 ;
        RECT 232.210 252.060 247.480 252.100 ;
        RECT 246.160 251.980 247.480 252.060 ;
        RECT 230.690 249.040 232.290 249.080 ;
        RECT 230.690 248.770 246.430 249.040 ;
        RECT 230.690 248.700 232.290 248.770 ;
        RECT 226.040 245.720 227.360 245.790 ;
        RECT 212.230 245.690 227.360 245.720 ;
        RECT 211.550 245.520 227.360 245.690 ;
        RECT 212.230 245.450 227.360 245.520 ;
        RECT 226.040 245.410 227.360 245.450 ;
        RECT 226.940 245.400 227.210 245.410 ;
        RECT 230.710 242.550 231.120 248.700 ;
        RECT 246.910 245.790 247.180 251.980 ;
        RECT 250.820 249.080 251.230 255.310 ;
        RECT 267.020 252.360 267.290 258.620 ;
        RECT 286.930 257.910 287.400 258.620 ;
        RECT 270.930 255.620 272.360 255.690 ;
        RECT 270.930 255.560 286.610 255.620 ;
        RECT 270.930 255.390 286.640 255.560 ;
        RECT 270.930 255.350 286.610 255.390 ;
        RECT 270.930 255.310 272.360 255.350 ;
        RECT 266.270 252.330 267.590 252.360 ;
        RECT 252.320 252.270 267.590 252.330 ;
        RECT 251.630 252.100 267.590 252.270 ;
        RECT 252.320 252.060 267.590 252.100 ;
        RECT 266.270 251.980 267.590 252.060 ;
        RECT 250.800 249.040 252.400 249.080 ;
        RECT 250.800 248.770 266.540 249.040 ;
        RECT 250.800 248.700 252.400 248.770 ;
        RECT 246.010 245.720 247.330 245.790 ;
        RECT 232.200 245.690 247.330 245.720 ;
        RECT 231.520 245.520 247.330 245.690 ;
        RECT 232.200 245.450 247.330 245.520 ;
        RECT 246.010 245.410 247.330 245.450 ;
        RECT 246.910 245.400 247.180 245.410 ;
        RECT 250.820 242.550 251.230 248.700 ;
        RECT 267.020 245.790 267.290 251.980 ;
        RECT 270.930 249.080 271.340 255.310 ;
        RECT 287.130 252.360 287.400 257.910 ;
        RECT 355.060 257.040 356.140 271.340 ;
        RECT 356.480 257.100 356.760 271.500 ;
        RECT 359.840 271.260 360.010 271.420 ;
        RECT 359.790 257.260 360.070 271.260 ;
        RECT 363.070 271.240 363.350 271.870 ;
        RECT 369.620 271.820 370.550 271.870 ;
        RECT 356.550 256.520 356.720 257.100 ;
        RECT 359.740 257.040 360.070 257.260 ;
        RECT 363.060 271.080 363.350 271.240 ;
        RECT 359.740 256.050 360.040 257.040 ;
        RECT 363.060 257.020 363.340 271.080 ;
        RECT 366.420 271.030 366.590 271.420 ;
        RECT 366.360 257.250 366.640 271.030 ;
        RECT 369.620 270.930 370.000 271.820 ;
        RECT 375.780 271.770 389.870 271.980 ;
        RECT 395.030 271.840 409.120 272.050 ;
        RECT 375.800 271.400 376.180 271.770 ;
        RECT 363.130 256.520 363.300 257.020 ;
        RECT 366.360 256.810 366.680 257.250 ;
        RECT 369.630 256.830 369.910 270.930 ;
        RECT 374.380 256.940 375.460 271.240 ;
        RECT 375.800 257.000 376.080 271.400 ;
        RECT 382.390 271.140 382.670 271.770 ;
        RECT 382.380 270.980 382.670 271.140 ;
        RECT 388.940 271.720 389.870 271.770 ;
        RECT 366.380 256.070 366.680 256.810 ;
        RECT 369.710 256.520 369.880 256.830 ;
        RECT 375.870 256.420 376.040 257.000 ;
        RECT 382.380 256.920 382.660 270.980 ;
        RECT 388.940 270.830 389.320 271.720 ;
        RECT 395.050 271.470 395.430 271.840 ;
        RECT 382.450 256.420 382.620 256.920 ;
        RECT 388.950 256.730 389.230 270.830 ;
        RECT 393.630 257.010 394.710 271.310 ;
        RECT 395.050 257.070 395.330 271.470 ;
        RECT 398.410 271.230 398.580 271.390 ;
        RECT 398.360 257.230 398.640 271.230 ;
        RECT 401.640 271.210 401.920 271.840 ;
        RECT 408.190 271.790 409.120 271.840 ;
        RECT 389.030 256.420 389.200 256.730 ;
        RECT 395.120 256.490 395.290 257.070 ;
        RECT 398.310 257.010 398.640 257.230 ;
        RECT 401.630 271.050 401.920 271.210 ;
        RECT 366.380 256.050 367.170 256.070 ;
        RECT 359.740 255.740 367.170 256.050 ;
        RECT 398.310 256.020 398.610 257.010 ;
        RECT 401.630 256.990 401.910 271.050 ;
        RECT 404.990 271.000 405.160 271.390 ;
        RECT 404.930 257.220 405.210 271.000 ;
        RECT 408.190 270.900 408.570 271.790 ;
        RECT 401.700 256.490 401.870 256.990 ;
        RECT 404.930 256.780 405.250 257.220 ;
        RECT 408.200 256.800 408.480 270.900 ;
        RECT 409.480 270.540 410.640 274.590 ;
        RECT 595.850 273.065 596.440 274.645 ;
        RECT 600.900 274.180 601.640 277.040 ;
        RECT 602.350 276.230 602.520 276.650 ;
        RECT 603.930 276.230 604.100 276.650 ;
        RECT 605.510 276.230 605.680 276.650 ;
        RECT 606.870 276.240 607.040 276.660 ;
        RECT 608.450 276.240 608.620 276.660 ;
        RECT 610.030 276.240 610.200 276.660 ;
        RECT 611.390 276.240 611.560 276.660 ;
        RECT 612.970 276.240 613.140 276.660 ;
        RECT 614.550 276.240 614.720 276.660 ;
        RECT 615.820 276.220 615.990 276.640 ;
        RECT 617.400 276.220 617.570 276.640 ;
        RECT 618.980 276.220 619.150 276.640 ;
        RECT 620.200 276.230 620.370 276.650 ;
        RECT 621.780 276.230 621.950 276.650 ;
        RECT 623.360 276.230 623.530 276.650 ;
        RECT 624.520 276.220 624.690 276.640 ;
        RECT 626.100 276.220 626.270 276.640 ;
        RECT 627.680 276.220 627.850 276.640 ;
        RECT 602.350 274.760 602.520 275.180 ;
        RECT 603.930 274.760 604.100 275.180 ;
        RECT 605.510 274.760 605.680 275.180 ;
        RECT 606.870 274.770 607.040 275.190 ;
        RECT 608.450 274.770 608.620 275.190 ;
        RECT 610.030 274.770 610.200 275.190 ;
        RECT 611.390 274.770 611.560 275.190 ;
        RECT 612.970 274.770 613.140 275.190 ;
        RECT 614.550 274.770 614.720 275.190 ;
        RECT 615.820 274.750 615.990 275.170 ;
        RECT 617.400 274.750 617.570 275.170 ;
        RECT 618.980 274.750 619.150 275.170 ;
        RECT 620.200 274.760 620.370 275.180 ;
        RECT 621.780 274.760 621.950 275.180 ;
        RECT 623.360 274.760 623.530 275.180 ;
        RECT 624.520 274.750 624.690 275.170 ;
        RECT 626.100 274.750 626.270 275.170 ;
        RECT 627.680 274.750 627.850 275.170 ;
        RECT 628.600 274.010 629.470 277.330 ;
        RECT 679.800 276.555 685.080 276.725 ;
        RECT 634.980 275.325 636.420 275.495 ;
        RECT 639.170 275.415 640.610 275.585 ;
        RECT 643.270 275.395 644.710 275.565 ;
        RECT 680.360 275.355 682.330 276.325 ;
        RECT 682.860 275.875 684.520 276.325 ;
        RECT 685.600 276.010 686.200 276.680 ;
        RECT 687.040 276.515 692.320 276.685 ;
        RECT 697.030 276.575 702.310 276.745 ;
        RECT 687.600 275.315 689.570 276.285 ;
        RECT 690.100 275.835 691.760 276.285 ;
        RECT 697.590 275.375 699.560 276.345 ;
        RECT 700.090 275.895 701.750 276.345 ;
        RECT 702.880 275.940 703.450 276.690 ;
        RECT 704.270 276.535 709.550 276.705 ;
        RECT 714.600 276.675 719.880 276.845 ;
        RECT 704.830 275.335 706.800 276.305 ;
        RECT 707.330 275.855 708.990 276.305 ;
        RECT 715.160 275.475 717.130 276.445 ;
        RECT 717.660 275.995 719.320 276.445 ;
        RECT 720.410 276.070 721.030 276.780 ;
        RECT 721.840 276.635 727.120 276.805 ;
        RECT 731.770 276.705 737.050 276.875 ;
        RECT 722.400 275.435 724.370 276.405 ;
        RECT 724.900 275.955 726.560 276.405 ;
        RECT 732.330 275.505 734.300 276.475 ;
        RECT 734.830 276.025 736.490 276.475 ;
        RECT 737.530 275.930 738.320 276.810 ;
        RECT 739.010 276.665 744.290 276.835 ;
        RECT 749.580 276.765 754.860 276.935 ;
        RECT 739.570 275.465 741.540 276.435 ;
        RECT 742.070 275.985 743.730 276.435 ;
        RECT 750.140 275.565 752.110 276.535 ;
        RECT 752.640 276.085 754.300 276.535 ;
        RECT 755.500 276.300 756.070 276.890 ;
        RECT 756.820 276.725 762.100 276.895 ;
        RECT 757.380 275.525 759.350 276.495 ;
        RECT 759.880 276.045 761.540 276.495 ;
        RECT 780.960 275.395 796.320 275.565 ;
        RECT 635.070 273.515 635.660 275.095 ;
        RECT 639.260 273.605 639.850 275.185 ;
        RECT 643.360 273.585 643.950 275.165 ;
        RECT 645.290 273.900 645.930 275.210 ;
        RECT 757.380 274.515 758.330 274.795 ;
        RECT 758.160 274.335 758.330 274.515 ;
        RECT 760.235 274.335 760.535 274.575 ;
        RECT 758.160 274.245 760.535 274.335 ;
        RECT 758.160 274.165 760.405 274.245 ;
        RECT 781.590 274.135 782.180 275.115 ;
        RECT 783.980 274.780 784.310 275.115 ;
        RECT 786.410 274.635 787.360 275.115 ;
        RECT 788.750 274.865 789.700 275.165 ;
        RECT 791.445 274.085 792.395 275.115 ;
        RECT 793.230 274.295 794.125 275.115 ;
        RECT 794.735 273.605 795.680 275.145 ;
        RECT 796.690 274.920 797.460 275.470 ;
        RECT 799.850 275.385 815.210 275.555 ;
        RECT 800.480 274.125 801.070 275.105 ;
        RECT 802.870 274.770 803.200 275.105 ;
        RECT 805.300 274.625 806.250 275.105 ;
        RECT 807.640 274.855 808.590 275.155 ;
        RECT 810.335 274.075 811.285 275.105 ;
        RECT 812.120 274.285 813.015 275.105 ;
        RECT 813.625 273.595 814.570 275.135 ;
        RECT 815.690 274.980 816.640 275.510 ;
        RECT 818.700 275.355 834.060 275.525 ;
        RECT 819.330 274.095 819.920 275.075 ;
        RECT 821.720 274.740 822.050 275.075 ;
        RECT 824.150 274.595 825.100 275.075 ;
        RECT 826.490 274.825 827.440 275.125 ;
        RECT 829.185 274.045 830.135 275.075 ;
        RECT 830.970 274.255 831.865 275.075 ;
        RECT 832.475 273.565 833.420 275.105 ;
        RECT 837.120 274.930 837.810 275.490 ;
        RECT 838.420 275.395 842.260 275.565 ;
        RECT 855.930 275.345 859.290 275.515 ;
        RECT 838.980 274.080 839.930 275.115 ;
        RECT 840.620 273.585 841.570 275.165 ;
        RECT 856.020 273.615 856.950 275.065 ;
        RECT 857.480 273.615 858.730 275.115 ;
        RECT 844.670 273.135 848.030 273.305 ;
        RECT 850.080 273.145 851.520 273.315 ;
        RECT 844.760 271.405 845.690 272.855 ;
        RECT 846.220 271.405 847.470 272.905 ;
        RECT 850.170 271.335 850.760 272.915 ;
        RECT 860.810 272.690 861.830 273.700 ;
        RECT 861.250 271.955 864.610 272.125 ;
        RECT 679.920 270.875 683.280 271.045 ;
        RECT 685.580 270.885 688.940 271.055 ;
        RECT 680.010 269.145 680.940 270.595 ;
        RECT 681.470 269.145 682.720 270.645 ;
        RECT 685.670 269.155 686.600 270.605 ;
        RECT 687.130 269.155 688.380 270.655 ;
        RECT 689.580 270.120 690.280 271.000 ;
        RECT 690.930 270.905 694.290 271.075 ;
        RECT 697.150 270.895 700.510 271.065 ;
        RECT 691.760 269.175 693.730 270.675 ;
        RECT 697.240 269.165 698.170 270.615 ;
        RECT 698.700 269.165 699.950 270.665 ;
        RECT 701.020 270.120 701.720 271.000 ;
        RECT 702.810 270.905 706.170 271.075 ;
        RECT 708.160 270.925 711.520 271.095 ;
        RECT 714.720 270.995 718.080 271.165 ;
        RECT 702.900 269.175 703.830 270.625 ;
        RECT 704.360 269.175 705.610 270.675 ;
        RECT 708.990 269.195 710.960 270.695 ;
        RECT 714.810 269.265 715.740 270.715 ;
        RECT 716.270 269.265 717.520 270.765 ;
        RECT 718.600 270.360 719.300 271.110 ;
        RECT 720.380 271.005 723.740 271.175 ;
        RECT 725.730 271.025 729.090 271.195 ;
        RECT 731.890 271.025 735.250 271.195 ;
        RECT 720.470 269.275 721.400 270.725 ;
        RECT 721.930 269.275 723.180 270.775 ;
        RECT 726.560 269.295 728.530 270.795 ;
        RECT 731.980 269.295 732.910 270.745 ;
        RECT 733.440 269.295 734.690 270.795 ;
        RECT 735.930 270.260 736.630 271.140 ;
        RECT 737.550 271.035 740.910 271.205 ;
        RECT 742.900 271.055 746.260 271.225 ;
        RECT 749.700 271.085 753.060 271.255 ;
        RECT 737.640 269.305 738.570 270.755 ;
        RECT 739.100 269.305 740.350 270.805 ;
        RECT 743.730 269.325 745.700 270.825 ;
        RECT 749.790 269.355 750.720 270.805 ;
        RECT 751.250 269.355 752.500 270.855 ;
        RECT 753.870 270.300 754.490 271.190 ;
        RECT 755.360 271.095 758.720 271.265 ;
        RECT 760.710 271.115 764.070 271.285 ;
        RECT 755.450 269.365 756.380 270.815 ;
        RECT 756.910 269.365 758.160 270.865 ;
        RECT 761.540 269.385 763.510 270.885 ;
        RECT 862.080 270.225 864.050 271.725 ;
        RECT 838.430 269.835 841.790 270.005 ;
        RECT 756.425 268.640 756.815 268.835 ;
        RECT 756.425 268.060 756.820 268.640 ;
        RECT 838.520 268.105 839.450 269.555 ;
        RECT 839.980 268.105 841.230 269.605 ;
        RECT 856.010 268.675 859.370 268.845 ;
        RECT 756.425 267.920 756.815 268.060 ;
        RECT 780.970 267.835 796.330 268.005 ;
        RECT 781.600 266.575 782.190 267.555 ;
        RECT 783.990 267.220 784.320 267.555 ;
        RECT 786.420 267.075 787.370 267.555 ;
        RECT 788.760 267.305 789.710 267.605 ;
        RECT 791.455 266.525 792.405 267.555 ;
        RECT 793.240 266.735 794.135 267.555 ;
        RECT 794.745 266.045 795.690 267.585 ;
        RECT 796.670 267.460 797.240 267.970 ;
        RECT 799.500 267.895 814.860 268.065 ;
        RECT 800.130 266.635 800.720 267.615 ;
        RECT 802.520 267.280 802.850 267.615 ;
        RECT 804.950 267.135 805.900 267.615 ;
        RECT 807.290 267.365 808.240 267.665 ;
        RECT 809.985 266.585 810.935 267.615 ;
        RECT 811.770 266.795 812.665 267.615 ;
        RECT 813.275 266.105 814.220 267.645 ;
        RECT 815.170 267.430 815.620 268.020 ;
        RECT 856.100 266.945 857.030 268.395 ;
        RECT 857.560 266.945 858.810 268.445 ;
        RECT 679.370 260.685 684.650 260.855 ;
        RECT 594.940 257.145 596.380 257.315 ;
        RECT 404.950 256.040 405.250 256.780 ;
        RECT 408.280 256.490 408.450 256.800 ;
        RECT 404.950 256.020 405.740 256.040 ;
        RECT 359.740 255.710 360.040 255.740 ;
        RECT 366.380 255.700 366.680 255.740 ;
        RECT 398.310 255.710 405.740 256.020 ;
        RECT 398.310 255.680 398.610 255.710 ;
        RECT 404.950 255.670 405.250 255.710 ;
        RECT 595.700 255.335 596.290 256.915 ;
        RECT 600.750 256.450 601.490 259.310 ;
        RECT 602.200 258.500 602.370 258.920 ;
        RECT 603.780 258.500 603.950 258.920 ;
        RECT 605.360 258.500 605.530 258.920 ;
        RECT 606.720 258.510 606.890 258.930 ;
        RECT 608.300 258.510 608.470 258.930 ;
        RECT 609.880 258.510 610.050 258.930 ;
        RECT 611.240 258.510 611.410 258.930 ;
        RECT 612.820 258.510 612.990 258.930 ;
        RECT 614.400 258.510 614.570 258.930 ;
        RECT 615.670 258.490 615.840 258.910 ;
        RECT 617.250 258.490 617.420 258.910 ;
        RECT 618.830 258.490 619.000 258.910 ;
        RECT 620.050 258.500 620.220 258.920 ;
        RECT 621.630 258.500 621.800 258.920 ;
        RECT 623.210 258.500 623.380 258.920 ;
        RECT 624.370 258.490 624.540 258.910 ;
        RECT 625.950 258.490 626.120 258.910 ;
        RECT 627.530 258.490 627.700 258.910 ;
        RECT 602.200 257.030 602.370 257.450 ;
        RECT 603.780 257.030 603.950 257.450 ;
        RECT 605.360 257.030 605.530 257.450 ;
        RECT 606.720 257.040 606.890 257.460 ;
        RECT 608.300 257.040 608.470 257.460 ;
        RECT 609.880 257.040 610.050 257.460 ;
        RECT 611.240 257.040 611.410 257.460 ;
        RECT 612.820 257.040 612.990 257.460 ;
        RECT 614.400 257.040 614.570 257.460 ;
        RECT 615.670 257.020 615.840 257.440 ;
        RECT 617.250 257.020 617.420 257.440 ;
        RECT 618.830 257.020 619.000 257.440 ;
        RECT 620.050 257.030 620.220 257.450 ;
        RECT 621.630 257.030 621.800 257.450 ;
        RECT 623.210 257.030 623.380 257.450 ;
        RECT 624.370 257.020 624.540 257.440 ;
        RECT 625.950 257.020 626.120 257.440 ;
        RECT 627.530 257.020 627.700 257.440 ;
        RECT 628.450 256.280 629.320 259.600 ;
        RECT 679.930 259.485 681.900 260.455 ;
        RECT 682.430 260.005 684.090 260.455 ;
        RECT 685.180 260.060 685.760 260.780 ;
        RECT 696.650 260.695 701.930 260.865 ;
        RECT 697.210 259.495 699.180 260.465 ;
        RECT 699.710 260.015 701.370 260.465 ;
        RECT 702.370 260.200 703.050 260.800 ;
        RECT 714.420 260.695 719.700 260.865 ;
        RECT 714.980 259.495 716.950 260.465 ;
        RECT 717.480 260.015 719.140 260.465 ;
        RECT 720.250 260.210 720.730 260.790 ;
        RECT 731.660 260.695 736.940 260.865 ;
        RECT 732.220 259.495 734.190 260.465 ;
        RECT 734.720 260.015 736.380 260.465 ;
        RECT 737.360 260.390 737.870 260.820 ;
        RECT 749.140 260.705 754.420 260.875 ;
        RECT 749.700 259.505 751.670 260.475 ;
        RECT 752.200 260.025 753.860 260.475 ;
        RECT 755.010 259.840 755.580 260.330 ;
        RECT 855.880 259.365 859.240 259.535 ;
        RECT 634.830 257.595 636.270 257.765 ;
        RECT 639.020 257.685 640.460 257.855 ;
        RECT 643.120 257.665 644.560 257.835 ;
        RECT 855.970 257.635 856.900 259.085 ;
        RECT 857.430 257.635 858.680 259.135 ;
        RECT 634.920 255.785 635.510 257.365 ;
        RECT 639.110 255.875 639.700 257.455 ;
        RECT 860.300 257.450 861.080 258.270 ;
        RECT 643.210 255.855 643.800 257.435 ;
        RECT 645.050 256.060 645.690 257.370 ;
        RECT 861.190 256.875 864.550 257.045 ;
        RECT 679.780 255.025 685.060 255.195 ;
        RECT 680.340 253.825 682.310 254.795 ;
        RECT 682.840 254.345 684.500 254.795 ;
        RECT 685.550 254.350 686.110 255.160 ;
        RECT 687.020 254.985 692.300 255.155 ;
        RECT 697.010 255.045 702.290 255.215 ;
        RECT 687.580 253.785 689.550 254.755 ;
        RECT 690.080 254.305 691.740 254.755 ;
        RECT 697.570 253.845 699.540 254.815 ;
        RECT 700.070 254.365 701.730 254.815 ;
        RECT 702.800 254.410 703.440 255.160 ;
        RECT 704.250 255.005 709.530 255.175 ;
        RECT 714.580 255.145 719.860 255.315 ;
        RECT 704.810 253.805 706.780 254.775 ;
        RECT 707.310 254.325 708.970 254.775 ;
        RECT 715.140 253.945 717.110 254.915 ;
        RECT 717.640 254.465 719.300 254.915 ;
        RECT 720.340 254.470 720.850 255.270 ;
        RECT 721.820 255.105 727.100 255.275 ;
        RECT 731.750 255.175 737.030 255.345 ;
        RECT 722.380 253.905 724.350 254.875 ;
        RECT 724.880 254.425 726.540 254.875 ;
        RECT 732.310 253.975 734.280 254.945 ;
        RECT 734.810 254.495 736.470 254.945 ;
        RECT 737.520 254.580 738.160 255.290 ;
        RECT 738.990 255.135 744.270 255.305 ;
        RECT 749.560 255.235 754.840 255.405 ;
        RECT 739.550 253.935 741.520 254.905 ;
        RECT 742.050 254.455 743.710 254.905 ;
        RECT 750.120 254.035 752.090 255.005 ;
        RECT 752.620 254.555 754.280 255.005 ;
        RECT 755.280 254.720 755.850 255.370 ;
        RECT 756.800 255.195 762.080 255.365 ;
        RECT 862.020 255.145 863.990 256.645 ;
        RECT 757.360 253.995 759.330 254.965 ;
        RECT 759.860 254.515 761.520 254.965 ;
        RECT 855.940 253.595 859.300 253.765 ;
        RECT 699.055 252.835 700.245 253.210 ;
        RECT 286.380 252.330 287.700 252.360 ;
        RECT 272.430 252.270 287.700 252.330 ;
        RECT 271.740 252.100 287.700 252.270 ;
        RECT 272.430 252.060 287.700 252.100 ;
        RECT 286.380 251.980 287.700 252.060 ;
        RECT 270.910 249.040 272.510 249.080 ;
        RECT 270.910 248.770 286.650 249.040 ;
        RECT 270.910 248.700 272.510 248.770 ;
        RECT 266.120 245.720 267.440 245.790 ;
        RECT 252.310 245.690 267.440 245.720 ;
        RECT 251.630 245.520 267.440 245.690 ;
        RECT 252.310 245.450 267.440 245.520 ;
        RECT 266.120 245.410 267.440 245.450 ;
        RECT 267.020 245.400 267.290 245.410 ;
        RECT 270.930 242.550 271.340 248.700 ;
        RECT 287.130 245.920 287.400 251.980 ;
        RECT 856.030 251.865 856.960 253.315 ;
        RECT 857.490 251.865 858.740 253.365 ;
        RECT 679.900 249.345 683.260 249.515 ;
        RECT 679.990 247.615 680.920 249.065 ;
        RECT 681.450 247.615 682.700 249.115 ;
        RECT 684.000 248.700 684.510 249.420 ;
        RECT 685.560 249.355 688.920 249.525 ;
        RECT 690.910 249.375 694.270 249.545 ;
        RECT 697.130 249.365 700.490 249.535 ;
        RECT 685.650 247.625 686.580 249.075 ;
        RECT 687.110 247.625 688.360 249.125 ;
        RECT 691.740 247.645 693.710 249.145 ;
        RECT 697.220 247.635 698.150 249.085 ;
        RECT 698.680 247.635 699.930 249.135 ;
        RECT 701.140 248.610 701.830 249.450 ;
        RECT 702.790 249.375 706.150 249.545 ;
        RECT 708.140 249.395 711.500 249.565 ;
        RECT 714.700 249.465 718.060 249.635 ;
        RECT 702.880 247.645 703.810 249.095 ;
        RECT 704.340 247.645 705.590 249.145 ;
        RECT 708.970 247.665 710.940 249.165 ;
        RECT 714.790 247.735 715.720 249.185 ;
        RECT 716.250 247.735 717.500 249.235 ;
        RECT 718.370 248.710 719.290 249.550 ;
        RECT 720.360 249.475 723.720 249.645 ;
        RECT 725.710 249.495 729.070 249.665 ;
        RECT 731.870 249.495 735.230 249.665 ;
        RECT 720.450 247.745 721.380 249.195 ;
        RECT 721.910 247.745 723.160 249.245 ;
        RECT 726.540 247.765 728.510 249.265 ;
        RECT 731.960 247.765 732.890 249.215 ;
        RECT 733.420 247.765 734.670 249.265 ;
        RECT 735.890 248.750 736.560 249.610 ;
        RECT 737.530 249.505 740.890 249.675 ;
        RECT 742.880 249.525 746.240 249.695 ;
        RECT 749.680 249.555 753.040 249.725 ;
        RECT 737.620 247.775 738.550 249.225 ;
        RECT 739.080 247.775 740.330 249.275 ;
        RECT 743.710 247.795 745.680 249.295 ;
        RECT 749.770 247.825 750.700 249.275 ;
        RECT 751.230 247.825 752.480 249.325 ;
        RECT 753.730 248.830 754.360 249.670 ;
        RECT 755.340 249.565 758.700 249.735 ;
        RECT 760.690 249.585 764.050 249.755 ;
        RECT 755.430 247.835 756.360 249.285 ;
        RECT 756.890 247.835 758.140 249.335 ;
        RECT 761.520 247.855 763.490 249.355 ;
        RECT 697.255 246.555 697.665 247.225 ;
        RECT 286.830 245.790 287.510 245.920 ;
        RECT 286.230 245.720 287.550 245.790 ;
        RECT 272.420 245.690 287.550 245.720 ;
        RECT 271.740 245.520 287.550 245.690 ;
        RECT 272.420 245.450 287.550 245.520 ;
        RECT 286.230 245.410 287.550 245.450 ;
        RECT 285.120 242.560 286.060 242.610 ;
        RECT 286.830 242.560 287.510 245.410 ;
        RECT 210.720 242.490 212.220 242.550 ;
        RECT 230.690 242.490 232.190 242.550 ;
        RECT 250.800 242.490 252.300 242.550 ;
        RECT 270.910 242.490 272.410 242.550 ;
        RECT 285.120 242.490 287.660 242.560 ;
        RECT 210.720 242.230 287.660 242.490 ;
        RECT 210.720 242.180 226.430 242.230 ;
        RECT 230.690 242.180 246.400 242.230 ;
        RECT 250.800 242.180 266.510 242.230 ;
        RECT 270.910 242.180 287.660 242.230 ;
        RECT 210.720 242.170 212.130 242.180 ;
        RECT 230.690 242.170 232.100 242.180 ;
        RECT 250.800 242.170 252.210 242.180 ;
        RECT 270.910 242.170 272.320 242.180 ;
        RECT 210.740 242.160 211.150 242.170 ;
        RECT 230.710 242.160 231.120 242.170 ;
        RECT 250.820 242.160 251.230 242.170 ;
        RECT 270.930 242.160 271.340 242.170 ;
        RECT 94.220 241.660 102.800 241.930 ;
        RECT 94.220 241.550 98.170 241.660 ;
        RECT 101.680 241.590 102.800 241.660 ;
        RECT 81.470 240.830 82.740 241.220 ;
        RECT 92.610 238.460 92.980 241.380 ;
        RECT 94.220 240.910 95.270 241.550 ;
        RECT 96.760 241.520 98.170 241.550 ;
        RECT 101.400 238.730 102.050 238.830 ;
        RECT 102.390 238.730 102.800 241.590 ;
        RECT 285.120 242.040 287.660 242.180 ;
        RECT 213.100 239.180 224.920 241.290 ;
        RECT 285.120 241.090 286.060 242.040 ;
        RECT 232.640 239.310 247.090 241.090 ;
        RECT 253.030 239.240 267.220 241.030 ;
        RECT 271.770 239.310 286.360 241.090 ;
        RECT 285.120 239.200 286.060 239.310 ;
        RECT 101.400 238.670 102.800 238.730 ;
        RECT 97.960 238.610 102.800 238.670 ;
        RECT 78.760 238.410 79.870 238.440 ;
        RECT 91.890 238.430 93.000 238.460 ;
        RECT 97.640 238.440 102.800 238.610 ;
        RECT 5.150 238.360 13.390 238.400 ;
        RECT 25.620 238.380 26.730 238.410 ;
        RECT 4.610 238.190 13.390 238.360 ;
        RECT 18.490 238.340 26.730 238.380 ;
        RECT 31.860 238.370 40.100 238.410 ;
        RECT 45.090 238.370 53.330 238.410 ;
        RECT 65.490 238.380 66.600 238.410 ;
        RECT 5.150 238.140 13.390 238.190 ;
        RECT 17.950 238.170 26.730 238.340 ;
        RECT 31.320 238.200 40.100 238.370 ;
        RECT 44.550 238.200 53.330 238.370 ;
        RECT 58.360 238.340 66.600 238.380 ;
        RECT 71.630 238.370 79.870 238.410 ;
        RECT 84.760 238.390 93.000 238.430 ;
        RECT 12.280 238.080 13.390 238.140 ;
        RECT 18.490 238.120 26.730 238.170 ;
        RECT 31.860 238.150 40.100 238.200 ;
        RECT 45.090 238.150 53.330 238.200 ;
        RECT 57.820 238.170 66.600 238.340 ;
        RECT 71.090 238.200 79.870 238.370 ;
        RECT 84.220 238.220 93.000 238.390 ;
        RECT 97.960 238.380 102.800 238.440 ;
        RECT 25.620 238.060 26.730 238.120 ;
        RECT 38.990 238.090 40.100 238.150 ;
        RECT 52.220 238.090 53.330 238.150 ;
        RECT 58.360 238.120 66.600 238.170 ;
        RECT 71.630 238.150 79.870 238.200 ;
        RECT 84.760 238.170 93.000 238.220 ;
        RECT 65.490 238.060 66.600 238.120 ;
        RECT 78.760 238.090 79.870 238.150 ;
        RECT 91.890 238.110 93.000 238.170 ;
        RECT -44.035 236.270 -43.855 236.660 ;
        RECT -51.725 236.250 -27.275 236.270 ;
        RECT -51.970 236.090 -26.880 236.250 ;
        RECT -51.970 236.080 -51.390 236.090 ;
        RECT -50.680 236.080 -50.100 236.090 ;
        RECT -49.390 236.080 -48.810 236.090 ;
        RECT -48.100 236.080 -47.520 236.090 ;
        RECT -46.810 236.080 -46.230 236.090 ;
        RECT -45.520 236.080 -44.940 236.090 ;
        RECT -44.230 236.080 -43.650 236.090 ;
        RECT -42.940 236.080 -42.360 236.090 ;
        RECT -41.650 236.080 -41.070 236.090 ;
        RECT -40.360 236.080 -39.780 236.090 ;
        RECT -39.070 236.080 -38.490 236.090 ;
        RECT -37.780 236.080 -37.200 236.090 ;
        RECT -36.490 236.080 -35.910 236.090 ;
        RECT -35.200 236.080 -34.620 236.090 ;
        RECT -33.910 236.080 -33.330 236.090 ;
        RECT -32.620 236.080 -32.040 236.090 ;
        RECT -31.330 236.080 -30.750 236.090 ;
        RECT -30.040 236.080 -29.460 236.090 ;
        RECT -28.750 236.080 -28.170 236.090 ;
        RECT -27.460 236.080 -26.880 236.090 ;
        RECT 12.300 236.050 22.080 237.000 ;
        RECT 45.190 236.010 53.170 237.150 ;
        RECT 70.820 235.940 78.480 237.080 ;
        RECT 84.810 236.030 92.070 237.170 ;
        RECT 101.400 237.060 102.050 238.380 ;
        RECT 102.390 238.350 102.800 238.380 ;
        RECT 97.030 235.950 102.620 237.060 ;
        RECT -53.080 231.975 -52.910 235.075 ;
        RECT -52.410 232.535 -52.240 234.155 ;
        RECT -49.830 232.535 -49.660 234.155 ;
        RECT -47.250 232.535 -47.080 234.155 ;
        RECT -44.670 232.535 -44.500 234.155 ;
        RECT -42.090 232.535 -41.920 234.155 ;
        RECT -39.510 232.535 -39.340 234.155 ;
        RECT -36.930 232.535 -36.760 234.155 ;
        RECT -34.350 232.535 -34.180 234.155 ;
        RECT -31.770 232.535 -31.600 234.155 ;
        RECT -29.190 232.535 -29.020 234.155 ;
        RECT -26.610 232.535 -26.440 234.155 ;
        RECT -25.940 231.975 -25.770 235.075 ;
        RECT -46.090 230.105 -32.760 230.275 ;
        RECT -46.010 224.550 -32.520 227.170 ;
        RECT -43.925 224.120 -43.745 224.550 ;
        RECT -51.615 224.100 -27.165 224.120 ;
        RECT -51.860 223.940 -26.770 224.100 ;
        RECT -51.860 223.930 -51.280 223.940 ;
        RECT -50.570 223.930 -49.990 223.940 ;
        RECT -49.280 223.930 -48.700 223.940 ;
        RECT -47.990 223.930 -47.410 223.940 ;
        RECT -46.700 223.930 -46.120 223.940 ;
        RECT -45.410 223.930 -44.830 223.940 ;
        RECT -44.120 223.930 -43.540 223.940 ;
        RECT -42.830 223.930 -42.250 223.940 ;
        RECT -41.540 223.930 -40.960 223.940 ;
        RECT -40.250 223.930 -39.670 223.940 ;
        RECT -38.960 223.930 -38.380 223.940 ;
        RECT -37.670 223.930 -37.090 223.940 ;
        RECT -36.380 223.930 -35.800 223.940 ;
        RECT -35.090 223.930 -34.510 223.940 ;
        RECT -33.800 223.930 -33.220 223.940 ;
        RECT -32.510 223.930 -31.930 223.940 ;
        RECT -31.220 223.930 -30.640 223.940 ;
        RECT -29.930 223.930 -29.350 223.940 ;
        RECT -28.640 223.930 -28.060 223.940 ;
        RECT -27.350 223.930 -26.770 223.940 ;
        RECT -52.970 219.825 -52.800 222.925 ;
        RECT -52.300 220.385 -52.130 222.005 ;
        RECT -49.720 220.385 -49.550 222.005 ;
        RECT -47.140 220.385 -46.970 222.005 ;
        RECT -44.560 220.385 -44.390 222.005 ;
        RECT -41.980 220.385 -41.810 222.005 ;
        RECT -39.400 220.385 -39.230 222.005 ;
        RECT -36.820 220.385 -36.650 222.005 ;
        RECT -34.240 220.385 -34.070 222.005 ;
        RECT -31.660 220.385 -31.490 222.005 ;
        RECT -29.080 220.385 -28.910 222.005 ;
        RECT -26.500 220.385 -26.330 222.005 ;
        RECT -25.830 219.825 -25.660 222.925 ;
        RECT -45.980 217.955 -32.650 218.125 ;
        RECT -46.010 137.145 -32.520 139.560 ;
        RECT -46.020 136.975 -32.520 137.145 ;
        RECT -46.010 136.940 -32.520 136.975 ;
        RECT -43.965 136.470 -43.785 136.940 ;
        RECT -51.655 136.450 -27.205 136.470 ;
        RECT -51.900 136.290 -26.810 136.450 ;
        RECT -51.900 136.280 -51.320 136.290 ;
        RECT -50.610 136.280 -50.030 136.290 ;
        RECT -49.320 136.280 -48.740 136.290 ;
        RECT -48.030 136.280 -47.450 136.290 ;
        RECT -46.740 136.280 -46.160 136.290 ;
        RECT -45.450 136.280 -44.870 136.290 ;
        RECT -44.160 136.280 -43.580 136.290 ;
        RECT -42.870 136.280 -42.290 136.290 ;
        RECT -41.580 136.280 -41.000 136.290 ;
        RECT -40.290 136.280 -39.710 136.290 ;
        RECT -39.000 136.280 -38.420 136.290 ;
        RECT -37.710 136.280 -37.130 136.290 ;
        RECT -36.420 136.280 -35.840 136.290 ;
        RECT -35.130 136.280 -34.550 136.290 ;
        RECT -33.840 136.280 -33.260 136.290 ;
        RECT -32.550 136.280 -31.970 136.290 ;
        RECT -31.260 136.280 -30.680 136.290 ;
        RECT -29.970 136.280 -29.390 136.290 ;
        RECT -28.680 136.280 -28.100 136.290 ;
        RECT -27.390 136.280 -26.810 136.290 ;
        RECT -53.010 132.175 -52.840 135.275 ;
        RECT -52.340 132.735 -52.170 134.355 ;
        RECT -49.760 132.735 -49.590 134.355 ;
        RECT -47.180 132.735 -47.010 134.355 ;
        RECT -44.600 132.735 -44.430 134.355 ;
        RECT -42.020 132.735 -41.850 134.355 ;
        RECT -39.440 132.735 -39.270 134.355 ;
        RECT -36.860 132.735 -36.690 134.355 ;
        RECT -34.280 132.735 -34.110 134.355 ;
        RECT -31.700 132.735 -31.530 134.355 ;
        RECT -29.120 132.735 -28.950 134.355 ;
        RECT -26.540 132.735 -26.370 134.355 ;
        RECT -25.870 132.175 -25.700 135.275 ;
        RECT -46.020 130.305 -32.690 130.475 ;
        RECT -45.890 17.705 -32.400 20.120 ;
        RECT -45.900 17.535 -32.400 17.705 ;
        RECT -45.890 17.500 -32.400 17.535 ;
        RECT -43.845 17.030 -43.665 17.500 ;
        RECT -51.535 17.010 -27.085 17.030 ;
        RECT -51.780 16.850 -26.690 17.010 ;
        RECT -51.780 16.840 -51.200 16.850 ;
        RECT -50.490 16.840 -49.910 16.850 ;
        RECT -49.200 16.840 -48.620 16.850 ;
        RECT -47.910 16.840 -47.330 16.850 ;
        RECT -46.620 16.840 -46.040 16.850 ;
        RECT -45.330 16.840 -44.750 16.850 ;
        RECT -44.040 16.840 -43.460 16.850 ;
        RECT -42.750 16.840 -42.170 16.850 ;
        RECT -41.460 16.840 -40.880 16.850 ;
        RECT -40.170 16.840 -39.590 16.850 ;
        RECT -38.880 16.840 -38.300 16.850 ;
        RECT -37.590 16.840 -37.010 16.850 ;
        RECT -36.300 16.840 -35.720 16.850 ;
        RECT -35.010 16.840 -34.430 16.850 ;
        RECT -33.720 16.840 -33.140 16.850 ;
        RECT -32.430 16.840 -31.850 16.850 ;
        RECT -31.140 16.840 -30.560 16.850 ;
        RECT -29.850 16.840 -29.270 16.850 ;
        RECT -28.560 16.840 -27.980 16.850 ;
        RECT -27.270 16.840 -26.690 16.850 ;
        RECT -52.890 12.735 -52.720 15.835 ;
        RECT -52.220 13.295 -52.050 14.915 ;
        RECT -49.640 13.295 -49.470 14.915 ;
        RECT -47.060 13.295 -46.890 14.915 ;
        RECT -44.480 13.295 -44.310 14.915 ;
        RECT -41.900 13.295 -41.730 14.915 ;
        RECT -39.320 13.295 -39.150 14.915 ;
        RECT -36.740 13.295 -36.570 14.915 ;
        RECT -34.160 13.295 -33.990 14.915 ;
        RECT -31.580 13.295 -31.410 14.915 ;
        RECT -29.000 13.295 -28.830 14.915 ;
        RECT -26.420 13.295 -26.250 14.915 ;
        RECT -25.750 12.735 -25.580 15.835 ;
        RECT -45.900 10.865 -32.570 11.035 ;
      LAYER mcon ;
        RECT 363.230 372.070 363.400 372.240 ;
        RECT 363.590 372.070 363.760 372.240 ;
        RECT 363.950 372.070 364.120 372.240 ;
        RECT 402.420 372.220 403.670 372.750 ;
        RECT 356.690 369.865 356.860 370.035 ;
        RECT 356.690 369.505 356.860 369.675 ;
        RECT 359.980 369.865 360.150 370.035 ;
        RECT 359.980 369.505 360.150 369.675 ;
        RECT 363.270 369.865 363.440 370.035 ;
        RECT 215.390 367.450 226.000 368.340 ;
        RECT 235.430 367.440 246.040 368.330 ;
        RECT 255.490 367.440 266.100 368.330 ;
        RECT 275.540 367.440 286.150 368.330 ;
        RECT 363.270 369.505 363.440 369.675 ;
        RECT 366.560 369.865 366.730 370.035 ;
        RECT 369.850 369.865 370.020 370.035 ;
        RECT 366.560 369.505 366.730 369.675 ;
        RECT 369.850 369.505 370.020 369.675 ;
        RECT 376.010 369.765 376.180 369.935 ;
        RECT 376.010 369.405 376.180 369.575 ;
        RECT 382.590 369.765 382.760 369.935 ;
        RECT 389.170 369.765 389.340 369.935 ;
        RECT 395.260 369.835 395.430 370.005 ;
        RECT 382.590 369.405 382.760 369.575 ;
        RECT 389.170 369.405 389.340 369.575 ;
        RECT 395.260 369.475 395.430 369.645 ;
        RECT 398.550 369.835 398.720 370.005 ;
        RECT 398.550 369.475 398.720 369.645 ;
        RECT 401.840 369.835 402.010 370.005 ;
        RECT 401.840 369.475 402.010 369.645 ;
        RECT 405.130 369.835 405.300 370.005 ;
        RECT 408.420 369.835 408.590 370.005 ;
        RECT 405.130 369.475 405.300 369.645 ;
        RECT 408.420 369.475 408.590 369.645 ;
        RECT 212.215 365.970 212.385 366.140 ;
        RECT 212.575 365.970 212.745 366.140 ;
        RECT 215.685 365.970 215.855 366.140 ;
        RECT 216.045 365.970 216.215 366.140 ;
        RECT 219.155 365.970 219.325 366.140 ;
        RECT 219.515 365.970 219.685 366.140 ;
        RECT 222.625 365.970 222.795 366.140 ;
        RECT 222.985 365.970 223.155 366.140 ;
        RECT 226.095 365.970 226.265 366.140 ;
        RECT 226.455 365.970 226.625 366.140 ;
        RECT 232.255 365.960 232.425 366.130 ;
        RECT 232.615 365.960 232.785 366.130 ;
        RECT 235.725 365.960 235.895 366.130 ;
        RECT 236.085 365.960 236.255 366.130 ;
        RECT 239.195 365.960 239.365 366.130 ;
        RECT 239.555 365.960 239.725 366.130 ;
        RECT 242.665 365.960 242.835 366.130 ;
        RECT 243.025 365.960 243.195 366.130 ;
        RECT 246.135 365.960 246.305 366.130 ;
        RECT 246.495 365.960 246.665 366.130 ;
        RECT 252.315 365.960 252.485 366.130 ;
        RECT 252.675 365.960 252.845 366.130 ;
        RECT 255.785 365.960 255.955 366.130 ;
        RECT 256.145 365.960 256.315 366.130 ;
        RECT 259.255 365.960 259.425 366.130 ;
        RECT 259.615 365.960 259.785 366.130 ;
        RECT 262.725 365.960 262.895 366.130 ;
        RECT 263.085 365.960 263.255 366.130 ;
        RECT 266.195 365.960 266.365 366.130 ;
        RECT 266.555 365.960 266.725 366.130 ;
        RECT 272.365 365.960 272.535 366.130 ;
        RECT 272.725 365.960 272.895 366.130 ;
        RECT 275.835 365.960 276.005 366.130 ;
        RECT 276.195 365.960 276.365 366.130 ;
        RECT 279.305 365.960 279.475 366.130 ;
        RECT 279.665 365.960 279.835 366.130 ;
        RECT 282.775 365.960 282.945 366.130 ;
        RECT 283.135 365.960 283.305 366.130 ;
        RECT 286.245 365.960 286.415 366.130 ;
        RECT 286.605 365.960 286.775 366.130 ;
        RECT 212.215 362.680 212.385 362.850 ;
        RECT 212.575 362.680 212.745 362.850 ;
        RECT 215.685 362.680 215.855 362.850 ;
        RECT 216.045 362.680 216.215 362.850 ;
        RECT 219.155 362.680 219.325 362.850 ;
        RECT 219.515 362.680 219.685 362.850 ;
        RECT 222.625 362.680 222.795 362.850 ;
        RECT 222.985 362.680 223.155 362.850 ;
        RECT 226.095 362.680 226.265 362.850 ;
        RECT 226.455 362.680 226.625 362.850 ;
        RECT -44.420 358.005 -34.530 359.615 ;
        RECT -51.775 357.460 -51.605 357.630 ;
        RECT -50.485 357.460 -50.315 357.630 ;
        RECT -49.195 357.460 -49.025 357.630 ;
        RECT -47.905 357.460 -47.735 357.630 ;
        RECT -46.615 357.460 -46.445 357.630 ;
        RECT -45.325 357.460 -45.155 357.630 ;
        RECT -44.035 357.460 -43.865 357.630 ;
        RECT -42.745 357.460 -42.575 357.630 ;
        RECT -41.455 357.460 -41.285 357.630 ;
        RECT -40.165 357.460 -39.995 357.630 ;
        RECT -38.875 357.460 -38.705 357.630 ;
        RECT -37.585 357.460 -37.415 357.630 ;
        RECT -36.295 357.460 -36.125 357.630 ;
        RECT -35.005 357.460 -34.835 357.630 ;
        RECT -33.715 357.460 -33.545 357.630 ;
        RECT -32.425 357.460 -32.255 357.630 ;
        RECT -31.135 357.460 -30.965 357.630 ;
        RECT -29.845 357.460 -29.675 357.630 ;
        RECT -28.555 357.460 -28.385 357.630 ;
        RECT -27.265 357.460 -27.095 357.630 ;
        RECT -52.420 355.180 -52.250 355.350 ;
        RECT -52.420 354.820 -52.250 354.990 ;
        RECT -52.420 354.460 -52.250 354.630 ;
        RECT -52.420 354.100 -52.250 354.270 ;
        RECT -49.840 355.180 -49.670 355.350 ;
        RECT -49.840 354.820 -49.670 354.990 ;
        RECT -49.840 354.460 -49.670 354.630 ;
        RECT -49.840 354.100 -49.670 354.270 ;
        RECT -47.260 355.180 -47.090 355.350 ;
        RECT -47.260 354.820 -47.090 354.990 ;
        RECT -47.260 354.460 -47.090 354.630 ;
        RECT -47.260 354.100 -47.090 354.270 ;
        RECT -44.680 355.180 -44.510 355.350 ;
        RECT -44.680 354.820 -44.510 354.990 ;
        RECT -44.680 354.460 -44.510 354.630 ;
        RECT -44.680 354.100 -44.510 354.270 ;
        RECT -42.100 355.180 -41.930 355.350 ;
        RECT -42.100 354.820 -41.930 354.990 ;
        RECT -42.100 354.460 -41.930 354.630 ;
        RECT -42.100 354.100 -41.930 354.270 ;
        RECT -39.520 355.180 -39.350 355.350 ;
        RECT -39.520 354.820 -39.350 354.990 ;
        RECT -39.520 354.460 -39.350 354.630 ;
        RECT -39.520 354.100 -39.350 354.270 ;
        RECT -36.940 355.180 -36.770 355.350 ;
        RECT -36.940 354.820 -36.770 354.990 ;
        RECT -36.940 354.460 -36.770 354.630 ;
        RECT -36.940 354.100 -36.770 354.270 ;
        RECT -34.360 355.180 -34.190 355.350 ;
        RECT -34.360 354.820 -34.190 354.990 ;
        RECT -34.360 354.460 -34.190 354.630 ;
        RECT -34.360 354.100 -34.190 354.270 ;
        RECT -31.780 355.180 -31.610 355.350 ;
        RECT -31.780 354.820 -31.610 354.990 ;
        RECT -31.780 354.460 -31.610 354.630 ;
        RECT -31.780 354.100 -31.610 354.270 ;
        RECT -29.200 355.180 -29.030 355.350 ;
        RECT -29.200 354.820 -29.030 354.990 ;
        RECT -29.200 354.460 -29.030 354.630 ;
        RECT -29.200 354.100 -29.030 354.270 ;
        RECT -26.620 355.180 -26.450 355.350 ;
        RECT -26.620 354.820 -26.450 354.990 ;
        RECT -26.620 354.460 -26.450 354.630 ;
        RECT -26.620 354.100 -26.450 354.270 ;
        RECT 232.255 362.670 232.425 362.840 ;
        RECT 232.615 362.670 232.785 362.840 ;
        RECT 235.725 362.670 235.895 362.840 ;
        RECT 236.085 362.670 236.255 362.840 ;
        RECT 239.195 362.670 239.365 362.840 ;
        RECT 239.555 362.670 239.725 362.840 ;
        RECT 242.665 362.670 242.835 362.840 ;
        RECT 243.025 362.670 243.195 362.840 ;
        RECT 246.135 362.670 246.305 362.840 ;
        RECT 246.495 362.670 246.665 362.840 ;
        RECT 212.215 359.390 212.385 359.560 ;
        RECT 212.575 359.390 212.745 359.560 ;
        RECT 215.685 359.390 215.855 359.560 ;
        RECT 216.045 359.390 216.215 359.560 ;
        RECT 219.155 359.390 219.325 359.560 ;
        RECT 219.515 359.390 219.685 359.560 ;
        RECT 222.625 359.390 222.795 359.560 ;
        RECT 222.985 359.390 223.155 359.560 ;
        RECT 226.095 359.390 226.265 359.560 ;
        RECT 226.455 359.390 226.625 359.560 ;
        RECT 212.215 356.100 212.385 356.270 ;
        RECT 212.575 356.100 212.745 356.270 ;
        RECT 215.685 356.100 215.855 356.270 ;
        RECT 216.045 356.100 216.215 356.270 ;
        RECT 219.155 356.100 219.325 356.270 ;
        RECT 219.515 356.100 219.685 356.270 ;
        RECT 222.625 356.100 222.795 356.270 ;
        RECT 222.985 356.100 223.155 356.270 ;
        RECT 226.095 356.100 226.265 356.270 ;
        RECT 226.455 356.100 226.625 356.270 ;
        RECT 252.315 362.670 252.485 362.840 ;
        RECT 252.675 362.670 252.845 362.840 ;
        RECT 255.785 362.670 255.955 362.840 ;
        RECT 256.145 362.670 256.315 362.840 ;
        RECT 259.255 362.670 259.425 362.840 ;
        RECT 259.615 362.670 259.785 362.840 ;
        RECT 262.725 362.670 262.895 362.840 ;
        RECT 263.085 362.670 263.255 362.840 ;
        RECT 266.195 362.670 266.365 362.840 ;
        RECT 266.555 362.670 266.725 362.840 ;
        RECT 232.255 359.380 232.425 359.550 ;
        RECT 232.615 359.380 232.785 359.550 ;
        RECT 235.725 359.380 235.895 359.550 ;
        RECT 236.085 359.380 236.255 359.550 ;
        RECT 239.195 359.380 239.365 359.550 ;
        RECT 239.555 359.380 239.725 359.550 ;
        RECT 242.665 359.380 242.835 359.550 ;
        RECT 243.025 359.380 243.195 359.550 ;
        RECT 246.135 359.380 246.305 359.550 ;
        RECT 246.495 359.380 246.665 359.550 ;
        RECT 232.255 356.090 232.425 356.260 ;
        RECT 232.615 356.090 232.785 356.260 ;
        RECT 235.725 356.090 235.895 356.260 ;
        RECT 236.085 356.090 236.255 356.260 ;
        RECT 239.195 356.090 239.365 356.260 ;
        RECT 239.555 356.090 239.725 356.260 ;
        RECT 242.665 356.090 242.835 356.260 ;
        RECT 243.025 356.090 243.195 356.260 ;
        RECT 246.135 356.090 246.305 356.260 ;
        RECT 246.495 356.090 246.665 356.260 ;
        RECT 212.215 352.810 212.385 352.980 ;
        RECT 212.575 352.810 212.745 352.980 ;
        RECT 215.685 352.810 215.855 352.980 ;
        RECT 216.045 352.810 216.215 352.980 ;
        RECT 219.155 352.810 219.325 352.980 ;
        RECT 219.515 352.810 219.685 352.980 ;
        RECT 222.625 352.810 222.795 352.980 ;
        RECT 222.985 352.810 223.155 352.980 ;
        RECT 226.095 352.810 226.265 352.980 ;
        RECT 226.455 352.810 226.625 352.980 ;
        RECT 272.365 362.670 272.535 362.840 ;
        RECT 272.725 362.670 272.895 362.840 ;
        RECT 275.835 362.670 276.005 362.840 ;
        RECT 276.195 362.670 276.365 362.840 ;
        RECT 279.305 362.670 279.475 362.840 ;
        RECT 279.665 362.670 279.835 362.840 ;
        RECT 282.775 362.670 282.945 362.840 ;
        RECT 283.135 362.670 283.305 362.840 ;
        RECT 286.245 362.670 286.415 362.840 ;
        RECT 286.605 362.670 286.775 362.840 ;
        RECT 252.315 359.380 252.485 359.550 ;
        RECT 252.675 359.380 252.845 359.550 ;
        RECT 255.785 359.380 255.955 359.550 ;
        RECT 256.145 359.380 256.315 359.550 ;
        RECT 259.255 359.380 259.425 359.550 ;
        RECT 259.615 359.380 259.785 359.550 ;
        RECT 262.725 359.380 262.895 359.550 ;
        RECT 263.085 359.380 263.255 359.550 ;
        RECT 266.195 359.380 266.365 359.550 ;
        RECT 266.555 359.380 266.725 359.550 ;
        RECT 252.315 356.090 252.485 356.260 ;
        RECT 252.675 356.090 252.845 356.260 ;
        RECT 255.785 356.090 255.955 356.260 ;
        RECT 256.145 356.090 256.315 356.260 ;
        RECT 259.255 356.090 259.425 356.260 ;
        RECT 259.615 356.090 259.785 356.260 ;
        RECT 262.725 356.090 262.895 356.260 ;
        RECT 263.085 356.090 263.255 356.260 ;
        RECT 266.195 356.090 266.365 356.260 ;
        RECT 266.555 356.090 266.725 356.260 ;
        RECT 232.255 352.800 232.425 352.970 ;
        RECT 232.615 352.800 232.785 352.970 ;
        RECT 235.725 352.800 235.895 352.970 ;
        RECT 236.085 352.800 236.255 352.970 ;
        RECT 239.195 352.800 239.365 352.970 ;
        RECT 239.555 352.800 239.725 352.970 ;
        RECT 242.665 352.800 242.835 352.970 ;
        RECT 243.025 352.800 243.195 352.970 ;
        RECT 246.135 352.800 246.305 352.970 ;
        RECT 246.495 352.800 246.665 352.970 ;
        RECT 355.455 364.695 355.625 364.865 ;
        RECT 355.455 364.335 355.625 364.505 ;
        RECT 355.455 363.975 355.625 364.145 ;
        RECT 355.455 363.615 355.625 363.785 ;
        RECT 356.550 365.295 356.720 365.465 ;
        RECT 356.550 364.935 356.720 365.105 ;
        RECT 355.455 363.255 355.625 363.425 ;
        RECT 355.455 362.895 355.625 363.065 ;
        RECT 355.455 362.535 355.625 362.705 ;
        RECT 355.455 362.175 355.625 362.345 ;
        RECT 355.455 361.815 355.625 361.985 ;
        RECT 355.455 361.455 355.625 361.625 ;
        RECT 355.455 361.095 355.625 361.265 ;
        RECT 355.455 360.735 355.625 360.905 ;
        RECT 355.455 360.375 355.625 360.545 ;
        RECT 355.455 360.015 355.625 360.185 ;
        RECT 355.455 359.655 355.625 359.825 ;
        RECT 272.365 359.380 272.535 359.550 ;
        RECT 272.725 359.380 272.895 359.550 ;
        RECT 275.835 359.380 276.005 359.550 ;
        RECT 276.195 359.380 276.365 359.550 ;
        RECT 279.305 359.380 279.475 359.550 ;
        RECT 279.665 359.380 279.835 359.550 ;
        RECT 282.775 359.380 282.945 359.550 ;
        RECT 283.135 359.380 283.305 359.550 ;
        RECT 286.245 359.380 286.415 359.550 ;
        RECT 286.605 359.380 286.775 359.550 ;
        RECT 355.455 359.295 355.625 359.465 ;
        RECT 272.365 356.090 272.535 356.260 ;
        RECT 272.725 356.090 272.895 356.260 ;
        RECT 275.835 356.090 276.005 356.260 ;
        RECT 276.195 356.090 276.365 356.260 ;
        RECT 279.305 356.090 279.475 356.260 ;
        RECT 279.665 356.090 279.835 356.260 ;
        RECT 282.775 356.090 282.945 356.260 ;
        RECT 283.135 356.090 283.305 356.260 ;
        RECT 286.245 356.090 286.415 356.260 ;
        RECT 286.605 356.090 286.775 356.260 ;
        RECT 252.315 352.800 252.485 352.970 ;
        RECT 252.675 352.800 252.845 352.970 ;
        RECT 255.785 352.800 255.955 352.970 ;
        RECT 256.145 352.800 256.315 352.970 ;
        RECT 259.255 352.800 259.425 352.970 ;
        RECT 259.615 352.800 259.785 352.970 ;
        RECT 262.725 352.800 262.895 352.970 ;
        RECT 263.085 352.800 263.255 352.970 ;
        RECT 266.195 352.800 266.365 352.970 ;
        RECT 266.555 352.800 266.725 352.970 ;
        RECT 355.455 358.935 355.625 359.105 ;
        RECT 355.455 358.575 355.625 358.745 ;
        RECT 355.455 358.215 355.625 358.385 ;
        RECT 355.455 357.855 355.625 358.025 ;
        RECT 355.455 357.495 355.625 357.665 ;
        RECT 355.455 357.135 355.625 357.305 ;
        RECT 355.455 356.775 355.625 356.945 ;
        RECT 355.455 356.415 355.625 356.585 ;
        RECT 355.455 356.055 355.625 356.225 ;
        RECT 355.455 355.695 355.625 355.865 ;
        RECT 355.455 355.335 355.625 355.505 ;
        RECT 355.455 354.975 355.625 355.145 ;
        RECT 355.455 354.615 355.625 354.785 ;
        RECT 355.455 354.255 355.625 354.425 ;
        RECT 355.455 353.895 355.625 354.065 ;
        RECT 355.455 353.535 355.625 353.705 ;
        RECT 355.455 353.175 355.625 353.345 ;
        RECT 272.365 352.800 272.535 352.970 ;
        RECT 272.725 352.800 272.895 352.970 ;
        RECT 275.835 352.800 276.005 352.970 ;
        RECT 276.195 352.800 276.365 352.970 ;
        RECT 279.305 352.800 279.475 352.970 ;
        RECT 279.665 352.800 279.835 352.970 ;
        RECT 282.775 352.800 282.945 352.970 ;
        RECT 283.135 352.800 283.305 352.970 ;
        RECT 286.245 352.800 286.415 352.970 ;
        RECT 286.605 352.800 286.775 352.970 ;
        RECT 355.455 352.815 355.625 352.985 ;
        RECT 212.215 349.520 212.385 349.690 ;
        RECT 212.575 349.520 212.745 349.690 ;
        RECT 215.685 349.520 215.855 349.690 ;
        RECT 216.045 349.520 216.215 349.690 ;
        RECT 219.155 349.520 219.325 349.690 ;
        RECT 219.515 349.520 219.685 349.690 ;
        RECT 222.625 349.520 222.795 349.690 ;
        RECT 222.985 349.520 223.155 349.690 ;
        RECT 226.095 349.520 226.265 349.690 ;
        RECT 226.455 349.520 226.625 349.690 ;
        RECT 232.255 349.510 232.425 349.680 ;
        RECT 232.615 349.510 232.785 349.680 ;
        RECT 235.725 349.510 235.895 349.680 ;
        RECT 236.085 349.510 236.255 349.680 ;
        RECT 239.195 349.510 239.365 349.680 ;
        RECT 239.555 349.510 239.725 349.680 ;
        RECT 242.665 349.510 242.835 349.680 ;
        RECT 243.025 349.510 243.195 349.680 ;
        RECT 246.135 349.510 246.305 349.680 ;
        RECT 246.495 349.510 246.665 349.680 ;
        RECT 252.315 349.510 252.485 349.680 ;
        RECT 252.675 349.510 252.845 349.680 ;
        RECT 255.785 349.510 255.955 349.680 ;
        RECT 256.145 349.510 256.315 349.680 ;
        RECT 259.255 349.510 259.425 349.680 ;
        RECT 259.615 349.510 259.785 349.680 ;
        RECT 262.725 349.510 262.895 349.680 ;
        RECT 263.085 349.510 263.255 349.680 ;
        RECT 266.195 349.510 266.365 349.680 ;
        RECT 266.555 349.510 266.725 349.680 ;
        RECT 272.365 349.510 272.535 349.680 ;
        RECT 272.725 349.510 272.895 349.680 ;
        RECT 275.835 349.510 276.005 349.680 ;
        RECT 276.195 349.510 276.365 349.680 ;
        RECT 279.305 349.510 279.475 349.680 ;
        RECT 279.665 349.510 279.835 349.680 ;
        RECT 282.775 349.510 282.945 349.680 ;
        RECT 283.135 349.510 283.305 349.680 ;
        RECT 286.245 349.510 286.415 349.680 ;
        RECT 286.605 349.510 286.775 349.680 ;
        RECT 355.455 352.455 355.625 352.625 ;
        RECT 355.455 352.095 355.625 352.265 ;
        RECT 356.550 361.825 356.720 361.995 ;
        RECT 356.550 361.465 356.720 361.635 ;
        RECT 356.550 358.355 356.720 358.525 ;
        RECT 356.550 357.995 356.720 358.165 ;
        RECT 356.550 354.885 356.720 355.055 ;
        RECT 356.550 354.525 356.720 354.695 ;
        RECT 356.550 351.415 356.720 351.585 ;
        RECT 359.840 365.295 360.010 365.465 ;
        RECT 359.840 364.935 360.010 365.105 ;
        RECT 359.840 361.825 360.010 361.995 ;
        RECT 359.840 361.465 360.010 361.635 ;
        RECT 359.840 358.355 360.010 358.525 ;
        RECT 359.840 357.995 360.010 358.165 ;
        RECT 359.840 354.885 360.010 355.055 ;
        RECT 359.840 354.525 360.010 354.695 ;
        RECT 359.840 351.415 360.010 351.585 ;
        RECT 356.550 351.055 356.720 351.225 ;
        RECT 288.875 348.135 289.045 348.305 ;
        RECT 215.350 346.460 225.960 347.350 ;
        RECT 235.320 346.460 245.930 347.350 ;
        RECT 255.430 346.460 266.040 347.350 ;
        RECT 275.540 346.460 286.150 347.350 ;
        RECT 288.875 347.775 289.045 347.945 ;
        RECT 288.875 347.415 289.045 347.585 ;
        RECT 363.130 365.295 363.300 365.465 ;
        RECT 363.130 364.935 363.300 365.105 ;
        RECT 363.130 361.825 363.300 361.995 ;
        RECT 363.130 361.465 363.300 361.635 ;
        RECT 363.130 358.355 363.300 358.525 ;
        RECT 363.130 357.995 363.300 358.165 ;
        RECT 363.130 354.885 363.300 355.055 ;
        RECT 363.130 354.525 363.300 354.695 ;
        RECT 363.130 351.415 363.300 351.585 ;
        RECT 366.420 365.295 366.590 365.465 ;
        RECT 369.710 365.295 369.880 365.465 ;
        RECT 366.420 364.935 366.590 365.105 ;
        RECT 366.420 361.825 366.590 361.995 ;
        RECT 366.420 361.465 366.590 361.635 ;
        RECT 366.420 358.355 366.590 358.525 ;
        RECT 366.420 357.995 366.590 358.165 ;
        RECT 366.420 354.885 366.590 355.055 ;
        RECT 366.420 354.525 366.590 354.695 ;
        RECT 366.420 351.415 366.590 351.585 ;
        RECT 369.710 364.935 369.880 365.105 ;
        RECT 369.710 361.825 369.880 361.995 ;
        RECT 369.710 361.465 369.880 361.635 ;
        RECT 369.710 358.355 369.880 358.525 ;
        RECT 369.710 357.995 369.880 358.165 ;
        RECT 369.710 354.885 369.880 355.055 ;
        RECT 369.710 354.525 369.880 354.695 ;
        RECT 359.840 351.055 360.010 351.225 ;
        RECT 363.130 351.055 363.300 351.225 ;
        RECT 366.420 351.055 366.590 351.225 ;
        RECT 369.710 351.415 369.880 351.585 ;
        RECT 374.775 364.595 374.945 364.765 ;
        RECT 374.775 364.235 374.945 364.405 ;
        RECT 374.775 363.875 374.945 364.045 ;
        RECT 374.775 363.515 374.945 363.685 ;
        RECT 374.775 363.155 374.945 363.325 ;
        RECT 374.775 362.795 374.945 362.965 ;
        RECT 374.775 362.435 374.945 362.605 ;
        RECT 374.775 362.075 374.945 362.245 ;
        RECT 374.775 361.715 374.945 361.885 ;
        RECT 374.775 361.355 374.945 361.525 ;
        RECT 374.775 360.995 374.945 361.165 ;
        RECT 374.775 360.635 374.945 360.805 ;
        RECT 374.775 360.275 374.945 360.445 ;
        RECT 374.775 359.915 374.945 360.085 ;
        RECT 374.775 359.555 374.945 359.725 ;
        RECT 374.775 359.195 374.945 359.365 ;
        RECT 374.775 358.835 374.945 359.005 ;
        RECT 374.775 358.475 374.945 358.645 ;
        RECT 374.775 358.115 374.945 358.285 ;
        RECT 374.775 357.755 374.945 357.925 ;
        RECT 374.775 357.395 374.945 357.565 ;
        RECT 374.775 357.035 374.945 357.205 ;
        RECT 374.775 356.675 374.945 356.845 ;
        RECT 374.775 356.315 374.945 356.485 ;
        RECT 374.775 355.955 374.945 356.125 ;
        RECT 374.775 355.595 374.945 355.765 ;
        RECT 374.775 355.235 374.945 355.405 ;
        RECT 374.775 354.875 374.945 355.045 ;
        RECT 374.775 354.515 374.945 354.685 ;
        RECT 374.775 354.155 374.945 354.325 ;
        RECT 374.775 353.795 374.945 353.965 ;
        RECT 374.775 353.435 374.945 353.605 ;
        RECT 374.775 353.075 374.945 353.245 ;
        RECT 374.775 352.715 374.945 352.885 ;
        RECT 374.775 352.355 374.945 352.525 ;
        RECT 374.775 351.995 374.945 352.165 ;
        RECT 375.870 365.195 376.040 365.365 ;
        RECT 375.870 364.835 376.040 365.005 ;
        RECT 375.870 361.725 376.040 361.895 ;
        RECT 375.870 361.365 376.040 361.535 ;
        RECT 375.870 358.255 376.040 358.425 ;
        RECT 375.870 357.895 376.040 358.065 ;
        RECT 375.870 354.785 376.040 354.955 ;
        RECT 375.870 354.425 376.040 354.595 ;
        RECT 375.870 351.315 376.040 351.485 ;
        RECT 382.450 365.195 382.620 365.365 ;
        RECT 389.030 365.195 389.200 365.365 ;
        RECT 382.450 364.835 382.620 365.005 ;
        RECT 382.450 361.725 382.620 361.895 ;
        RECT 382.450 361.365 382.620 361.535 ;
        RECT 382.450 358.255 382.620 358.425 ;
        RECT 382.450 357.895 382.620 358.065 ;
        RECT 382.450 354.785 382.620 354.955 ;
        RECT 382.450 354.425 382.620 354.595 ;
        RECT 382.450 351.315 382.620 351.485 ;
        RECT 369.710 351.055 369.880 351.225 ;
        RECT 389.030 364.835 389.200 365.005 ;
        RECT 389.030 361.725 389.200 361.895 ;
        RECT 389.030 361.365 389.200 361.535 ;
        RECT 389.030 358.255 389.200 358.425 ;
        RECT 389.030 357.895 389.200 358.065 ;
        RECT 389.030 354.785 389.200 354.955 ;
        RECT 389.030 354.425 389.200 354.595 ;
        RECT 389.030 351.315 389.200 351.485 ;
        RECT 375.870 350.955 376.040 351.125 ;
        RECT 212.175 344.980 212.345 345.150 ;
        RECT 212.535 344.980 212.705 345.150 ;
        RECT 215.645 344.980 215.815 345.150 ;
        RECT 216.005 344.980 216.175 345.150 ;
        RECT 219.115 344.980 219.285 345.150 ;
        RECT 219.475 344.980 219.645 345.150 ;
        RECT 222.585 344.980 222.755 345.150 ;
        RECT 222.945 344.980 223.115 345.150 ;
        RECT 226.055 344.980 226.225 345.150 ;
        RECT 226.415 344.980 226.585 345.150 ;
        RECT 232.145 344.980 232.315 345.150 ;
        RECT 232.505 344.980 232.675 345.150 ;
        RECT 235.615 344.980 235.785 345.150 ;
        RECT 235.975 344.980 236.145 345.150 ;
        RECT 239.085 344.980 239.255 345.150 ;
        RECT 239.445 344.980 239.615 345.150 ;
        RECT 242.555 344.980 242.725 345.150 ;
        RECT 242.915 344.980 243.085 345.150 ;
        RECT 246.025 344.980 246.195 345.150 ;
        RECT 246.385 344.980 246.555 345.150 ;
        RECT 252.255 344.980 252.425 345.150 ;
        RECT 252.615 344.980 252.785 345.150 ;
        RECT 255.725 344.980 255.895 345.150 ;
        RECT 256.085 344.980 256.255 345.150 ;
        RECT 259.195 344.980 259.365 345.150 ;
        RECT 259.555 344.980 259.725 345.150 ;
        RECT 262.665 344.980 262.835 345.150 ;
        RECT 263.025 344.980 263.195 345.150 ;
        RECT 266.135 344.980 266.305 345.150 ;
        RECT 266.495 344.980 266.665 345.150 ;
        RECT 272.365 344.980 272.535 345.150 ;
        RECT 272.725 344.980 272.895 345.150 ;
        RECT 275.835 344.980 276.005 345.150 ;
        RECT 276.195 344.980 276.365 345.150 ;
        RECT 279.305 344.980 279.475 345.150 ;
        RECT 279.665 344.980 279.835 345.150 ;
        RECT 282.775 344.980 282.945 345.150 ;
        RECT 283.135 344.980 283.305 345.150 ;
        RECT 286.245 344.980 286.415 345.150 ;
        RECT 286.605 344.980 286.775 345.150 ;
        RECT 355.435 345.815 355.605 345.985 ;
        RECT 355.435 345.455 355.605 345.625 ;
        RECT 355.435 345.095 355.605 345.265 ;
        RECT 212.175 341.690 212.345 341.860 ;
        RECT 212.535 341.690 212.705 341.860 ;
        RECT 215.645 341.690 215.815 341.860 ;
        RECT 216.005 341.690 216.175 341.860 ;
        RECT 219.115 341.690 219.285 341.860 ;
        RECT 219.475 341.690 219.645 341.860 ;
        RECT 222.585 341.690 222.755 341.860 ;
        RECT 222.945 341.690 223.115 341.860 ;
        RECT 226.055 341.690 226.225 341.860 ;
        RECT 226.415 341.690 226.585 341.860 ;
        RECT 232.145 341.690 232.315 341.860 ;
        RECT 232.505 341.690 232.675 341.860 ;
        RECT 235.615 341.690 235.785 341.860 ;
        RECT 235.975 341.690 236.145 341.860 ;
        RECT 239.085 341.690 239.255 341.860 ;
        RECT 239.445 341.690 239.615 341.860 ;
        RECT 242.555 341.690 242.725 341.860 ;
        RECT 242.915 341.690 243.085 341.860 ;
        RECT 246.025 341.690 246.195 341.860 ;
        RECT 246.385 341.690 246.555 341.860 ;
        RECT 212.175 338.400 212.345 338.570 ;
        RECT 212.535 338.400 212.705 338.570 ;
        RECT 215.645 338.400 215.815 338.570 ;
        RECT 216.005 338.400 216.175 338.570 ;
        RECT 219.115 338.400 219.285 338.570 ;
        RECT 219.475 338.400 219.645 338.570 ;
        RECT 222.585 338.400 222.755 338.570 ;
        RECT 222.945 338.400 223.115 338.570 ;
        RECT 226.055 338.400 226.225 338.570 ;
        RECT 226.415 338.400 226.585 338.570 ;
        RECT 212.175 335.110 212.345 335.280 ;
        RECT 212.535 335.110 212.705 335.280 ;
        RECT 215.645 335.110 215.815 335.280 ;
        RECT 216.005 335.110 216.175 335.280 ;
        RECT 219.115 335.110 219.285 335.280 ;
        RECT 219.475 335.110 219.645 335.280 ;
        RECT 222.585 335.110 222.755 335.280 ;
        RECT 222.945 335.110 223.115 335.280 ;
        RECT 226.055 335.110 226.225 335.280 ;
        RECT 226.415 335.110 226.585 335.280 ;
        RECT 5.435 329.260 5.605 329.430 ;
        RECT 5.795 329.260 5.965 329.430 ;
        RECT 6.155 329.260 6.325 329.430 ;
        RECT 6.515 329.260 6.685 329.430 ;
        RECT 6.875 329.260 7.045 329.430 ;
        RECT 7.235 329.260 7.405 329.430 ;
        RECT 7.595 329.260 7.765 329.430 ;
        RECT 7.955 329.260 8.125 329.430 ;
        RECT 8.315 329.260 8.485 329.430 ;
        RECT 8.675 329.260 8.845 329.430 ;
        RECT 9.035 329.260 9.205 329.430 ;
        RECT 9.395 329.260 9.565 329.430 ;
        RECT 9.755 329.260 9.925 329.430 ;
        RECT 10.115 329.260 10.285 329.430 ;
        RECT 10.475 329.260 10.645 329.430 ;
        RECT 10.835 329.260 11.005 329.430 ;
        RECT 11.195 329.260 11.365 329.430 ;
        RECT 11.555 329.260 11.725 329.430 ;
        RECT 11.915 329.260 12.085 329.430 ;
        RECT 12.275 329.260 12.445 329.430 ;
        RECT 18.775 329.240 18.945 329.410 ;
        RECT 19.135 329.240 19.305 329.410 ;
        RECT 19.495 329.240 19.665 329.410 ;
        RECT 19.855 329.240 20.025 329.410 ;
        RECT 20.215 329.240 20.385 329.410 ;
        RECT 20.575 329.240 20.745 329.410 ;
        RECT 20.935 329.240 21.105 329.410 ;
        RECT 21.295 329.240 21.465 329.410 ;
        RECT 21.655 329.240 21.825 329.410 ;
        RECT 22.015 329.240 22.185 329.410 ;
        RECT 22.375 329.240 22.545 329.410 ;
        RECT 22.735 329.240 22.905 329.410 ;
        RECT 23.095 329.240 23.265 329.410 ;
        RECT 23.455 329.240 23.625 329.410 ;
        RECT 23.815 329.240 23.985 329.410 ;
        RECT 24.175 329.240 24.345 329.410 ;
        RECT 24.535 329.240 24.705 329.410 ;
        RECT 24.895 329.240 25.065 329.410 ;
        RECT 25.255 329.240 25.425 329.410 ;
        RECT 25.615 329.240 25.785 329.410 ;
        RECT 32.145 329.270 32.315 329.440 ;
        RECT 32.505 329.270 32.675 329.440 ;
        RECT 32.865 329.270 33.035 329.440 ;
        RECT 33.225 329.270 33.395 329.440 ;
        RECT 33.585 329.270 33.755 329.440 ;
        RECT 33.945 329.270 34.115 329.440 ;
        RECT 34.305 329.270 34.475 329.440 ;
        RECT 34.665 329.270 34.835 329.440 ;
        RECT 35.025 329.270 35.195 329.440 ;
        RECT 35.385 329.270 35.555 329.440 ;
        RECT 35.745 329.270 35.915 329.440 ;
        RECT 36.105 329.270 36.275 329.440 ;
        RECT 36.465 329.270 36.635 329.440 ;
        RECT 36.825 329.270 36.995 329.440 ;
        RECT 37.185 329.270 37.355 329.440 ;
        RECT 37.545 329.270 37.715 329.440 ;
        RECT 37.905 329.270 38.075 329.440 ;
        RECT 38.265 329.270 38.435 329.440 ;
        RECT 38.625 329.270 38.795 329.440 ;
        RECT 38.985 329.270 39.155 329.440 ;
        RECT 45.375 329.270 45.545 329.440 ;
        RECT 45.735 329.270 45.905 329.440 ;
        RECT 46.095 329.270 46.265 329.440 ;
        RECT 46.455 329.270 46.625 329.440 ;
        RECT 46.815 329.270 46.985 329.440 ;
        RECT 47.175 329.270 47.345 329.440 ;
        RECT 47.535 329.270 47.705 329.440 ;
        RECT 47.895 329.270 48.065 329.440 ;
        RECT 48.255 329.270 48.425 329.440 ;
        RECT 48.615 329.270 48.785 329.440 ;
        RECT 48.975 329.270 49.145 329.440 ;
        RECT 49.335 329.270 49.505 329.440 ;
        RECT 49.695 329.270 49.865 329.440 ;
        RECT 50.055 329.270 50.225 329.440 ;
        RECT 50.415 329.270 50.585 329.440 ;
        RECT 50.775 329.270 50.945 329.440 ;
        RECT 51.135 329.270 51.305 329.440 ;
        RECT 51.495 329.270 51.665 329.440 ;
        RECT 51.855 329.270 52.025 329.440 ;
        RECT 52.215 329.270 52.385 329.440 ;
        RECT 58.645 329.240 58.815 329.410 ;
        RECT 59.005 329.240 59.175 329.410 ;
        RECT 59.365 329.240 59.535 329.410 ;
        RECT 59.725 329.240 59.895 329.410 ;
        RECT 60.085 329.240 60.255 329.410 ;
        RECT 60.445 329.240 60.615 329.410 ;
        RECT 60.805 329.240 60.975 329.410 ;
        RECT 61.165 329.240 61.335 329.410 ;
        RECT 61.525 329.240 61.695 329.410 ;
        RECT 61.885 329.240 62.055 329.410 ;
        RECT 62.245 329.240 62.415 329.410 ;
        RECT 62.605 329.240 62.775 329.410 ;
        RECT 62.965 329.240 63.135 329.410 ;
        RECT 63.325 329.240 63.495 329.410 ;
        RECT 63.685 329.240 63.855 329.410 ;
        RECT 64.045 329.240 64.215 329.410 ;
        RECT 64.405 329.240 64.575 329.410 ;
        RECT 64.765 329.240 64.935 329.410 ;
        RECT 65.125 329.240 65.295 329.410 ;
        RECT 65.485 329.240 65.655 329.410 ;
        RECT 71.915 329.270 72.085 329.440 ;
        RECT 72.275 329.270 72.445 329.440 ;
        RECT 72.635 329.270 72.805 329.440 ;
        RECT 72.995 329.270 73.165 329.440 ;
        RECT 73.355 329.270 73.525 329.440 ;
        RECT 73.715 329.270 73.885 329.440 ;
        RECT 74.075 329.270 74.245 329.440 ;
        RECT 74.435 329.270 74.605 329.440 ;
        RECT 74.795 329.270 74.965 329.440 ;
        RECT 75.155 329.270 75.325 329.440 ;
        RECT 75.515 329.270 75.685 329.440 ;
        RECT 75.875 329.270 76.045 329.440 ;
        RECT 76.235 329.270 76.405 329.440 ;
        RECT 76.595 329.270 76.765 329.440 ;
        RECT 76.955 329.270 77.125 329.440 ;
        RECT 77.315 329.270 77.485 329.440 ;
        RECT 77.675 329.270 77.845 329.440 ;
        RECT 78.035 329.270 78.205 329.440 ;
        RECT 78.395 329.270 78.565 329.440 ;
        RECT 78.755 329.270 78.925 329.440 ;
        RECT 85.045 329.290 85.215 329.460 ;
        RECT 85.405 329.290 85.575 329.460 ;
        RECT 85.765 329.290 85.935 329.460 ;
        RECT 86.125 329.290 86.295 329.460 ;
        RECT 86.485 329.290 86.655 329.460 ;
        RECT 86.845 329.290 87.015 329.460 ;
        RECT 87.205 329.290 87.375 329.460 ;
        RECT 87.565 329.290 87.735 329.460 ;
        RECT 87.925 329.290 88.095 329.460 ;
        RECT 88.285 329.290 88.455 329.460 ;
        RECT 88.645 329.290 88.815 329.460 ;
        RECT 89.005 329.290 89.175 329.460 ;
        RECT 89.365 329.290 89.535 329.460 ;
        RECT 89.725 329.290 89.895 329.460 ;
        RECT 90.085 329.290 90.255 329.460 ;
        RECT 90.445 329.290 90.615 329.460 ;
        RECT 90.805 329.290 90.975 329.460 ;
        RECT 91.165 329.290 91.335 329.460 ;
        RECT 91.525 329.290 91.695 329.460 ;
        RECT 91.885 329.290 92.055 329.460 ;
        RECT 97.960 329.085 102.450 329.615 ;
        RECT 252.255 341.690 252.425 341.860 ;
        RECT 252.615 341.690 252.785 341.860 ;
        RECT 255.725 341.690 255.895 341.860 ;
        RECT 256.085 341.690 256.255 341.860 ;
        RECT 259.195 341.690 259.365 341.860 ;
        RECT 259.555 341.690 259.725 341.860 ;
        RECT 262.665 341.690 262.835 341.860 ;
        RECT 263.025 341.690 263.195 341.860 ;
        RECT 266.135 341.690 266.305 341.860 ;
        RECT 266.495 341.690 266.665 341.860 ;
        RECT 232.145 338.400 232.315 338.570 ;
        RECT 232.505 338.400 232.675 338.570 ;
        RECT 235.615 338.400 235.785 338.570 ;
        RECT 235.975 338.400 236.145 338.570 ;
        RECT 239.085 338.400 239.255 338.570 ;
        RECT 239.445 338.400 239.615 338.570 ;
        RECT 242.555 338.400 242.725 338.570 ;
        RECT 242.915 338.400 243.085 338.570 ;
        RECT 246.025 338.400 246.195 338.570 ;
        RECT 246.385 338.400 246.555 338.570 ;
        RECT 232.145 335.110 232.315 335.280 ;
        RECT 232.505 335.110 232.675 335.280 ;
        RECT 235.615 335.110 235.785 335.280 ;
        RECT 235.975 335.110 236.145 335.280 ;
        RECT 239.085 335.110 239.255 335.280 ;
        RECT 239.445 335.110 239.615 335.280 ;
        RECT 242.555 335.110 242.725 335.280 ;
        RECT 242.915 335.110 243.085 335.280 ;
        RECT 246.025 335.110 246.195 335.280 ;
        RECT 246.385 335.110 246.555 335.280 ;
        RECT 212.175 331.820 212.345 331.990 ;
        RECT 212.535 331.820 212.705 331.990 ;
        RECT 215.645 331.820 215.815 331.990 ;
        RECT 216.005 331.820 216.175 331.990 ;
        RECT 219.115 331.820 219.285 331.990 ;
        RECT 219.475 331.820 219.645 331.990 ;
        RECT 222.585 331.820 222.755 331.990 ;
        RECT 222.945 331.820 223.115 331.990 ;
        RECT 226.055 331.820 226.225 331.990 ;
        RECT 226.415 331.820 226.585 331.990 ;
        RECT 272.365 341.690 272.535 341.860 ;
        RECT 272.725 341.690 272.895 341.860 ;
        RECT 275.835 341.690 276.005 341.860 ;
        RECT 276.195 341.690 276.365 341.860 ;
        RECT 279.305 341.690 279.475 341.860 ;
        RECT 279.665 341.690 279.835 341.860 ;
        RECT 282.775 341.690 282.945 341.860 ;
        RECT 283.135 341.690 283.305 341.860 ;
        RECT 286.245 341.690 286.415 341.860 ;
        RECT 286.605 341.690 286.775 341.860 ;
        RECT 252.255 338.400 252.425 338.570 ;
        RECT 252.615 338.400 252.785 338.570 ;
        RECT 255.725 338.400 255.895 338.570 ;
        RECT 256.085 338.400 256.255 338.570 ;
        RECT 259.195 338.400 259.365 338.570 ;
        RECT 259.555 338.400 259.725 338.570 ;
        RECT 262.665 338.400 262.835 338.570 ;
        RECT 263.025 338.400 263.195 338.570 ;
        RECT 266.135 338.400 266.305 338.570 ;
        RECT 266.495 338.400 266.665 338.570 ;
        RECT 252.255 335.110 252.425 335.280 ;
        RECT 252.615 335.110 252.785 335.280 ;
        RECT 255.725 335.110 255.895 335.280 ;
        RECT 256.085 335.110 256.255 335.280 ;
        RECT 259.195 335.110 259.365 335.280 ;
        RECT 259.555 335.110 259.725 335.280 ;
        RECT 262.665 335.110 262.835 335.280 ;
        RECT 263.025 335.110 263.195 335.280 ;
        RECT 266.135 335.110 266.305 335.280 ;
        RECT 266.495 335.110 266.665 335.280 ;
        RECT 232.145 331.820 232.315 331.990 ;
        RECT 232.505 331.820 232.675 331.990 ;
        RECT 235.615 331.820 235.785 331.990 ;
        RECT 235.975 331.820 236.145 331.990 ;
        RECT 239.085 331.820 239.255 331.990 ;
        RECT 239.445 331.820 239.615 331.990 ;
        RECT 242.555 331.820 242.725 331.990 ;
        RECT 242.915 331.820 243.085 331.990 ;
        RECT 246.025 331.820 246.195 331.990 ;
        RECT 246.385 331.820 246.555 331.990 ;
        RECT 355.435 344.735 355.605 344.905 ;
        RECT 355.435 344.375 355.605 344.545 ;
        RECT 355.435 344.015 355.605 344.185 ;
        RECT 355.435 343.655 355.605 343.825 ;
        RECT 355.435 343.295 355.605 343.465 ;
        RECT 355.435 342.935 355.605 343.105 ;
        RECT 355.435 342.575 355.605 342.745 ;
        RECT 355.435 342.215 355.605 342.385 ;
        RECT 355.435 341.855 355.605 342.025 ;
        RECT 355.435 341.495 355.605 341.665 ;
        RECT 355.435 341.135 355.605 341.305 ;
        RECT 355.435 340.775 355.605 340.945 ;
        RECT 355.435 340.415 355.605 340.585 ;
        RECT 355.435 340.055 355.605 340.225 ;
        RECT 355.435 339.695 355.605 339.865 ;
        RECT 355.435 339.335 355.605 339.505 ;
        RECT 355.435 338.975 355.605 339.145 ;
        RECT 272.365 338.400 272.535 338.570 ;
        RECT 272.725 338.400 272.895 338.570 ;
        RECT 275.835 338.400 276.005 338.570 ;
        RECT 276.195 338.400 276.365 338.570 ;
        RECT 279.305 338.400 279.475 338.570 ;
        RECT 279.665 338.400 279.835 338.570 ;
        RECT 282.775 338.400 282.945 338.570 ;
        RECT 283.135 338.400 283.305 338.570 ;
        RECT 286.245 338.400 286.415 338.570 ;
        RECT 286.605 338.400 286.775 338.570 ;
        RECT 355.435 338.615 355.605 338.785 ;
        RECT 272.365 335.110 272.535 335.280 ;
        RECT 272.725 335.110 272.895 335.280 ;
        RECT 275.835 335.110 276.005 335.280 ;
        RECT 276.195 335.110 276.365 335.280 ;
        RECT 279.305 335.110 279.475 335.280 ;
        RECT 279.665 335.110 279.835 335.280 ;
        RECT 282.775 335.110 282.945 335.280 ;
        RECT 283.135 335.110 283.305 335.280 ;
        RECT 286.245 335.110 286.415 335.280 ;
        RECT 286.605 335.110 286.775 335.280 ;
        RECT 252.255 331.820 252.425 331.990 ;
        RECT 252.615 331.820 252.785 331.990 ;
        RECT 255.725 331.820 255.895 331.990 ;
        RECT 256.085 331.820 256.255 331.990 ;
        RECT 259.195 331.820 259.365 331.990 ;
        RECT 259.555 331.820 259.725 331.990 ;
        RECT 262.665 331.820 262.835 331.990 ;
        RECT 263.025 331.820 263.195 331.990 ;
        RECT 266.135 331.820 266.305 331.990 ;
        RECT 266.495 331.820 266.665 331.990 ;
        RECT 355.435 338.255 355.605 338.425 ;
        RECT 355.435 337.895 355.605 338.065 ;
        RECT 355.435 337.535 355.605 337.705 ;
        RECT 355.435 337.175 355.605 337.345 ;
        RECT 355.435 336.815 355.605 336.985 ;
        RECT 355.435 336.455 355.605 336.625 ;
        RECT 355.435 336.095 355.605 336.265 ;
        RECT 355.435 335.735 355.605 335.905 ;
        RECT 355.435 335.375 355.605 335.545 ;
        RECT 355.435 335.015 355.605 335.185 ;
        RECT 355.435 334.655 355.605 334.825 ;
        RECT 355.435 334.295 355.605 334.465 ;
        RECT 355.435 333.935 355.605 334.105 ;
        RECT 355.435 333.575 355.605 333.745 ;
        RECT 355.435 333.215 355.605 333.385 ;
        RECT 356.530 346.415 356.700 346.585 ;
        RECT 356.530 346.055 356.700 346.225 ;
        RECT 356.530 342.945 356.700 343.115 ;
        RECT 356.530 342.585 356.700 342.755 ;
        RECT 356.530 339.475 356.700 339.645 ;
        RECT 356.530 339.115 356.700 339.285 ;
        RECT 356.530 336.005 356.700 336.175 ;
        RECT 356.530 335.645 356.700 335.815 ;
        RECT 382.450 350.955 382.620 351.125 ;
        RECT 394.025 364.665 394.195 364.835 ;
        RECT 394.025 364.305 394.195 364.475 ;
        RECT 395.120 365.265 395.290 365.435 ;
        RECT 395.120 364.905 395.290 365.075 ;
        RECT 394.025 363.945 394.195 364.115 ;
        RECT 394.025 363.585 394.195 363.755 ;
        RECT 394.025 363.225 394.195 363.395 ;
        RECT 394.025 362.865 394.195 363.035 ;
        RECT 394.025 362.505 394.195 362.675 ;
        RECT 394.025 362.145 394.195 362.315 ;
        RECT 394.025 361.785 394.195 361.955 ;
        RECT 394.025 361.425 394.195 361.595 ;
        RECT 394.025 361.065 394.195 361.235 ;
        RECT 394.025 360.705 394.195 360.875 ;
        RECT 394.025 360.345 394.195 360.515 ;
        RECT 394.025 359.985 394.195 360.155 ;
        RECT 394.025 359.625 394.195 359.795 ;
        RECT 394.025 359.265 394.195 359.435 ;
        RECT 394.025 358.905 394.195 359.075 ;
        RECT 394.025 358.545 394.195 358.715 ;
        RECT 394.025 358.185 394.195 358.355 ;
        RECT 394.025 357.825 394.195 357.995 ;
        RECT 394.025 357.465 394.195 357.635 ;
        RECT 394.025 357.105 394.195 357.275 ;
        RECT 394.025 356.745 394.195 356.915 ;
        RECT 394.025 356.385 394.195 356.555 ;
        RECT 394.025 356.025 394.195 356.195 ;
        RECT 394.025 355.665 394.195 355.835 ;
        RECT 394.025 355.305 394.195 355.475 ;
        RECT 394.025 354.945 394.195 355.115 ;
        RECT 394.025 354.585 394.195 354.755 ;
        RECT 394.025 354.225 394.195 354.395 ;
        RECT 394.025 353.865 394.195 354.035 ;
        RECT 394.025 353.505 394.195 353.675 ;
        RECT 394.025 353.145 394.195 353.315 ;
        RECT 394.025 352.785 394.195 352.955 ;
        RECT 394.025 352.425 394.195 352.595 ;
        RECT 394.025 352.065 394.195 352.235 ;
        RECT 395.120 361.795 395.290 361.965 ;
        RECT 395.120 361.435 395.290 361.605 ;
        RECT 395.120 358.325 395.290 358.495 ;
        RECT 395.120 357.965 395.290 358.135 ;
        RECT 395.120 354.855 395.290 355.025 ;
        RECT 395.120 354.495 395.290 354.665 ;
        RECT 395.120 351.385 395.290 351.555 ;
        RECT 398.410 365.265 398.580 365.435 ;
        RECT 398.410 364.905 398.580 365.075 ;
        RECT 398.410 361.795 398.580 361.965 ;
        RECT 398.410 361.435 398.580 361.605 ;
        RECT 398.410 358.325 398.580 358.495 ;
        RECT 398.410 357.965 398.580 358.135 ;
        RECT 398.410 354.855 398.580 355.025 ;
        RECT 398.410 354.495 398.580 354.665 ;
        RECT 398.410 351.385 398.580 351.555 ;
        RECT 389.030 350.955 389.200 351.125 ;
        RECT 395.120 351.025 395.290 351.195 ;
        RECT 359.820 346.415 359.990 346.585 ;
        RECT 359.820 346.055 359.990 346.225 ;
        RECT 359.820 342.945 359.990 343.115 ;
        RECT 359.820 342.585 359.990 342.755 ;
        RECT 359.820 339.475 359.990 339.645 ;
        RECT 359.820 339.115 359.990 339.285 ;
        RECT 359.820 336.005 359.990 336.175 ;
        RECT 359.820 335.645 359.990 335.815 ;
        RECT 356.530 332.535 356.700 332.705 ;
        RECT 356.530 332.175 356.700 332.345 ;
        RECT 272.365 331.820 272.535 331.990 ;
        RECT 272.725 331.820 272.895 331.990 ;
        RECT 275.835 331.820 276.005 331.990 ;
        RECT 276.195 331.820 276.365 331.990 ;
        RECT 279.305 331.820 279.475 331.990 ;
        RECT 279.665 331.820 279.835 331.990 ;
        RECT 282.775 331.820 282.945 331.990 ;
        RECT 283.135 331.820 283.305 331.990 ;
        RECT 286.245 331.820 286.415 331.990 ;
        RECT 286.605 331.820 286.775 331.990 ;
        RECT 212.175 328.530 212.345 328.700 ;
        RECT 212.535 328.530 212.705 328.700 ;
        RECT 215.645 328.530 215.815 328.700 ;
        RECT 216.005 328.530 216.175 328.700 ;
        RECT 219.115 328.530 219.285 328.700 ;
        RECT 219.475 328.530 219.645 328.700 ;
        RECT 222.585 328.530 222.755 328.700 ;
        RECT 222.945 328.530 223.115 328.700 ;
        RECT 226.055 328.530 226.225 328.700 ;
        RECT 226.415 328.530 226.585 328.700 ;
        RECT 232.145 328.530 232.315 328.700 ;
        RECT 232.505 328.530 232.675 328.700 ;
        RECT 235.615 328.530 235.785 328.700 ;
        RECT 235.975 328.530 236.145 328.700 ;
        RECT 239.085 328.530 239.255 328.700 ;
        RECT 239.445 328.530 239.615 328.700 ;
        RECT 242.555 328.530 242.725 328.700 ;
        RECT 242.915 328.530 243.085 328.700 ;
        RECT 246.025 328.530 246.195 328.700 ;
        RECT 246.385 328.530 246.555 328.700 ;
        RECT 252.255 328.530 252.425 328.700 ;
        RECT 252.615 328.530 252.785 328.700 ;
        RECT 255.725 328.530 255.895 328.700 ;
        RECT 256.085 328.530 256.255 328.700 ;
        RECT 259.195 328.530 259.365 328.700 ;
        RECT 259.555 328.530 259.725 328.700 ;
        RECT 262.665 328.530 262.835 328.700 ;
        RECT 263.025 328.530 263.195 328.700 ;
        RECT 266.135 328.530 266.305 328.700 ;
        RECT 266.495 328.530 266.665 328.700 ;
        RECT 272.365 328.530 272.535 328.700 ;
        RECT 272.725 328.530 272.895 328.700 ;
        RECT 275.835 328.530 276.005 328.700 ;
        RECT 276.195 328.530 276.365 328.700 ;
        RECT 279.305 328.530 279.475 328.700 ;
        RECT 279.665 328.530 279.835 328.700 ;
        RECT 282.775 328.530 282.945 328.700 ;
        RECT 283.135 328.530 283.305 328.700 ;
        RECT 286.245 328.530 286.415 328.700 ;
        RECT 286.605 328.530 286.775 328.700 ;
        RECT 359.820 332.535 359.990 332.705 ;
        RECT 363.110 346.415 363.280 346.585 ;
        RECT 363.110 346.055 363.280 346.225 ;
        RECT 363.110 342.945 363.280 343.115 ;
        RECT 363.110 342.585 363.280 342.755 ;
        RECT 363.110 339.475 363.280 339.645 ;
        RECT 363.110 339.115 363.280 339.285 ;
        RECT 363.110 336.005 363.280 336.175 ;
        RECT 363.110 335.645 363.280 335.815 ;
        RECT 363.110 332.535 363.280 332.705 ;
        RECT 366.400 346.415 366.570 346.585 ;
        RECT 369.690 346.415 369.860 346.585 ;
        RECT 366.400 346.055 366.570 346.225 ;
        RECT 366.400 342.945 366.570 343.115 ;
        RECT 366.400 342.585 366.570 342.755 ;
        RECT 366.400 339.475 366.570 339.645 ;
        RECT 366.400 339.115 366.570 339.285 ;
        RECT 366.400 336.005 366.570 336.175 ;
        RECT 366.400 335.645 366.570 335.815 ;
        RECT 366.400 332.535 366.570 332.705 ;
        RECT 369.690 346.055 369.860 346.225 ;
        RECT 369.690 342.945 369.860 343.115 ;
        RECT 369.690 342.585 369.860 342.755 ;
        RECT 369.690 339.475 369.860 339.645 ;
        RECT 369.690 339.115 369.860 339.285 ;
        RECT 369.690 336.005 369.860 336.175 ;
        RECT 369.690 335.645 369.860 335.815 ;
        RECT 359.820 332.175 359.990 332.345 ;
        RECT 363.110 332.175 363.280 332.345 ;
        RECT 366.400 332.175 366.570 332.345 ;
        RECT 369.690 332.535 369.860 332.705 ;
        RECT 374.755 345.715 374.925 345.885 ;
        RECT 374.755 345.355 374.925 345.525 ;
        RECT 374.755 344.995 374.925 345.165 ;
        RECT 374.755 344.635 374.925 344.805 ;
        RECT 374.755 344.275 374.925 344.445 ;
        RECT 374.755 343.915 374.925 344.085 ;
        RECT 374.755 343.555 374.925 343.725 ;
        RECT 374.755 343.195 374.925 343.365 ;
        RECT 374.755 342.835 374.925 343.005 ;
        RECT 374.755 342.475 374.925 342.645 ;
        RECT 374.755 342.115 374.925 342.285 ;
        RECT 374.755 341.755 374.925 341.925 ;
        RECT 374.755 341.395 374.925 341.565 ;
        RECT 374.755 341.035 374.925 341.205 ;
        RECT 374.755 340.675 374.925 340.845 ;
        RECT 374.755 340.315 374.925 340.485 ;
        RECT 374.755 339.955 374.925 340.125 ;
        RECT 374.755 339.595 374.925 339.765 ;
        RECT 374.755 339.235 374.925 339.405 ;
        RECT 374.755 338.875 374.925 339.045 ;
        RECT 374.755 338.515 374.925 338.685 ;
        RECT 374.755 338.155 374.925 338.325 ;
        RECT 374.755 337.795 374.925 337.965 ;
        RECT 374.755 337.435 374.925 337.605 ;
        RECT 374.755 337.075 374.925 337.245 ;
        RECT 374.755 336.715 374.925 336.885 ;
        RECT 374.755 336.355 374.925 336.525 ;
        RECT 374.755 335.995 374.925 336.165 ;
        RECT 374.755 335.635 374.925 335.805 ;
        RECT 374.755 335.275 374.925 335.445 ;
        RECT 374.755 334.915 374.925 335.085 ;
        RECT 374.755 334.555 374.925 334.725 ;
        RECT 374.755 334.195 374.925 334.365 ;
        RECT 374.755 333.835 374.925 334.005 ;
        RECT 374.755 333.475 374.925 333.645 ;
        RECT 374.755 333.115 374.925 333.285 ;
        RECT 375.850 346.315 376.020 346.485 ;
        RECT 375.850 345.955 376.020 346.125 ;
        RECT 375.850 342.845 376.020 343.015 ;
        RECT 375.850 342.485 376.020 342.655 ;
        RECT 375.850 339.375 376.020 339.545 ;
        RECT 375.850 339.015 376.020 339.185 ;
        RECT 375.850 335.905 376.020 336.075 ;
        RECT 375.850 335.545 376.020 335.715 ;
        RECT 382.430 346.315 382.600 346.485 ;
        RECT 401.700 365.265 401.870 365.435 ;
        RECT 401.700 364.905 401.870 365.075 ;
        RECT 401.700 361.795 401.870 361.965 ;
        RECT 401.700 361.435 401.870 361.605 ;
        RECT 401.700 358.325 401.870 358.495 ;
        RECT 401.700 357.965 401.870 358.135 ;
        RECT 401.700 354.855 401.870 355.025 ;
        RECT 401.700 354.495 401.870 354.665 ;
        RECT 401.700 351.385 401.870 351.555 ;
        RECT 404.990 365.265 405.160 365.435 ;
        RECT 408.280 365.265 408.450 365.435 ;
        RECT 404.990 364.905 405.160 365.075 ;
        RECT 404.990 361.795 405.160 361.965 ;
        RECT 404.990 361.435 405.160 361.605 ;
        RECT 404.990 358.325 405.160 358.495 ;
        RECT 404.990 357.965 405.160 358.135 ;
        RECT 404.990 354.855 405.160 355.025 ;
        RECT 404.990 354.495 405.160 354.665 ;
        RECT 404.990 351.385 405.160 351.555 ;
        RECT 408.280 364.905 408.450 365.075 ;
        RECT 408.280 361.795 408.450 361.965 ;
        RECT 408.280 361.435 408.450 361.605 ;
        RECT 408.280 358.325 408.450 358.495 ;
        RECT 408.280 357.965 408.450 358.135 ;
        RECT 408.280 354.855 408.450 355.025 ;
        RECT 654.125 354.845 654.295 355.015 ;
        RECT 654.605 354.845 654.775 355.015 ;
        RECT 655.085 354.845 655.255 355.015 ;
        RECT 408.280 354.495 408.450 354.665 ;
        RECT 654.760 354.365 654.930 354.535 ;
        RECT 655.120 354.365 655.290 354.535 ;
        RECT 657.705 354.835 657.875 355.005 ;
        RECT 658.185 354.835 658.355 355.005 ;
        RECT 658.665 354.835 658.835 355.005 ;
        RECT 659.145 354.835 659.315 355.005 ;
        RECT 659.625 354.835 659.795 355.005 ;
        RECT 660.105 354.835 660.275 355.005 ;
        RECT 660.585 354.835 660.755 355.005 ;
        RECT 661.065 354.835 661.235 355.005 ;
        RECT 661.545 354.835 661.715 355.005 ;
        RECT 662.025 354.835 662.195 355.005 ;
        RECT 662.505 354.835 662.675 355.005 ;
        RECT 662.985 354.835 663.155 355.005 ;
        RECT 663.465 354.835 663.635 355.005 ;
        RECT 663.945 354.835 664.115 355.005 ;
        RECT 664.425 354.835 664.595 355.005 ;
        RECT 664.905 354.835 665.075 355.005 ;
        RECT 665.385 354.835 665.555 355.005 ;
        RECT 665.865 354.835 666.035 355.005 ;
        RECT 666.345 354.835 666.515 355.005 ;
        RECT 666.825 354.835 666.995 355.005 ;
        RECT 667.305 354.835 667.475 355.005 ;
        RECT 667.785 354.835 667.955 355.005 ;
        RECT 668.265 354.835 668.435 355.005 ;
        RECT 668.745 354.835 668.915 355.005 ;
        RECT 669.225 354.835 669.395 355.005 ;
        RECT 669.705 354.835 669.875 355.005 ;
        RECT 670.185 354.835 670.355 355.005 ;
        RECT 670.665 354.835 670.835 355.005 ;
        RECT 671.145 354.835 671.315 355.005 ;
        RECT 671.625 354.835 671.795 355.005 ;
        RECT 672.105 354.835 672.275 355.005 ;
        RECT 672.585 354.835 672.755 355.005 ;
        RECT 658.220 354.355 658.390 354.525 ;
        RECT 658.580 354.355 658.750 354.525 ;
        RECT 658.940 354.355 659.110 354.525 ;
        RECT 659.750 354.355 659.920 354.525 ;
        RECT 660.110 354.355 660.280 354.525 ;
        RECT 660.470 354.355 660.640 354.525 ;
        RECT 661.505 354.355 661.675 354.525 ;
        RECT 661.865 354.355 662.035 354.525 ;
        RECT 662.225 354.355 662.395 354.525 ;
        RECT 664.200 354.355 664.370 354.525 ;
        RECT 664.560 354.355 664.730 354.525 ;
        RECT 664.920 354.355 665.090 354.525 ;
        RECT 666.540 354.355 666.710 354.525 ;
        RECT 666.900 354.355 667.070 354.525 ;
        RECT 667.260 354.355 667.430 354.525 ;
        RECT 669.690 354.355 669.860 354.525 ;
        RECT 671.720 354.355 671.890 354.525 ;
        RECT 672.080 354.355 672.250 354.525 ;
        RECT 675.755 354.795 675.925 354.965 ;
        RECT 676.235 354.795 676.405 354.965 ;
        RECT 676.715 354.795 676.885 354.965 ;
        RECT 677.195 354.795 677.365 354.965 ;
        RECT 677.675 354.795 677.845 354.965 ;
        RECT 678.155 354.795 678.325 354.965 ;
        RECT 678.635 354.795 678.805 354.965 ;
        RECT 679.115 354.795 679.285 354.965 ;
        RECT 679.595 354.795 679.765 354.965 ;
        RECT 680.075 354.795 680.245 354.965 ;
        RECT 680.555 354.795 680.725 354.965 ;
        RECT 681.035 354.795 681.205 354.965 ;
        RECT 681.515 354.795 681.685 354.965 ;
        RECT 681.995 354.795 682.165 354.965 ;
        RECT 682.475 354.795 682.645 354.965 ;
        RECT 682.955 354.795 683.125 354.965 ;
        RECT 683.435 354.795 683.605 354.965 ;
        RECT 683.915 354.795 684.085 354.965 ;
        RECT 684.395 354.795 684.565 354.965 ;
        RECT 684.875 354.795 685.045 354.965 ;
        RECT 685.355 354.795 685.525 354.965 ;
        RECT 685.835 354.795 686.005 354.965 ;
        RECT 686.315 354.795 686.485 354.965 ;
        RECT 686.795 354.795 686.965 354.965 ;
        RECT 687.275 354.795 687.445 354.965 ;
        RECT 687.755 354.795 687.925 354.965 ;
        RECT 688.235 354.795 688.405 354.965 ;
        RECT 688.715 354.795 688.885 354.965 ;
        RECT 689.195 354.795 689.365 354.965 ;
        RECT 689.675 354.795 689.845 354.965 ;
        RECT 690.155 354.795 690.325 354.965 ;
        RECT 690.635 354.795 690.805 354.965 ;
        RECT 676.270 354.315 676.440 354.485 ;
        RECT 676.630 354.315 676.800 354.485 ;
        RECT 676.990 354.315 677.160 354.485 ;
        RECT 677.800 354.315 677.970 354.485 ;
        RECT 678.160 354.315 678.330 354.485 ;
        RECT 678.520 354.315 678.690 354.485 ;
        RECT 679.555 354.315 679.725 354.485 ;
        RECT 679.915 354.315 680.085 354.485 ;
        RECT 680.275 354.315 680.445 354.485 ;
        RECT 682.250 354.315 682.420 354.485 ;
        RECT 682.610 354.315 682.780 354.485 ;
        RECT 682.970 354.315 683.140 354.485 ;
        RECT 684.590 354.315 684.760 354.485 ;
        RECT 684.950 354.315 685.120 354.485 ;
        RECT 685.310 354.315 685.480 354.485 ;
        RECT 687.740 354.315 687.910 354.485 ;
        RECT 689.770 354.315 689.940 354.485 ;
        RECT 690.130 354.315 690.300 354.485 ;
        RECT 693.345 354.815 693.515 354.985 ;
        RECT 693.825 354.815 693.995 354.985 ;
        RECT 694.305 354.815 694.475 354.985 ;
        RECT 694.785 354.815 694.955 354.985 ;
        RECT 695.265 354.815 695.435 354.985 ;
        RECT 695.745 354.815 695.915 354.985 ;
        RECT 696.225 354.815 696.395 354.985 ;
        RECT 696.705 354.815 696.875 354.985 ;
        RECT 697.185 354.815 697.355 354.985 ;
        RECT 697.665 354.815 697.835 354.985 ;
        RECT 698.145 354.815 698.315 354.985 ;
        RECT 698.625 354.815 698.795 354.985 ;
        RECT 699.105 354.815 699.275 354.985 ;
        RECT 699.585 354.815 699.755 354.985 ;
        RECT 700.065 354.815 700.235 354.985 ;
        RECT 700.545 354.815 700.715 354.985 ;
        RECT 701.025 354.815 701.195 354.985 ;
        RECT 701.505 354.815 701.675 354.985 ;
        RECT 701.985 354.815 702.155 354.985 ;
        RECT 702.465 354.815 702.635 354.985 ;
        RECT 702.945 354.815 703.115 354.985 ;
        RECT 703.425 354.815 703.595 354.985 ;
        RECT 703.905 354.815 704.075 354.985 ;
        RECT 704.385 354.815 704.555 354.985 ;
        RECT 704.865 354.815 705.035 354.985 ;
        RECT 705.345 354.815 705.515 354.985 ;
        RECT 705.825 354.815 705.995 354.985 ;
        RECT 706.305 354.815 706.475 354.985 ;
        RECT 706.785 354.815 706.955 354.985 ;
        RECT 707.265 354.815 707.435 354.985 ;
        RECT 707.745 354.815 707.915 354.985 ;
        RECT 708.225 354.815 708.395 354.985 ;
        RECT 693.860 354.335 694.030 354.505 ;
        RECT 694.220 354.335 694.390 354.505 ;
        RECT 694.580 354.335 694.750 354.505 ;
        RECT 695.390 354.335 695.560 354.505 ;
        RECT 695.750 354.335 695.920 354.505 ;
        RECT 696.110 354.335 696.280 354.505 ;
        RECT 697.145 354.335 697.315 354.505 ;
        RECT 697.505 354.335 697.675 354.505 ;
        RECT 697.865 354.335 698.035 354.505 ;
        RECT 699.840 354.335 700.010 354.505 ;
        RECT 700.200 354.335 700.370 354.505 ;
        RECT 700.560 354.335 700.730 354.505 ;
        RECT 702.180 354.335 702.350 354.505 ;
        RECT 702.540 354.335 702.710 354.505 ;
        RECT 702.900 354.335 703.070 354.505 ;
        RECT 705.330 354.335 705.500 354.505 ;
        RECT 707.360 354.335 707.530 354.505 ;
        RECT 707.720 354.335 707.890 354.505 ;
        RECT 711.195 354.815 711.365 354.985 ;
        RECT 711.675 354.815 711.845 354.985 ;
        RECT 712.155 354.815 712.325 354.985 ;
        RECT 712.635 354.815 712.805 354.985 ;
        RECT 713.115 354.815 713.285 354.985 ;
        RECT 713.595 354.815 713.765 354.985 ;
        RECT 714.075 354.815 714.245 354.985 ;
        RECT 714.555 354.815 714.725 354.985 ;
        RECT 715.035 354.815 715.205 354.985 ;
        RECT 715.515 354.815 715.685 354.985 ;
        RECT 715.995 354.815 716.165 354.985 ;
        RECT 716.475 354.815 716.645 354.985 ;
        RECT 716.955 354.815 717.125 354.985 ;
        RECT 717.435 354.815 717.605 354.985 ;
        RECT 717.915 354.815 718.085 354.985 ;
        RECT 718.395 354.815 718.565 354.985 ;
        RECT 718.875 354.815 719.045 354.985 ;
        RECT 719.355 354.815 719.525 354.985 ;
        RECT 719.835 354.815 720.005 354.985 ;
        RECT 720.315 354.815 720.485 354.985 ;
        RECT 720.795 354.815 720.965 354.985 ;
        RECT 721.275 354.815 721.445 354.985 ;
        RECT 721.755 354.815 721.925 354.985 ;
        RECT 722.235 354.815 722.405 354.985 ;
        RECT 722.715 354.815 722.885 354.985 ;
        RECT 723.195 354.815 723.365 354.985 ;
        RECT 723.675 354.815 723.845 354.985 ;
        RECT 724.155 354.815 724.325 354.985 ;
        RECT 724.635 354.815 724.805 354.985 ;
        RECT 725.115 354.815 725.285 354.985 ;
        RECT 725.595 354.815 725.765 354.985 ;
        RECT 726.075 354.815 726.245 354.985 ;
        RECT 711.710 354.335 711.880 354.505 ;
        RECT 712.070 354.335 712.240 354.505 ;
        RECT 712.430 354.335 712.600 354.505 ;
        RECT 713.240 354.335 713.410 354.505 ;
        RECT 713.600 354.335 713.770 354.505 ;
        RECT 713.960 354.335 714.130 354.505 ;
        RECT 714.995 354.335 715.165 354.505 ;
        RECT 715.355 354.335 715.525 354.505 ;
        RECT 715.715 354.335 715.885 354.505 ;
        RECT 717.690 354.335 717.860 354.505 ;
        RECT 718.050 354.335 718.220 354.505 ;
        RECT 718.410 354.335 718.580 354.505 ;
        RECT 720.030 354.335 720.200 354.505 ;
        RECT 720.390 354.335 720.560 354.505 ;
        RECT 720.750 354.335 720.920 354.505 ;
        RECT 723.180 354.335 723.350 354.505 ;
        RECT 725.210 354.335 725.380 354.505 ;
        RECT 725.570 354.335 725.740 354.505 ;
        RECT 729.455 354.815 729.625 354.985 ;
        RECT 729.935 354.815 730.105 354.985 ;
        RECT 730.415 354.815 730.585 354.985 ;
        RECT 730.895 354.815 731.065 354.985 ;
        RECT 731.375 354.815 731.545 354.985 ;
        RECT 731.855 354.815 732.025 354.985 ;
        RECT 732.335 354.815 732.505 354.985 ;
        RECT 732.815 354.815 732.985 354.985 ;
        RECT 733.295 354.815 733.465 354.985 ;
        RECT 733.775 354.815 733.945 354.985 ;
        RECT 734.255 354.815 734.425 354.985 ;
        RECT 734.735 354.815 734.905 354.985 ;
        RECT 735.215 354.815 735.385 354.985 ;
        RECT 735.695 354.815 735.865 354.985 ;
        RECT 736.175 354.815 736.345 354.985 ;
        RECT 736.655 354.815 736.825 354.985 ;
        RECT 737.135 354.815 737.305 354.985 ;
        RECT 737.615 354.815 737.785 354.985 ;
        RECT 738.095 354.815 738.265 354.985 ;
        RECT 738.575 354.815 738.745 354.985 ;
        RECT 739.055 354.815 739.225 354.985 ;
        RECT 739.535 354.815 739.705 354.985 ;
        RECT 740.015 354.815 740.185 354.985 ;
        RECT 740.495 354.815 740.665 354.985 ;
        RECT 740.975 354.815 741.145 354.985 ;
        RECT 741.455 354.815 741.625 354.985 ;
        RECT 741.935 354.815 742.105 354.985 ;
        RECT 742.415 354.815 742.585 354.985 ;
        RECT 742.895 354.815 743.065 354.985 ;
        RECT 743.375 354.815 743.545 354.985 ;
        RECT 743.855 354.815 744.025 354.985 ;
        RECT 744.335 354.815 744.505 354.985 ;
        RECT 729.970 354.335 730.140 354.505 ;
        RECT 730.330 354.335 730.500 354.505 ;
        RECT 730.690 354.335 730.860 354.505 ;
        RECT 731.500 354.335 731.670 354.505 ;
        RECT 731.860 354.335 732.030 354.505 ;
        RECT 732.220 354.335 732.390 354.505 ;
        RECT 733.255 354.335 733.425 354.505 ;
        RECT 733.615 354.335 733.785 354.505 ;
        RECT 733.975 354.335 734.145 354.505 ;
        RECT 735.950 354.335 736.120 354.505 ;
        RECT 736.310 354.335 736.480 354.505 ;
        RECT 736.670 354.335 736.840 354.505 ;
        RECT 738.290 354.335 738.460 354.505 ;
        RECT 738.650 354.335 738.820 354.505 ;
        RECT 739.010 354.335 739.180 354.505 ;
        RECT 741.440 354.335 741.610 354.505 ;
        RECT 743.470 354.335 743.640 354.505 ;
        RECT 743.830 354.335 744.000 354.505 ;
        RECT 747.225 354.785 747.395 354.955 ;
        RECT 747.705 354.785 747.875 354.955 ;
        RECT 748.185 354.785 748.355 354.955 ;
        RECT 748.665 354.785 748.835 354.955 ;
        RECT 749.145 354.785 749.315 354.955 ;
        RECT 749.625 354.785 749.795 354.955 ;
        RECT 750.105 354.785 750.275 354.955 ;
        RECT 750.585 354.785 750.755 354.955 ;
        RECT 751.065 354.785 751.235 354.955 ;
        RECT 751.545 354.785 751.715 354.955 ;
        RECT 752.025 354.785 752.195 354.955 ;
        RECT 752.505 354.785 752.675 354.955 ;
        RECT 752.985 354.785 753.155 354.955 ;
        RECT 753.465 354.785 753.635 354.955 ;
        RECT 753.945 354.785 754.115 354.955 ;
        RECT 754.425 354.785 754.595 354.955 ;
        RECT 754.905 354.785 755.075 354.955 ;
        RECT 755.385 354.785 755.555 354.955 ;
        RECT 755.865 354.785 756.035 354.955 ;
        RECT 756.345 354.785 756.515 354.955 ;
        RECT 756.825 354.785 756.995 354.955 ;
        RECT 757.305 354.785 757.475 354.955 ;
        RECT 757.785 354.785 757.955 354.955 ;
        RECT 758.265 354.785 758.435 354.955 ;
        RECT 758.745 354.785 758.915 354.955 ;
        RECT 759.225 354.785 759.395 354.955 ;
        RECT 759.705 354.785 759.875 354.955 ;
        RECT 760.185 354.785 760.355 354.955 ;
        RECT 760.665 354.785 760.835 354.955 ;
        RECT 761.145 354.785 761.315 354.955 ;
        RECT 761.625 354.785 761.795 354.955 ;
        RECT 762.105 354.785 762.275 354.955 ;
        RECT 747.740 354.305 747.910 354.475 ;
        RECT 748.100 354.305 748.270 354.475 ;
        RECT 748.460 354.305 748.630 354.475 ;
        RECT 749.270 354.305 749.440 354.475 ;
        RECT 749.630 354.305 749.800 354.475 ;
        RECT 749.990 354.305 750.160 354.475 ;
        RECT 751.025 354.305 751.195 354.475 ;
        RECT 751.385 354.305 751.555 354.475 ;
        RECT 751.745 354.305 751.915 354.475 ;
        RECT 753.720 354.305 753.890 354.475 ;
        RECT 754.080 354.305 754.250 354.475 ;
        RECT 754.440 354.305 754.610 354.475 ;
        RECT 756.060 354.305 756.230 354.475 ;
        RECT 756.420 354.305 756.590 354.475 ;
        RECT 756.780 354.305 756.950 354.475 ;
        RECT 759.210 354.305 759.380 354.475 ;
        RECT 761.240 354.305 761.410 354.475 ;
        RECT 761.600 354.305 761.770 354.475 ;
        RECT 765.265 354.705 765.435 354.875 ;
        RECT 765.745 354.705 765.915 354.875 ;
        RECT 766.225 354.705 766.395 354.875 ;
        RECT 766.705 354.705 766.875 354.875 ;
        RECT 767.185 354.705 767.355 354.875 ;
        RECT 767.665 354.705 767.835 354.875 ;
        RECT 768.145 354.705 768.315 354.875 ;
        RECT 768.625 354.705 768.795 354.875 ;
        RECT 769.105 354.705 769.275 354.875 ;
        RECT 769.585 354.705 769.755 354.875 ;
        RECT 770.065 354.705 770.235 354.875 ;
        RECT 770.545 354.705 770.715 354.875 ;
        RECT 771.025 354.705 771.195 354.875 ;
        RECT 771.505 354.705 771.675 354.875 ;
        RECT 771.985 354.705 772.155 354.875 ;
        RECT 772.465 354.705 772.635 354.875 ;
        RECT 772.945 354.705 773.115 354.875 ;
        RECT 773.425 354.705 773.595 354.875 ;
        RECT 773.905 354.705 774.075 354.875 ;
        RECT 774.385 354.705 774.555 354.875 ;
        RECT 774.865 354.705 775.035 354.875 ;
        RECT 775.345 354.705 775.515 354.875 ;
        RECT 775.825 354.705 775.995 354.875 ;
        RECT 776.305 354.705 776.475 354.875 ;
        RECT 776.785 354.705 776.955 354.875 ;
        RECT 777.265 354.705 777.435 354.875 ;
        RECT 777.745 354.705 777.915 354.875 ;
        RECT 778.225 354.705 778.395 354.875 ;
        RECT 778.705 354.705 778.875 354.875 ;
        RECT 779.185 354.705 779.355 354.875 ;
        RECT 779.665 354.705 779.835 354.875 ;
        RECT 780.145 354.705 780.315 354.875 ;
        RECT 765.780 354.225 765.950 354.395 ;
        RECT 766.140 354.225 766.310 354.395 ;
        RECT 766.500 354.225 766.670 354.395 ;
        RECT 767.310 354.225 767.480 354.395 ;
        RECT 767.670 354.225 767.840 354.395 ;
        RECT 768.030 354.225 768.200 354.395 ;
        RECT 769.065 354.225 769.235 354.395 ;
        RECT 769.425 354.225 769.595 354.395 ;
        RECT 769.785 354.225 769.955 354.395 ;
        RECT 771.760 354.225 771.930 354.395 ;
        RECT 772.120 354.225 772.290 354.395 ;
        RECT 772.480 354.225 772.650 354.395 ;
        RECT 774.100 354.225 774.270 354.395 ;
        RECT 774.460 354.225 774.630 354.395 ;
        RECT 774.820 354.225 774.990 354.395 ;
        RECT 777.250 354.225 777.420 354.395 ;
        RECT 779.280 354.225 779.450 354.395 ;
        RECT 779.640 354.225 779.810 354.395 ;
        RECT 783.425 354.745 783.595 354.915 ;
        RECT 783.905 354.745 784.075 354.915 ;
        RECT 784.385 354.745 784.555 354.915 ;
        RECT 784.865 354.745 785.035 354.915 ;
        RECT 785.345 354.745 785.515 354.915 ;
        RECT 785.825 354.745 785.995 354.915 ;
        RECT 786.305 354.745 786.475 354.915 ;
        RECT 786.785 354.745 786.955 354.915 ;
        RECT 787.265 354.745 787.435 354.915 ;
        RECT 787.745 354.745 787.915 354.915 ;
        RECT 788.225 354.745 788.395 354.915 ;
        RECT 788.705 354.745 788.875 354.915 ;
        RECT 789.185 354.745 789.355 354.915 ;
        RECT 789.665 354.745 789.835 354.915 ;
        RECT 790.145 354.745 790.315 354.915 ;
        RECT 790.625 354.745 790.795 354.915 ;
        RECT 791.105 354.745 791.275 354.915 ;
        RECT 791.585 354.745 791.755 354.915 ;
        RECT 792.065 354.745 792.235 354.915 ;
        RECT 792.545 354.745 792.715 354.915 ;
        RECT 793.025 354.745 793.195 354.915 ;
        RECT 793.505 354.745 793.675 354.915 ;
        RECT 793.985 354.745 794.155 354.915 ;
        RECT 794.465 354.745 794.635 354.915 ;
        RECT 794.945 354.745 795.115 354.915 ;
        RECT 795.425 354.745 795.595 354.915 ;
        RECT 795.905 354.745 796.075 354.915 ;
        RECT 796.385 354.745 796.555 354.915 ;
        RECT 796.865 354.745 797.035 354.915 ;
        RECT 797.345 354.745 797.515 354.915 ;
        RECT 797.825 354.745 797.995 354.915 ;
        RECT 798.305 354.745 798.475 354.915 ;
        RECT 783.940 354.265 784.110 354.435 ;
        RECT 784.300 354.265 784.470 354.435 ;
        RECT 784.660 354.265 784.830 354.435 ;
        RECT 785.470 354.265 785.640 354.435 ;
        RECT 785.830 354.265 786.000 354.435 ;
        RECT 786.190 354.265 786.360 354.435 ;
        RECT 787.225 354.265 787.395 354.435 ;
        RECT 787.585 354.265 787.755 354.435 ;
        RECT 787.945 354.265 788.115 354.435 ;
        RECT 789.920 354.265 790.090 354.435 ;
        RECT 790.280 354.265 790.450 354.435 ;
        RECT 790.640 354.265 790.810 354.435 ;
        RECT 792.260 354.265 792.430 354.435 ;
        RECT 792.620 354.265 792.790 354.435 ;
        RECT 792.980 354.265 793.150 354.435 ;
        RECT 795.410 354.265 795.580 354.435 ;
        RECT 797.440 354.265 797.610 354.435 ;
        RECT 797.800 354.265 797.970 354.435 ;
        RECT 801.805 354.755 801.975 354.925 ;
        RECT 802.285 354.755 802.455 354.925 ;
        RECT 802.765 354.755 802.935 354.925 ;
        RECT 803.245 354.755 803.415 354.925 ;
        RECT 803.725 354.755 803.895 354.925 ;
        RECT 804.205 354.755 804.375 354.925 ;
        RECT 804.685 354.755 804.855 354.925 ;
        RECT 805.165 354.755 805.335 354.925 ;
        RECT 805.645 354.755 805.815 354.925 ;
        RECT 806.125 354.755 806.295 354.925 ;
        RECT 806.605 354.755 806.775 354.925 ;
        RECT 807.085 354.755 807.255 354.925 ;
        RECT 807.565 354.755 807.735 354.925 ;
        RECT 808.045 354.755 808.215 354.925 ;
        RECT 808.525 354.755 808.695 354.925 ;
        RECT 809.005 354.755 809.175 354.925 ;
        RECT 809.485 354.755 809.655 354.925 ;
        RECT 809.965 354.755 810.135 354.925 ;
        RECT 810.445 354.755 810.615 354.925 ;
        RECT 810.925 354.755 811.095 354.925 ;
        RECT 811.405 354.755 811.575 354.925 ;
        RECT 811.885 354.755 812.055 354.925 ;
        RECT 812.365 354.755 812.535 354.925 ;
        RECT 812.845 354.755 813.015 354.925 ;
        RECT 813.325 354.755 813.495 354.925 ;
        RECT 813.805 354.755 813.975 354.925 ;
        RECT 814.285 354.755 814.455 354.925 ;
        RECT 814.765 354.755 814.935 354.925 ;
        RECT 815.245 354.755 815.415 354.925 ;
        RECT 815.725 354.755 815.895 354.925 ;
        RECT 816.205 354.755 816.375 354.925 ;
        RECT 816.685 354.755 816.855 354.925 ;
        RECT 802.320 354.275 802.490 354.445 ;
        RECT 802.680 354.275 802.850 354.445 ;
        RECT 803.040 354.275 803.210 354.445 ;
        RECT 803.850 354.275 804.020 354.445 ;
        RECT 804.210 354.275 804.380 354.445 ;
        RECT 804.570 354.275 804.740 354.445 ;
        RECT 805.605 354.275 805.775 354.445 ;
        RECT 805.965 354.275 806.135 354.445 ;
        RECT 806.325 354.275 806.495 354.445 ;
        RECT 808.300 354.275 808.470 354.445 ;
        RECT 808.660 354.275 808.830 354.445 ;
        RECT 809.020 354.275 809.190 354.445 ;
        RECT 810.640 354.275 810.810 354.445 ;
        RECT 811.000 354.275 811.170 354.445 ;
        RECT 811.360 354.275 811.530 354.445 ;
        RECT 813.790 354.275 813.960 354.445 ;
        RECT 815.820 354.275 815.990 354.445 ;
        RECT 816.180 354.275 816.350 354.445 ;
        RECT 820.605 354.735 820.775 354.905 ;
        RECT 821.085 354.735 821.255 354.905 ;
        RECT 821.565 354.735 821.735 354.905 ;
        RECT 822.045 354.735 822.215 354.905 ;
        RECT 822.525 354.735 822.695 354.905 ;
        RECT 823.005 354.735 823.175 354.905 ;
        RECT 823.485 354.735 823.655 354.905 ;
        RECT 823.965 354.735 824.135 354.905 ;
        RECT 824.445 354.735 824.615 354.905 ;
        RECT 824.925 354.735 825.095 354.905 ;
        RECT 825.405 354.735 825.575 354.905 ;
        RECT 825.885 354.735 826.055 354.905 ;
        RECT 826.365 354.735 826.535 354.905 ;
        RECT 826.845 354.735 827.015 354.905 ;
        RECT 827.325 354.735 827.495 354.905 ;
        RECT 827.805 354.735 827.975 354.905 ;
        RECT 828.285 354.735 828.455 354.905 ;
        RECT 828.765 354.735 828.935 354.905 ;
        RECT 829.245 354.735 829.415 354.905 ;
        RECT 829.725 354.735 829.895 354.905 ;
        RECT 830.205 354.735 830.375 354.905 ;
        RECT 830.685 354.735 830.855 354.905 ;
        RECT 831.165 354.735 831.335 354.905 ;
        RECT 831.645 354.735 831.815 354.905 ;
        RECT 832.125 354.735 832.295 354.905 ;
        RECT 832.605 354.735 832.775 354.905 ;
        RECT 833.085 354.735 833.255 354.905 ;
        RECT 833.565 354.735 833.735 354.905 ;
        RECT 834.045 354.735 834.215 354.905 ;
        RECT 834.525 354.735 834.695 354.905 ;
        RECT 835.005 354.735 835.175 354.905 ;
        RECT 835.485 354.735 835.655 354.905 ;
        RECT 821.120 354.255 821.290 354.425 ;
        RECT 821.480 354.255 821.650 354.425 ;
        RECT 821.840 354.255 822.010 354.425 ;
        RECT 822.650 354.255 822.820 354.425 ;
        RECT 823.010 354.255 823.180 354.425 ;
        RECT 823.370 354.255 823.540 354.425 ;
        RECT 824.405 354.255 824.575 354.425 ;
        RECT 824.765 354.255 824.935 354.425 ;
        RECT 825.125 354.255 825.295 354.425 ;
        RECT 827.100 354.255 827.270 354.425 ;
        RECT 827.460 354.255 827.630 354.425 ;
        RECT 827.820 354.255 827.990 354.425 ;
        RECT 829.440 354.255 829.610 354.425 ;
        RECT 829.800 354.255 829.970 354.425 ;
        RECT 830.160 354.255 830.330 354.425 ;
        RECT 832.590 354.255 832.760 354.425 ;
        RECT 834.620 354.255 834.790 354.425 ;
        RECT 834.980 354.255 835.150 354.425 ;
        RECT 839.075 354.715 839.245 354.885 ;
        RECT 839.555 354.715 839.725 354.885 ;
        RECT 840.035 354.715 840.205 354.885 ;
        RECT 839.710 354.235 839.880 354.405 ;
        RECT 840.070 354.235 840.240 354.405 ;
        RECT 832.145 352.045 832.315 352.215 ;
        RECT 398.410 351.025 398.580 351.195 ;
        RECT 401.700 351.025 401.870 351.195 ;
        RECT 404.990 351.025 405.160 351.195 ;
        RECT 408.280 351.385 408.450 351.555 ;
        RECT 408.280 351.025 408.450 351.195 ;
        RECT 389.010 346.315 389.180 346.485 ;
        RECT 382.430 345.955 382.600 346.125 ;
        RECT 382.430 342.845 382.600 343.015 ;
        RECT 382.430 342.485 382.600 342.655 ;
        RECT 382.430 339.375 382.600 339.545 ;
        RECT 382.430 339.015 382.600 339.185 ;
        RECT 382.430 335.905 382.600 336.075 ;
        RECT 382.430 335.545 382.600 335.715 ;
        RECT 375.850 332.435 376.020 332.605 ;
        RECT 369.690 332.175 369.860 332.345 ;
        RECT 382.430 332.435 382.600 332.605 ;
        RECT 389.010 345.955 389.180 346.125 ;
        RECT 389.010 342.845 389.180 343.015 ;
        RECT 389.010 342.485 389.180 342.655 ;
        RECT 389.010 339.375 389.180 339.545 ;
        RECT 389.010 339.015 389.180 339.185 ;
        RECT 389.010 335.905 389.180 336.075 ;
        RECT 389.010 335.545 389.180 335.715 ;
        RECT 389.010 332.435 389.180 332.605 ;
        RECT 375.850 332.075 376.020 332.245 ;
        RECT 98.025 327.930 98.195 328.100 ;
        RECT 98.385 327.930 98.555 328.100 ;
        RECT 101.495 327.930 101.665 328.100 ;
        RECT 101.855 327.930 102.025 328.100 ;
        RECT 4.995 327.680 5.165 327.850 ;
        RECT 5.355 327.680 5.525 327.850 ;
        RECT 8.465 327.680 8.635 327.850 ;
        RECT 8.825 327.680 8.995 327.850 ;
        RECT 11.935 327.680 12.105 327.850 ;
        RECT 12.295 327.680 12.465 327.850 ;
        RECT 18.335 327.660 18.505 327.830 ;
        RECT 18.695 327.660 18.865 327.830 ;
        RECT 21.805 327.660 21.975 327.830 ;
        RECT 22.165 327.660 22.335 327.830 ;
        RECT 25.275 327.660 25.445 327.830 ;
        RECT 25.635 327.660 25.805 327.830 ;
        RECT 31.705 327.690 31.875 327.860 ;
        RECT 32.065 327.690 32.235 327.860 ;
        RECT 35.175 327.690 35.345 327.860 ;
        RECT 35.535 327.690 35.705 327.860 ;
        RECT 38.645 327.690 38.815 327.860 ;
        RECT 39.005 327.690 39.175 327.860 ;
        RECT 44.935 327.690 45.105 327.860 ;
        RECT 45.295 327.690 45.465 327.860 ;
        RECT 48.405 327.690 48.575 327.860 ;
        RECT 48.765 327.690 48.935 327.860 ;
        RECT 51.875 327.690 52.045 327.860 ;
        RECT 52.235 327.690 52.405 327.860 ;
        RECT 58.205 327.660 58.375 327.830 ;
        RECT 58.565 327.660 58.735 327.830 ;
        RECT 61.675 327.660 61.845 327.830 ;
        RECT 62.035 327.660 62.205 327.830 ;
        RECT 65.145 327.660 65.315 327.830 ;
        RECT 65.505 327.660 65.675 327.830 ;
        RECT 71.475 327.690 71.645 327.860 ;
        RECT 71.835 327.690 72.005 327.860 ;
        RECT 74.945 327.690 75.115 327.860 ;
        RECT 75.305 327.690 75.475 327.860 ;
        RECT 78.415 327.690 78.585 327.860 ;
        RECT 78.775 327.690 78.945 327.860 ;
        RECT 84.605 327.710 84.775 327.880 ;
        RECT 84.965 327.710 85.135 327.880 ;
        RECT 88.075 327.710 88.245 327.880 ;
        RECT 88.435 327.710 88.605 327.880 ;
        RECT 91.545 327.710 91.715 327.880 ;
        RECT 91.905 327.710 92.075 327.880 ;
        RECT 4.995 324.390 5.165 324.560 ;
        RECT 5.355 324.390 5.525 324.560 ;
        RECT 8.465 324.390 8.635 324.560 ;
        RECT 8.825 324.390 8.995 324.560 ;
        RECT 11.935 324.390 12.105 324.560 ;
        RECT 12.295 324.390 12.465 324.560 ;
        RECT 4.995 321.100 5.165 321.270 ;
        RECT 5.355 321.100 5.525 321.270 ;
        RECT 8.465 321.100 8.635 321.270 ;
        RECT 8.825 321.100 8.995 321.270 ;
        RECT 11.935 321.100 12.105 321.270 ;
        RECT 12.295 321.100 12.465 321.270 ;
        RECT 4.995 317.810 5.165 317.980 ;
        RECT 5.355 317.810 5.525 317.980 ;
        RECT 8.465 317.810 8.635 317.980 ;
        RECT 8.825 317.810 8.995 317.980 ;
        RECT 11.935 317.810 12.105 317.980 ;
        RECT 12.295 317.810 12.465 317.980 ;
        RECT 4.995 314.520 5.165 314.690 ;
        RECT 5.355 314.520 5.525 314.690 ;
        RECT 8.465 314.520 8.635 314.690 ;
        RECT 8.825 314.520 8.995 314.690 ;
        RECT 11.935 314.520 12.105 314.690 ;
        RECT 12.295 314.520 12.465 314.690 ;
        RECT 4.995 311.230 5.165 311.400 ;
        RECT 5.355 311.230 5.525 311.400 ;
        RECT 8.465 311.230 8.635 311.400 ;
        RECT 8.825 311.230 8.995 311.400 ;
        RECT 11.935 311.230 12.105 311.400 ;
        RECT 12.295 311.230 12.465 311.400 ;
        RECT 18.335 324.370 18.505 324.540 ;
        RECT 18.695 324.370 18.865 324.540 ;
        RECT 21.805 324.370 21.975 324.540 ;
        RECT 22.165 324.370 22.335 324.540 ;
        RECT 25.275 324.370 25.445 324.540 ;
        RECT 25.635 324.370 25.805 324.540 ;
        RECT 18.335 321.080 18.505 321.250 ;
        RECT 18.695 321.080 18.865 321.250 ;
        RECT 21.805 321.080 21.975 321.250 ;
        RECT 22.165 321.080 22.335 321.250 ;
        RECT 25.275 321.080 25.445 321.250 ;
        RECT 25.635 321.080 25.805 321.250 ;
        RECT 18.335 317.790 18.505 317.960 ;
        RECT 18.695 317.790 18.865 317.960 ;
        RECT 21.805 317.790 21.975 317.960 ;
        RECT 22.165 317.790 22.335 317.960 ;
        RECT 25.275 317.790 25.445 317.960 ;
        RECT 25.635 317.790 25.805 317.960 ;
        RECT 18.335 314.500 18.505 314.670 ;
        RECT 18.695 314.500 18.865 314.670 ;
        RECT 21.805 314.500 21.975 314.670 ;
        RECT 22.165 314.500 22.335 314.670 ;
        RECT 25.275 314.500 25.445 314.670 ;
        RECT 25.635 314.500 25.805 314.670 ;
        RECT 18.335 311.210 18.505 311.380 ;
        RECT 18.695 311.210 18.865 311.380 ;
        RECT 21.805 311.210 21.975 311.380 ;
        RECT 22.165 311.210 22.335 311.380 ;
        RECT 25.275 311.210 25.445 311.380 ;
        RECT 25.635 311.210 25.805 311.380 ;
        RECT 4.995 307.940 5.165 308.110 ;
        RECT 5.355 307.940 5.525 308.110 ;
        RECT 8.465 307.940 8.635 308.110 ;
        RECT 8.825 307.940 8.995 308.110 ;
        RECT 11.935 307.940 12.105 308.110 ;
        RECT 12.295 307.940 12.465 308.110 ;
        RECT 4.995 304.650 5.165 304.820 ;
        RECT 5.355 304.650 5.525 304.820 ;
        RECT 8.465 304.650 8.635 304.820 ;
        RECT 8.825 304.650 8.995 304.820 ;
        RECT 11.935 304.650 12.105 304.820 ;
        RECT 12.295 304.650 12.465 304.820 ;
        RECT 15.530 303.660 16.420 305.270 ;
        RECT 31.705 324.400 31.875 324.570 ;
        RECT 32.065 324.400 32.235 324.570 ;
        RECT 35.175 324.400 35.345 324.570 ;
        RECT 35.535 324.400 35.705 324.570 ;
        RECT 38.645 324.400 38.815 324.570 ;
        RECT 39.005 324.400 39.175 324.570 ;
        RECT 31.705 321.110 31.875 321.280 ;
        RECT 32.065 321.110 32.235 321.280 ;
        RECT 35.175 321.110 35.345 321.280 ;
        RECT 35.535 321.110 35.705 321.280 ;
        RECT 38.645 321.110 38.815 321.280 ;
        RECT 39.005 321.110 39.175 321.280 ;
        RECT 31.705 317.820 31.875 317.990 ;
        RECT 32.065 317.820 32.235 317.990 ;
        RECT 35.175 317.820 35.345 317.990 ;
        RECT 35.535 317.820 35.705 317.990 ;
        RECT 38.645 317.820 38.815 317.990 ;
        RECT 39.005 317.820 39.175 317.990 ;
        RECT 31.705 314.530 31.875 314.700 ;
        RECT 32.065 314.530 32.235 314.700 ;
        RECT 35.175 314.530 35.345 314.700 ;
        RECT 35.535 314.530 35.705 314.700 ;
        RECT 38.645 314.530 38.815 314.700 ;
        RECT 39.005 314.530 39.175 314.700 ;
        RECT 31.705 311.240 31.875 311.410 ;
        RECT 32.065 311.240 32.235 311.410 ;
        RECT 35.175 311.240 35.345 311.410 ;
        RECT 35.535 311.240 35.705 311.410 ;
        RECT 38.645 311.240 38.815 311.410 ;
        RECT 39.005 311.240 39.175 311.410 ;
        RECT 18.335 307.920 18.505 308.090 ;
        RECT 18.695 307.920 18.865 308.090 ;
        RECT 21.805 307.920 21.975 308.090 ;
        RECT 22.165 307.920 22.335 308.090 ;
        RECT 25.275 307.920 25.445 308.090 ;
        RECT 25.635 307.920 25.805 308.090 ;
        RECT 18.335 304.630 18.505 304.800 ;
        RECT 18.695 304.630 18.865 304.800 ;
        RECT 21.805 304.630 21.975 304.800 ;
        RECT 22.165 304.630 22.335 304.800 ;
        RECT 25.275 304.630 25.445 304.800 ;
        RECT 25.635 304.630 25.805 304.800 ;
        RECT 28.745 303.810 29.635 305.420 ;
        RECT 44.935 324.400 45.105 324.570 ;
        RECT 45.295 324.400 45.465 324.570 ;
        RECT 48.405 324.400 48.575 324.570 ;
        RECT 48.765 324.400 48.935 324.570 ;
        RECT 51.875 324.400 52.045 324.570 ;
        RECT 52.235 324.400 52.405 324.570 ;
        RECT 44.935 321.110 45.105 321.280 ;
        RECT 45.295 321.110 45.465 321.280 ;
        RECT 48.405 321.110 48.575 321.280 ;
        RECT 48.765 321.110 48.935 321.280 ;
        RECT 51.875 321.110 52.045 321.280 ;
        RECT 52.235 321.110 52.405 321.280 ;
        RECT 44.935 317.820 45.105 317.990 ;
        RECT 45.295 317.820 45.465 317.990 ;
        RECT 48.405 317.820 48.575 317.990 ;
        RECT 48.765 317.820 48.935 317.990 ;
        RECT 51.875 317.820 52.045 317.990 ;
        RECT 52.235 317.820 52.405 317.990 ;
        RECT 44.935 314.530 45.105 314.700 ;
        RECT 45.295 314.530 45.465 314.700 ;
        RECT 48.405 314.530 48.575 314.700 ;
        RECT 48.765 314.530 48.935 314.700 ;
        RECT 51.875 314.530 52.045 314.700 ;
        RECT 52.235 314.530 52.405 314.700 ;
        RECT 44.935 311.240 45.105 311.410 ;
        RECT 45.295 311.240 45.465 311.410 ;
        RECT 48.405 311.240 48.575 311.410 ;
        RECT 48.765 311.240 48.935 311.410 ;
        RECT 51.875 311.240 52.045 311.410 ;
        RECT 52.235 311.240 52.405 311.410 ;
        RECT 31.705 307.950 31.875 308.120 ;
        RECT 32.065 307.950 32.235 308.120 ;
        RECT 35.175 307.950 35.345 308.120 ;
        RECT 35.535 307.950 35.705 308.120 ;
        RECT 38.645 307.950 38.815 308.120 ;
        RECT 39.005 307.950 39.175 308.120 ;
        RECT 31.705 304.660 31.875 304.830 ;
        RECT 32.065 304.660 32.235 304.830 ;
        RECT 35.175 304.660 35.345 304.830 ;
        RECT 35.535 304.660 35.705 304.830 ;
        RECT 38.645 304.660 38.815 304.830 ;
        RECT 39.005 304.660 39.175 304.830 ;
        RECT 41.960 303.515 42.850 305.845 ;
        RECT 58.205 324.370 58.375 324.540 ;
        RECT 58.565 324.370 58.735 324.540 ;
        RECT 61.675 324.370 61.845 324.540 ;
        RECT 62.035 324.370 62.205 324.540 ;
        RECT 65.145 324.370 65.315 324.540 ;
        RECT 65.505 324.370 65.675 324.540 ;
        RECT 58.205 321.080 58.375 321.250 ;
        RECT 58.565 321.080 58.735 321.250 ;
        RECT 61.675 321.080 61.845 321.250 ;
        RECT 62.035 321.080 62.205 321.250 ;
        RECT 65.145 321.080 65.315 321.250 ;
        RECT 65.505 321.080 65.675 321.250 ;
        RECT 58.205 317.790 58.375 317.960 ;
        RECT 58.565 317.790 58.735 317.960 ;
        RECT 61.675 317.790 61.845 317.960 ;
        RECT 62.035 317.790 62.205 317.960 ;
        RECT 65.145 317.790 65.315 317.960 ;
        RECT 65.505 317.790 65.675 317.960 ;
        RECT 58.205 314.500 58.375 314.670 ;
        RECT 58.565 314.500 58.735 314.670 ;
        RECT 61.675 314.500 61.845 314.670 ;
        RECT 62.035 314.500 62.205 314.670 ;
        RECT 65.145 314.500 65.315 314.670 ;
        RECT 65.505 314.500 65.675 314.670 ;
        RECT 58.205 311.210 58.375 311.380 ;
        RECT 58.565 311.210 58.735 311.380 ;
        RECT 61.675 311.210 61.845 311.380 ;
        RECT 62.035 311.210 62.205 311.380 ;
        RECT 65.145 311.210 65.315 311.380 ;
        RECT 65.505 311.210 65.675 311.380 ;
        RECT 44.935 307.950 45.105 308.120 ;
        RECT 45.295 307.950 45.465 308.120 ;
        RECT 48.405 307.950 48.575 308.120 ;
        RECT 48.765 307.950 48.935 308.120 ;
        RECT 51.875 307.950 52.045 308.120 ;
        RECT 52.235 307.950 52.405 308.120 ;
        RECT 44.935 304.660 45.105 304.830 ;
        RECT 45.295 304.660 45.465 304.830 ;
        RECT 48.405 304.660 48.575 304.830 ;
        RECT 48.765 304.660 48.935 304.830 ;
        RECT 51.875 304.660 52.045 304.830 ;
        RECT 52.235 304.660 52.405 304.830 ;
        RECT 55.380 303.400 56.270 305.370 ;
        RECT 71.475 324.400 71.645 324.570 ;
        RECT 71.835 324.400 72.005 324.570 ;
        RECT 74.945 324.400 75.115 324.570 ;
        RECT 75.305 324.400 75.475 324.570 ;
        RECT 78.415 324.400 78.585 324.570 ;
        RECT 78.775 324.400 78.945 324.570 ;
        RECT 71.475 321.110 71.645 321.280 ;
        RECT 71.835 321.110 72.005 321.280 ;
        RECT 74.945 321.110 75.115 321.280 ;
        RECT 75.305 321.110 75.475 321.280 ;
        RECT 78.415 321.110 78.585 321.280 ;
        RECT 78.775 321.110 78.945 321.280 ;
        RECT 71.475 317.820 71.645 317.990 ;
        RECT 71.835 317.820 72.005 317.990 ;
        RECT 74.945 317.820 75.115 317.990 ;
        RECT 75.305 317.820 75.475 317.990 ;
        RECT 78.415 317.820 78.585 317.990 ;
        RECT 78.775 317.820 78.945 317.990 ;
        RECT 71.475 314.530 71.645 314.700 ;
        RECT 71.835 314.530 72.005 314.700 ;
        RECT 74.945 314.530 75.115 314.700 ;
        RECT 75.305 314.530 75.475 314.700 ;
        RECT 78.415 314.530 78.585 314.700 ;
        RECT 78.775 314.530 78.945 314.700 ;
        RECT 71.475 311.240 71.645 311.410 ;
        RECT 71.835 311.240 72.005 311.410 ;
        RECT 74.945 311.240 75.115 311.410 ;
        RECT 75.305 311.240 75.475 311.410 ;
        RECT 78.415 311.240 78.585 311.410 ;
        RECT 78.775 311.240 78.945 311.410 ;
        RECT 58.205 307.920 58.375 308.090 ;
        RECT 58.565 307.920 58.735 308.090 ;
        RECT 61.675 307.920 61.845 308.090 ;
        RECT 62.035 307.920 62.205 308.090 ;
        RECT 65.145 307.920 65.315 308.090 ;
        RECT 65.505 307.920 65.675 308.090 ;
        RECT 58.205 304.630 58.375 304.800 ;
        RECT 58.565 304.630 58.735 304.800 ;
        RECT 61.675 304.630 61.845 304.800 ;
        RECT 62.035 304.630 62.205 304.800 ;
        RECT 65.145 304.630 65.315 304.800 ;
        RECT 65.505 304.630 65.675 304.800 ;
        RECT 68.685 303.585 69.215 305.555 ;
        RECT 84.605 324.420 84.775 324.590 ;
        RECT 84.965 324.420 85.135 324.590 ;
        RECT 88.075 324.420 88.245 324.590 ;
        RECT 88.435 324.420 88.605 324.590 ;
        RECT 91.545 324.420 91.715 324.590 ;
        RECT 91.905 324.420 92.075 324.590 ;
        RECT 355.435 326.965 355.605 327.135 ;
        RECT 355.435 326.605 355.605 326.775 ;
        RECT 355.435 326.245 355.605 326.415 ;
        RECT 355.435 325.885 355.605 326.055 ;
        RECT 355.435 325.525 355.605 325.695 ;
        RECT 98.025 324.640 98.195 324.810 ;
        RECT 98.385 324.640 98.555 324.810 ;
        RECT 101.495 324.640 101.665 324.810 ;
        RECT 101.855 324.640 102.025 324.810 ;
        RECT 84.605 321.130 84.775 321.300 ;
        RECT 84.965 321.130 85.135 321.300 ;
        RECT 88.075 321.130 88.245 321.300 ;
        RECT 88.435 321.130 88.605 321.300 ;
        RECT 91.545 321.130 91.715 321.300 ;
        RECT 91.905 321.130 92.075 321.300 ;
        RECT 84.605 317.840 84.775 318.010 ;
        RECT 84.965 317.840 85.135 318.010 ;
        RECT 88.075 317.840 88.245 318.010 ;
        RECT 88.435 317.840 88.605 318.010 ;
        RECT 91.545 317.840 91.715 318.010 ;
        RECT 91.905 317.840 92.075 318.010 ;
        RECT 84.605 314.550 84.775 314.720 ;
        RECT 84.965 314.550 85.135 314.720 ;
        RECT 88.075 314.550 88.245 314.720 ;
        RECT 88.435 314.550 88.605 314.720 ;
        RECT 91.545 314.550 91.715 314.720 ;
        RECT 91.905 314.550 92.075 314.720 ;
        RECT 84.605 311.260 84.775 311.430 ;
        RECT 84.965 311.260 85.135 311.430 ;
        RECT 88.075 311.260 88.245 311.430 ;
        RECT 88.435 311.260 88.605 311.430 ;
        RECT 91.545 311.260 91.715 311.430 ;
        RECT 91.905 311.260 92.075 311.430 ;
        RECT 71.475 307.950 71.645 308.120 ;
        RECT 71.835 307.950 72.005 308.120 ;
        RECT 74.945 307.950 75.115 308.120 ;
        RECT 75.305 307.950 75.475 308.120 ;
        RECT 78.415 307.950 78.585 308.120 ;
        RECT 78.775 307.950 78.945 308.120 ;
        RECT 71.475 304.660 71.645 304.830 ;
        RECT 71.835 304.660 72.005 304.830 ;
        RECT 74.945 304.660 75.115 304.830 ;
        RECT 75.305 304.660 75.475 304.830 ;
        RECT 78.415 304.660 78.585 304.830 ;
        RECT 78.775 304.660 78.945 304.830 ;
        RECT 81.620 304.050 82.870 305.300 ;
        RECT 215.290 324.090 225.900 324.980 ;
        RECT 235.330 324.080 245.940 324.970 ;
        RECT 255.390 324.080 266.000 324.970 ;
        RECT 275.440 324.080 286.050 324.970 ;
        RECT 355.435 325.165 355.605 325.335 ;
        RECT 355.435 324.805 355.605 324.975 ;
        RECT 355.435 324.445 355.605 324.615 ;
        RECT 355.435 324.085 355.605 324.255 ;
        RECT 355.435 323.725 355.605 323.895 ;
        RECT 355.435 323.365 355.605 323.535 ;
        RECT 355.435 323.005 355.605 323.175 ;
        RECT 212.115 322.610 212.285 322.780 ;
        RECT 212.475 322.610 212.645 322.780 ;
        RECT 215.585 322.610 215.755 322.780 ;
        RECT 215.945 322.610 216.115 322.780 ;
        RECT 219.055 322.610 219.225 322.780 ;
        RECT 219.415 322.610 219.585 322.780 ;
        RECT 222.525 322.610 222.695 322.780 ;
        RECT 222.885 322.610 223.055 322.780 ;
        RECT 225.995 322.610 226.165 322.780 ;
        RECT 226.355 322.610 226.525 322.780 ;
        RECT 232.155 322.600 232.325 322.770 ;
        RECT 232.515 322.600 232.685 322.770 ;
        RECT 235.625 322.600 235.795 322.770 ;
        RECT 235.985 322.600 236.155 322.770 ;
        RECT 239.095 322.600 239.265 322.770 ;
        RECT 239.455 322.600 239.625 322.770 ;
        RECT 242.565 322.600 242.735 322.770 ;
        RECT 242.925 322.600 243.095 322.770 ;
        RECT 246.035 322.600 246.205 322.770 ;
        RECT 246.395 322.600 246.565 322.770 ;
        RECT 252.215 322.600 252.385 322.770 ;
        RECT 252.575 322.600 252.745 322.770 ;
        RECT 255.685 322.600 255.855 322.770 ;
        RECT 256.045 322.600 256.215 322.770 ;
        RECT 259.155 322.600 259.325 322.770 ;
        RECT 259.515 322.600 259.685 322.770 ;
        RECT 262.625 322.600 262.795 322.770 ;
        RECT 262.985 322.600 263.155 322.770 ;
        RECT 266.095 322.600 266.265 322.770 ;
        RECT 266.455 322.600 266.625 322.770 ;
        RECT 272.265 322.600 272.435 322.770 ;
        RECT 272.625 322.600 272.795 322.770 ;
        RECT 275.735 322.600 275.905 322.770 ;
        RECT 276.095 322.600 276.265 322.770 ;
        RECT 279.205 322.600 279.375 322.770 ;
        RECT 279.565 322.600 279.735 322.770 ;
        RECT 282.675 322.600 282.845 322.770 ;
        RECT 283.035 322.600 283.205 322.770 ;
        RECT 286.145 322.600 286.315 322.770 ;
        RECT 286.505 322.600 286.675 322.770 ;
        RECT 98.025 321.350 98.195 321.520 ;
        RECT 98.385 321.350 98.555 321.520 ;
        RECT 101.495 321.350 101.665 321.520 ;
        RECT 101.855 321.350 102.025 321.520 ;
        RECT 103.700 320.380 103.870 320.550 ;
        RECT 98.025 318.060 98.195 318.230 ;
        RECT 98.385 318.060 98.555 318.230 ;
        RECT 101.495 318.060 101.665 318.230 ;
        RECT 101.855 318.060 102.025 318.230 ;
        RECT 355.435 322.645 355.605 322.815 ;
        RECT 355.435 322.285 355.605 322.455 ;
        RECT 355.435 321.925 355.605 322.095 ;
        RECT 355.435 321.565 355.605 321.735 ;
        RECT 355.435 321.205 355.605 321.375 ;
        RECT 355.435 320.845 355.605 321.015 ;
        RECT 355.435 320.485 355.605 320.655 ;
        RECT 355.435 320.125 355.605 320.295 ;
        RECT 355.435 319.765 355.605 319.935 ;
        RECT 355.435 319.405 355.605 319.575 ;
        RECT 355.435 319.045 355.605 319.215 ;
        RECT 355.435 318.685 355.605 318.855 ;
        RECT 355.435 318.325 355.605 318.495 ;
        RECT 355.435 317.965 355.605 318.135 ;
        RECT 355.435 317.605 355.605 317.775 ;
        RECT 355.435 317.245 355.605 317.415 ;
        RECT 355.435 316.885 355.605 317.055 ;
        RECT 355.435 316.525 355.605 316.695 ;
        RECT 212.115 316.030 212.285 316.200 ;
        RECT 212.475 316.030 212.645 316.200 ;
        RECT 215.585 316.030 215.755 316.200 ;
        RECT 215.945 316.030 216.115 316.200 ;
        RECT 219.055 316.030 219.225 316.200 ;
        RECT 219.415 316.030 219.585 316.200 ;
        RECT 222.525 316.030 222.695 316.200 ;
        RECT 222.885 316.030 223.055 316.200 ;
        RECT 225.995 316.030 226.165 316.200 ;
        RECT 226.355 316.030 226.525 316.200 ;
        RECT 232.155 316.020 232.325 316.190 ;
        RECT 232.515 316.020 232.685 316.190 ;
        RECT 235.625 316.020 235.795 316.190 ;
        RECT 235.985 316.020 236.155 316.190 ;
        RECT 239.095 316.020 239.265 316.190 ;
        RECT 239.455 316.020 239.625 316.190 ;
        RECT 242.565 316.020 242.735 316.190 ;
        RECT 242.925 316.020 243.095 316.190 ;
        RECT 246.035 316.020 246.205 316.190 ;
        RECT 246.395 316.020 246.565 316.190 ;
        RECT 252.215 316.020 252.385 316.190 ;
        RECT 252.575 316.020 252.745 316.190 ;
        RECT 255.685 316.020 255.855 316.190 ;
        RECT 256.045 316.020 256.215 316.190 ;
        RECT 259.155 316.020 259.325 316.190 ;
        RECT 259.515 316.020 259.685 316.190 ;
        RECT 262.625 316.020 262.795 316.190 ;
        RECT 262.985 316.020 263.155 316.190 ;
        RECT 266.095 316.020 266.265 316.190 ;
        RECT 266.455 316.020 266.625 316.190 ;
        RECT 272.265 316.020 272.435 316.190 ;
        RECT 272.625 316.020 272.795 316.190 ;
        RECT 275.735 316.020 275.905 316.190 ;
        RECT 276.095 316.020 276.265 316.190 ;
        RECT 279.205 316.020 279.375 316.190 ;
        RECT 279.565 316.020 279.735 316.190 ;
        RECT 282.675 316.020 282.845 316.190 ;
        RECT 283.035 316.020 283.205 316.190 ;
        RECT 286.145 316.020 286.315 316.190 ;
        RECT 286.505 316.020 286.675 316.190 ;
        RECT 98.025 314.770 98.195 314.940 ;
        RECT 98.385 314.770 98.555 314.940 ;
        RECT 101.495 314.770 101.665 314.940 ;
        RECT 101.855 314.770 102.025 314.940 ;
        RECT 98.025 311.480 98.195 311.650 ;
        RECT 98.385 311.480 98.555 311.650 ;
        RECT 101.495 311.480 101.665 311.650 ;
        RECT 101.855 311.480 102.025 311.650 ;
        RECT 84.605 307.970 84.775 308.140 ;
        RECT 84.965 307.970 85.135 308.140 ;
        RECT 88.075 307.970 88.245 308.140 ;
        RECT 88.435 307.970 88.605 308.140 ;
        RECT 91.545 307.970 91.715 308.140 ;
        RECT 91.905 307.970 92.075 308.140 ;
        RECT 84.605 304.680 84.775 304.850 ;
        RECT 84.965 304.680 85.135 304.850 ;
        RECT 88.075 304.680 88.245 304.850 ;
        RECT 88.435 304.680 88.605 304.850 ;
        RECT 91.545 304.680 91.715 304.850 ;
        RECT 91.905 304.680 92.075 304.850 ;
        RECT 94.440 304.140 95.330 305.750 ;
        RECT 355.435 316.165 355.605 316.335 ;
        RECT 355.435 315.805 355.605 315.975 ;
        RECT 355.435 315.445 355.605 315.615 ;
        RECT 355.435 315.085 355.605 315.255 ;
        RECT 355.435 314.725 355.605 314.895 ;
        RECT 355.435 314.365 355.605 314.535 ;
        RECT 356.530 327.565 356.700 327.735 ;
        RECT 356.530 327.205 356.700 327.375 ;
        RECT 356.530 324.095 356.700 324.265 ;
        RECT 356.530 323.735 356.700 323.905 ;
        RECT 356.530 320.625 356.700 320.795 ;
        RECT 356.530 320.265 356.700 320.435 ;
        RECT 356.530 317.155 356.700 317.325 ;
        RECT 356.530 316.795 356.700 316.965 ;
        RECT 356.530 313.685 356.700 313.855 ;
        RECT 382.430 332.075 382.600 332.245 ;
        RECT 394.005 345.785 394.175 345.955 ;
        RECT 394.005 345.425 394.175 345.595 ;
        RECT 394.005 345.065 394.175 345.235 ;
        RECT 394.005 344.705 394.175 344.875 ;
        RECT 394.005 344.345 394.175 344.515 ;
        RECT 394.005 343.985 394.175 344.155 ;
        RECT 394.005 343.625 394.175 343.795 ;
        RECT 394.005 343.265 394.175 343.435 ;
        RECT 394.005 342.905 394.175 343.075 ;
        RECT 394.005 342.545 394.175 342.715 ;
        RECT 394.005 342.185 394.175 342.355 ;
        RECT 394.005 341.825 394.175 341.995 ;
        RECT 394.005 341.465 394.175 341.635 ;
        RECT 394.005 341.105 394.175 341.275 ;
        RECT 394.005 340.745 394.175 340.915 ;
        RECT 394.005 340.385 394.175 340.555 ;
        RECT 394.005 340.025 394.175 340.195 ;
        RECT 394.005 339.665 394.175 339.835 ;
        RECT 394.005 339.305 394.175 339.475 ;
        RECT 394.005 338.945 394.175 339.115 ;
        RECT 394.005 338.585 394.175 338.755 ;
        RECT 394.005 338.225 394.175 338.395 ;
        RECT 394.005 337.865 394.175 338.035 ;
        RECT 394.005 337.505 394.175 337.675 ;
        RECT 394.005 337.145 394.175 337.315 ;
        RECT 394.005 336.785 394.175 336.955 ;
        RECT 394.005 336.425 394.175 336.595 ;
        RECT 394.005 336.065 394.175 336.235 ;
        RECT 394.005 335.705 394.175 335.875 ;
        RECT 394.005 335.345 394.175 335.515 ;
        RECT 394.005 334.985 394.175 335.155 ;
        RECT 394.005 334.625 394.175 334.795 ;
        RECT 394.005 334.265 394.175 334.435 ;
        RECT 394.005 333.905 394.175 334.075 ;
        RECT 394.005 333.545 394.175 333.715 ;
        RECT 394.005 333.185 394.175 333.355 ;
        RECT 395.100 346.385 395.270 346.555 ;
        RECT 395.100 346.025 395.270 346.195 ;
        RECT 395.100 342.915 395.270 343.085 ;
        RECT 395.100 342.555 395.270 342.725 ;
        RECT 395.100 339.445 395.270 339.615 ;
        RECT 395.100 339.085 395.270 339.255 ;
        RECT 395.100 335.975 395.270 336.145 ;
        RECT 395.100 335.615 395.270 335.785 ;
        RECT 398.390 346.385 398.560 346.555 ;
        RECT 398.390 346.025 398.560 346.195 ;
        RECT 398.390 342.915 398.560 343.085 ;
        RECT 398.390 342.555 398.560 342.725 ;
        RECT 398.390 339.445 398.560 339.615 ;
        RECT 398.390 339.085 398.560 339.255 ;
        RECT 398.390 335.975 398.560 336.145 ;
        RECT 398.390 335.615 398.560 335.785 ;
        RECT 395.100 332.505 395.270 332.675 ;
        RECT 389.010 332.075 389.180 332.245 ;
        RECT 395.100 332.145 395.270 332.315 ;
        RECT 398.390 332.505 398.560 332.675 ;
        RECT 401.680 346.385 401.850 346.555 ;
        RECT 401.680 346.025 401.850 346.195 ;
        RECT 401.680 342.915 401.850 343.085 ;
        RECT 401.680 342.555 401.850 342.725 ;
        RECT 401.680 339.445 401.850 339.615 ;
        RECT 401.680 339.085 401.850 339.255 ;
        RECT 401.680 335.975 401.850 336.145 ;
        RECT 401.680 335.615 401.850 335.785 ;
        RECT 401.680 332.505 401.850 332.675 ;
        RECT 404.970 346.385 405.140 346.555 ;
        RECT 783.985 346.575 784.155 346.745 ;
        RECT 784.465 346.575 784.635 346.745 ;
        RECT 784.945 346.575 785.115 346.745 ;
        RECT 785.425 346.575 785.595 346.745 ;
        RECT 785.905 346.575 786.075 346.745 ;
        RECT 786.385 346.575 786.555 346.745 ;
        RECT 786.865 346.575 787.035 346.745 ;
        RECT 408.260 346.385 408.430 346.555 ;
        RECT 404.970 346.025 405.140 346.195 ;
        RECT 404.970 342.915 405.140 343.085 ;
        RECT 404.970 342.555 405.140 342.725 ;
        RECT 404.970 339.445 405.140 339.615 ;
        RECT 404.970 339.085 405.140 339.255 ;
        RECT 404.970 335.975 405.140 336.145 ;
        RECT 404.970 335.615 405.140 335.785 ;
        RECT 404.970 332.505 405.140 332.675 ;
        RECT 408.260 346.025 408.430 346.195 ;
        RECT 784.390 346.095 784.560 346.265 ;
        RECT 784.750 346.095 784.920 346.265 ;
        RECT 785.110 346.095 785.280 346.265 ;
        RECT 785.470 346.095 785.640 346.265 ;
        RECT 786.190 346.095 786.360 346.265 ;
        RECT 786.550 346.095 786.720 346.265 ;
        RECT 786.910 346.095 787.080 346.265 ;
        RECT 790.545 346.605 790.715 346.775 ;
        RECT 791.025 346.605 791.195 346.775 ;
        RECT 791.505 346.605 791.675 346.775 ;
        RECT 791.180 346.125 791.350 346.295 ;
        RECT 791.540 346.125 791.710 346.295 ;
        RECT 794.005 346.665 794.175 346.835 ;
        RECT 794.485 346.665 794.655 346.835 ;
        RECT 794.965 346.665 795.135 346.835 ;
        RECT 795.445 346.665 795.615 346.835 ;
        RECT 795.925 346.665 796.095 346.835 ;
        RECT 796.405 346.665 796.575 346.835 ;
        RECT 796.885 346.665 797.055 346.835 ;
        RECT 797.365 346.665 797.535 346.835 ;
        RECT 797.845 346.665 798.015 346.835 ;
        RECT 798.325 346.665 798.495 346.835 ;
        RECT 798.805 346.665 798.975 346.835 ;
        RECT 799.285 346.665 799.455 346.835 ;
        RECT 799.765 346.665 799.935 346.835 ;
        RECT 800.245 346.665 800.415 346.835 ;
        RECT 800.725 346.665 800.895 346.835 ;
        RECT 801.205 346.665 801.375 346.835 ;
        RECT 801.685 346.665 801.855 346.835 ;
        RECT 802.165 346.665 802.335 346.835 ;
        RECT 802.645 346.665 802.815 346.835 ;
        RECT 803.125 346.665 803.295 346.835 ;
        RECT 803.605 346.665 803.775 346.835 ;
        RECT 804.085 346.665 804.255 346.835 ;
        RECT 804.565 346.665 804.735 346.835 ;
        RECT 805.045 346.665 805.215 346.835 ;
        RECT 805.525 346.665 805.695 346.835 ;
        RECT 806.005 346.665 806.175 346.835 ;
        RECT 806.485 346.665 806.655 346.835 ;
        RECT 806.965 346.665 807.135 346.835 ;
        RECT 807.445 346.665 807.615 346.835 ;
        RECT 807.925 346.665 808.095 346.835 ;
        RECT 808.405 346.665 808.575 346.835 ;
        RECT 808.885 346.665 809.055 346.835 ;
        RECT 794.520 346.185 794.690 346.355 ;
        RECT 794.880 346.185 795.050 346.355 ;
        RECT 795.240 346.185 795.410 346.355 ;
        RECT 796.050 346.185 796.220 346.355 ;
        RECT 796.410 346.185 796.580 346.355 ;
        RECT 796.770 346.185 796.940 346.355 ;
        RECT 797.805 346.185 797.975 346.355 ;
        RECT 798.165 346.185 798.335 346.355 ;
        RECT 798.525 346.185 798.695 346.355 ;
        RECT 800.500 346.185 800.670 346.355 ;
        RECT 800.860 346.185 801.030 346.355 ;
        RECT 801.220 346.185 801.390 346.355 ;
        RECT 802.840 346.185 803.010 346.355 ;
        RECT 803.200 346.185 803.370 346.355 ;
        RECT 803.560 346.185 803.730 346.355 ;
        RECT 805.990 346.185 806.160 346.355 ;
        RECT 808.020 346.185 808.190 346.355 ;
        RECT 808.380 346.185 808.550 346.355 ;
        RECT 813.365 346.575 813.535 346.745 ;
        RECT 813.845 346.575 814.015 346.745 ;
        RECT 814.325 346.575 814.495 346.745 ;
        RECT 814.805 346.575 814.975 346.745 ;
        RECT 815.285 346.575 815.455 346.745 ;
        RECT 815.765 346.575 815.935 346.745 ;
        RECT 816.245 346.575 816.415 346.745 ;
        RECT 816.725 346.575 816.895 346.745 ;
        RECT 817.205 346.575 817.375 346.745 ;
        RECT 817.685 346.575 817.855 346.745 ;
        RECT 818.165 346.575 818.335 346.745 ;
        RECT 818.645 346.575 818.815 346.745 ;
        RECT 819.125 346.575 819.295 346.745 ;
        RECT 819.605 346.575 819.775 346.745 ;
        RECT 820.085 346.575 820.255 346.745 ;
        RECT 820.565 346.575 820.735 346.745 ;
        RECT 821.045 346.575 821.215 346.745 ;
        RECT 821.525 346.575 821.695 346.745 ;
        RECT 822.005 346.575 822.175 346.745 ;
        RECT 822.485 346.575 822.655 346.745 ;
        RECT 822.965 346.575 823.135 346.745 ;
        RECT 823.445 346.575 823.615 346.745 ;
        RECT 823.925 346.575 824.095 346.745 ;
        RECT 824.405 346.575 824.575 346.745 ;
        RECT 824.885 346.575 825.055 346.745 ;
        RECT 825.365 346.575 825.535 346.745 ;
        RECT 825.845 346.575 826.015 346.745 ;
        RECT 826.325 346.575 826.495 346.745 ;
        RECT 826.805 346.575 826.975 346.745 ;
        RECT 827.285 346.575 827.455 346.745 ;
        RECT 827.765 346.575 827.935 346.745 ;
        RECT 828.245 346.575 828.415 346.745 ;
        RECT 813.880 346.095 814.050 346.265 ;
        RECT 814.240 346.095 814.410 346.265 ;
        RECT 814.600 346.095 814.770 346.265 ;
        RECT 815.410 346.095 815.580 346.265 ;
        RECT 815.770 346.095 815.940 346.265 ;
        RECT 816.130 346.095 816.300 346.265 ;
        RECT 817.165 346.095 817.335 346.265 ;
        RECT 817.525 346.095 817.695 346.265 ;
        RECT 817.885 346.095 818.055 346.265 ;
        RECT 819.860 346.095 820.030 346.265 ;
        RECT 820.220 346.095 820.390 346.265 ;
        RECT 820.580 346.095 820.750 346.265 ;
        RECT 822.200 346.095 822.370 346.265 ;
        RECT 822.560 346.095 822.730 346.265 ;
        RECT 822.920 346.095 823.090 346.265 ;
        RECT 825.350 346.095 825.520 346.265 ;
        RECT 827.380 346.095 827.550 346.265 ;
        RECT 827.740 346.095 827.910 346.265 ;
        RECT 408.260 342.915 408.430 343.085 ;
        RECT 408.260 342.555 408.430 342.725 ;
        RECT 408.260 339.445 408.430 339.615 ;
        RECT 408.260 339.085 408.430 339.255 ;
        RECT 408.260 335.975 408.430 336.145 ;
        RECT 408.260 335.615 408.430 335.785 ;
        RECT 398.390 332.145 398.560 332.315 ;
        RECT 401.680 332.145 401.850 332.315 ;
        RECT 404.970 332.145 405.140 332.315 ;
        RECT 408.260 332.505 408.430 332.675 ;
        RECT 408.260 332.145 408.430 332.315 ;
        RECT 601.450 332.165 601.620 332.335 ;
        RECT 602.630 332.175 602.800 332.345 ;
        RECT 604.210 332.175 604.380 332.345 ;
        RECT 605.790 332.175 605.960 332.345 ;
        RECT 607.150 332.185 607.320 332.355 ;
        RECT 608.730 332.185 608.900 332.355 ;
        RECT 610.310 332.185 610.480 332.355 ;
        RECT 611.670 332.185 611.840 332.355 ;
        RECT 613.250 332.185 613.420 332.355 ;
        RECT 614.830 332.185 615.000 332.355 ;
        RECT 616.100 332.165 616.270 332.335 ;
        RECT 617.680 332.165 617.850 332.335 ;
        RECT 619.260 332.165 619.430 332.335 ;
        RECT 620.480 332.175 620.650 332.345 ;
        RECT 622.060 332.175 622.230 332.345 ;
        RECT 623.640 332.175 623.810 332.345 ;
        RECT 624.800 332.165 624.970 332.335 ;
        RECT 626.380 332.165 626.550 332.335 ;
        RECT 627.960 332.165 628.130 332.335 ;
        RECT 629.180 332.395 629.350 332.565 ;
        RECT 663.345 332.485 663.515 332.655 ;
        RECT 663.825 332.485 663.995 332.655 ;
        RECT 664.305 332.485 664.475 332.655 ;
        RECT 664.785 332.485 664.955 332.655 ;
        RECT 665.265 332.485 665.435 332.655 ;
        RECT 665.745 332.485 665.915 332.655 ;
        RECT 666.225 332.485 666.395 332.655 ;
        RECT 668.975 332.485 669.145 332.655 ;
        RECT 669.455 332.485 669.625 332.655 ;
        RECT 669.935 332.485 670.105 332.655 ;
        RECT 670.415 332.485 670.585 332.655 ;
        RECT 670.895 332.485 671.065 332.655 ;
        RECT 671.375 332.485 671.545 332.655 ;
        RECT 671.855 332.485 672.025 332.655 ;
        RECT 674.735 332.385 674.905 332.555 ;
        RECT 675.215 332.385 675.385 332.555 ;
        RECT 675.695 332.385 675.865 332.555 ;
        RECT 676.175 332.385 676.345 332.555 ;
        RECT 676.655 332.385 676.825 332.555 ;
        RECT 677.135 332.385 677.305 332.555 ;
        RECT 677.615 332.385 677.785 332.555 ;
        RECT 681.765 332.425 681.935 332.595 ;
        RECT 682.245 332.425 682.415 332.595 ;
        RECT 682.725 332.425 682.895 332.595 ;
        RECT 683.205 332.425 683.375 332.595 ;
        RECT 683.685 332.425 683.855 332.595 ;
        RECT 684.165 332.425 684.335 332.595 ;
        RECT 684.645 332.425 684.815 332.595 ;
        RECT 685.125 332.425 685.295 332.595 ;
        RECT 687.625 332.435 687.795 332.605 ;
        RECT 688.105 332.435 688.275 332.605 ;
        RECT 688.585 332.435 688.755 332.605 ;
        RECT 689.065 332.435 689.235 332.605 ;
        RECT 689.545 332.435 689.715 332.605 ;
        RECT 690.025 332.435 690.195 332.605 ;
        RECT 690.505 332.435 690.675 332.605 ;
        RECT 601.450 331.805 601.620 331.975 ;
        RECT 601.450 331.445 601.620 331.615 ;
        RECT 601.450 331.085 601.620 331.255 ;
        RECT 629.180 332.035 629.350 332.205 ;
        RECT 629.180 331.675 629.350 331.845 ;
        RECT 629.180 331.315 629.350 331.485 ;
        RECT 663.300 332.005 663.470 332.175 ;
        RECT 663.660 332.005 663.830 332.175 ;
        RECT 664.020 332.005 664.190 332.175 ;
        RECT 635.415 331.145 635.585 331.315 ;
        RECT 635.895 331.145 636.065 331.315 ;
        RECT 636.375 331.145 636.545 331.315 ;
        RECT 639.605 331.235 639.775 331.405 ;
        RECT 640.085 331.235 640.255 331.405 ;
        RECT 640.565 331.235 640.735 331.405 ;
        RECT 643.705 331.215 643.875 331.385 ;
        RECT 644.185 331.215 644.355 331.385 ;
        RECT 644.665 331.215 644.835 331.385 ;
        RECT 595.525 330.695 595.695 330.865 ;
        RECT 596.005 330.695 596.175 330.865 ;
        RECT 596.485 330.695 596.655 330.865 ;
        RECT 601.450 330.725 601.620 330.895 ;
        RECT 596.160 330.215 596.330 330.385 ;
        RECT 596.520 330.215 596.690 330.385 ;
        RECT 602.630 330.705 602.800 330.875 ;
        RECT 604.210 330.705 604.380 330.875 ;
        RECT 605.790 330.705 605.960 330.875 ;
        RECT 607.150 330.715 607.320 330.885 ;
        RECT 608.730 330.715 608.900 330.885 ;
        RECT 610.310 330.715 610.480 330.885 ;
        RECT 611.670 330.715 611.840 330.885 ;
        RECT 613.250 330.715 613.420 330.885 ;
        RECT 614.830 330.715 615.000 330.885 ;
        RECT 616.100 330.695 616.270 330.865 ;
        RECT 617.680 330.695 617.850 330.865 ;
        RECT 619.260 330.695 619.430 330.865 ;
        RECT 620.480 330.705 620.650 330.875 ;
        RECT 622.060 330.705 622.230 330.875 ;
        RECT 623.640 330.705 623.810 330.875 ;
        RECT 624.800 330.695 624.970 330.865 ;
        RECT 626.380 330.695 626.550 330.865 ;
        RECT 627.960 330.695 628.130 330.865 ;
        RECT 629.180 330.955 629.350 331.125 ;
        RECT 629.180 330.595 629.350 330.765 ;
        RECT 635.380 330.665 635.550 330.835 ;
        RECT 635.740 330.665 635.910 330.835 ;
        RECT 639.570 330.755 639.740 330.925 ;
        RECT 639.930 330.755 640.100 330.925 ;
        RECT 643.670 330.735 643.840 330.905 ;
        RECT 644.030 330.735 644.200 330.905 ;
        RECT 664.740 332.005 664.910 332.175 ;
        RECT 665.100 332.005 665.270 332.175 ;
        RECT 665.460 332.005 665.630 332.175 ;
        RECT 665.820 332.005 665.990 332.175 ;
        RECT 668.930 332.005 669.100 332.175 ;
        RECT 669.290 332.005 669.460 332.175 ;
        RECT 669.650 332.005 669.820 332.175 ;
        RECT 670.370 332.005 670.540 332.175 ;
        RECT 670.730 332.005 670.900 332.175 ;
        RECT 671.090 332.005 671.260 332.175 ;
        RECT 671.450 332.005 671.620 332.175 ;
        RECT 675.410 331.905 675.580 332.075 ;
        RECT 675.770 331.905 675.940 332.075 ;
        RECT 676.130 331.905 676.300 332.075 ;
        RECT 676.490 331.905 676.660 332.075 ;
        RECT 676.850 331.905 677.020 332.075 ;
        RECT 677.210 331.905 677.380 332.075 ;
        RECT 682.200 331.945 682.370 332.115 ;
        RECT 682.560 331.945 682.730 332.115 ;
        RECT 682.920 331.945 683.090 332.115 ;
        RECT 683.840 331.945 684.010 332.115 ;
        RECT 684.200 331.945 684.370 332.115 ;
        RECT 684.560 331.945 684.730 332.115 ;
        RECT 687.580 331.955 687.750 332.125 ;
        RECT 687.940 331.955 688.110 332.125 ;
        RECT 688.300 331.955 688.470 332.125 ;
        RECT 689.020 331.955 689.190 332.125 ;
        RECT 689.380 331.955 689.550 332.125 ;
        RECT 689.740 331.955 689.910 332.125 ;
        RECT 690.100 331.955 690.270 332.125 ;
        RECT 862.550 329.310 863.440 330.920 ;
        RECT 359.820 327.565 359.990 327.735 ;
        RECT 359.820 327.205 359.990 327.375 ;
        RECT 359.820 324.095 359.990 324.265 ;
        RECT 359.820 323.735 359.990 323.905 ;
        RECT 359.820 320.625 359.990 320.795 ;
        RECT 359.820 320.265 359.990 320.435 ;
        RECT 359.820 317.155 359.990 317.325 ;
        RECT 359.820 316.795 359.990 316.965 ;
        RECT 356.530 313.325 356.700 313.495 ;
        RECT 359.820 313.685 359.990 313.855 ;
        RECT 363.110 327.565 363.280 327.735 ;
        RECT 363.110 327.205 363.280 327.375 ;
        RECT 363.110 324.095 363.280 324.265 ;
        RECT 363.110 323.735 363.280 323.905 ;
        RECT 363.110 320.625 363.280 320.795 ;
        RECT 363.110 320.265 363.280 320.435 ;
        RECT 363.110 317.155 363.280 317.325 ;
        RECT 363.110 316.795 363.280 316.965 ;
        RECT 363.110 313.685 363.280 313.855 ;
        RECT 366.400 327.565 366.570 327.735 ;
        RECT 369.690 327.565 369.860 327.735 ;
        RECT 366.400 327.205 366.570 327.375 ;
        RECT 366.400 324.095 366.570 324.265 ;
        RECT 366.400 323.735 366.570 323.905 ;
        RECT 366.400 320.625 366.570 320.795 ;
        RECT 366.400 320.265 366.570 320.435 ;
        RECT 366.400 317.155 366.570 317.325 ;
        RECT 366.400 316.795 366.570 316.965 ;
        RECT 366.400 313.685 366.570 313.855 ;
        RECT 369.690 327.205 369.860 327.375 ;
        RECT 369.690 324.095 369.860 324.265 ;
        RECT 369.690 323.735 369.860 323.905 ;
        RECT 369.690 320.625 369.860 320.795 ;
        RECT 369.690 320.265 369.860 320.435 ;
        RECT 369.690 317.155 369.860 317.325 ;
        RECT 369.690 316.795 369.860 316.965 ;
        RECT 359.820 313.325 359.990 313.495 ;
        RECT 363.110 313.325 363.280 313.495 ;
        RECT 366.400 313.325 366.570 313.495 ;
        RECT 369.690 313.685 369.860 313.855 ;
        RECT 374.755 326.865 374.925 327.035 ;
        RECT 374.755 326.505 374.925 326.675 ;
        RECT 374.755 326.145 374.925 326.315 ;
        RECT 374.755 325.785 374.925 325.955 ;
        RECT 374.755 325.425 374.925 325.595 ;
        RECT 374.755 325.065 374.925 325.235 ;
        RECT 374.755 324.705 374.925 324.875 ;
        RECT 374.755 324.345 374.925 324.515 ;
        RECT 374.755 323.985 374.925 324.155 ;
        RECT 374.755 323.625 374.925 323.795 ;
        RECT 374.755 323.265 374.925 323.435 ;
        RECT 374.755 322.905 374.925 323.075 ;
        RECT 374.755 322.545 374.925 322.715 ;
        RECT 374.755 322.185 374.925 322.355 ;
        RECT 374.755 321.825 374.925 321.995 ;
        RECT 374.755 321.465 374.925 321.635 ;
        RECT 374.755 321.105 374.925 321.275 ;
        RECT 374.755 320.745 374.925 320.915 ;
        RECT 374.755 320.385 374.925 320.555 ;
        RECT 374.755 320.025 374.925 320.195 ;
        RECT 374.755 319.665 374.925 319.835 ;
        RECT 374.755 319.305 374.925 319.475 ;
        RECT 374.755 318.945 374.925 319.115 ;
        RECT 374.755 318.585 374.925 318.755 ;
        RECT 374.755 318.225 374.925 318.395 ;
        RECT 374.755 317.865 374.925 318.035 ;
        RECT 374.755 317.505 374.925 317.675 ;
        RECT 374.755 317.145 374.925 317.315 ;
        RECT 374.755 316.785 374.925 316.955 ;
        RECT 374.755 316.425 374.925 316.595 ;
        RECT 374.755 316.065 374.925 316.235 ;
        RECT 374.755 315.705 374.925 315.875 ;
        RECT 374.755 315.345 374.925 315.515 ;
        RECT 374.755 314.985 374.925 315.155 ;
        RECT 374.755 314.625 374.925 314.795 ;
        RECT 374.755 314.265 374.925 314.435 ;
        RECT 375.850 327.465 376.020 327.635 ;
        RECT 375.850 327.105 376.020 327.275 ;
        RECT 375.850 323.995 376.020 324.165 ;
        RECT 375.850 323.635 376.020 323.805 ;
        RECT 375.850 320.525 376.020 320.695 ;
        RECT 375.850 320.165 376.020 320.335 ;
        RECT 375.850 317.055 376.020 317.225 ;
        RECT 375.850 316.695 376.020 316.865 ;
        RECT 375.850 313.585 376.020 313.755 ;
        RECT 369.690 313.325 369.860 313.495 ;
        RECT 382.430 327.465 382.600 327.635 ;
        RECT 389.010 327.465 389.180 327.635 ;
        RECT 382.430 327.105 382.600 327.275 ;
        RECT 382.430 323.995 382.600 324.165 ;
        RECT 382.430 323.635 382.600 323.805 ;
        RECT 382.430 320.525 382.600 320.695 ;
        RECT 382.430 320.165 382.600 320.335 ;
        RECT 382.430 317.055 382.600 317.225 ;
        RECT 382.430 316.695 382.600 316.865 ;
        RECT 382.430 313.585 382.600 313.755 ;
        RECT 389.010 327.105 389.180 327.275 ;
        RECT 389.010 323.995 389.180 324.165 ;
        RECT 389.010 323.635 389.180 323.805 ;
        RECT 389.010 320.525 389.180 320.695 ;
        RECT 389.010 320.165 389.180 320.335 ;
        RECT 389.010 317.055 389.180 317.225 ;
        RECT 389.010 316.695 389.180 316.865 ;
        RECT 389.010 313.585 389.180 313.755 ;
        RECT 375.850 313.225 376.020 313.395 ;
        RECT 212.115 309.450 212.285 309.620 ;
        RECT 212.475 309.450 212.645 309.620 ;
        RECT 215.585 309.450 215.755 309.620 ;
        RECT 215.945 309.450 216.115 309.620 ;
        RECT 219.055 309.450 219.225 309.620 ;
        RECT 219.415 309.450 219.585 309.620 ;
        RECT 222.525 309.450 222.695 309.620 ;
        RECT 222.885 309.450 223.055 309.620 ;
        RECT 225.995 309.450 226.165 309.620 ;
        RECT 226.355 309.450 226.525 309.620 ;
        RECT 232.155 309.440 232.325 309.610 ;
        RECT 232.515 309.440 232.685 309.610 ;
        RECT 235.625 309.440 235.795 309.610 ;
        RECT 235.985 309.440 236.155 309.610 ;
        RECT 239.095 309.440 239.265 309.610 ;
        RECT 239.455 309.440 239.625 309.610 ;
        RECT 242.565 309.440 242.735 309.610 ;
        RECT 242.925 309.440 243.095 309.610 ;
        RECT 246.035 309.440 246.205 309.610 ;
        RECT 246.395 309.440 246.565 309.610 ;
        RECT 252.215 309.440 252.385 309.610 ;
        RECT 252.575 309.440 252.745 309.610 ;
        RECT 255.685 309.440 255.855 309.610 ;
        RECT 256.045 309.440 256.215 309.610 ;
        RECT 259.155 309.440 259.325 309.610 ;
        RECT 259.515 309.440 259.685 309.610 ;
        RECT 262.625 309.440 262.795 309.610 ;
        RECT 262.985 309.440 263.155 309.610 ;
        RECT 266.095 309.440 266.265 309.610 ;
        RECT 266.455 309.440 266.625 309.610 ;
        RECT 272.265 309.440 272.435 309.610 ;
        RECT 272.625 309.440 272.795 309.610 ;
        RECT 275.735 309.440 275.905 309.610 ;
        RECT 276.095 309.440 276.265 309.610 ;
        RECT 279.205 309.440 279.375 309.610 ;
        RECT 279.565 309.440 279.735 309.610 ;
        RECT 282.675 309.440 282.845 309.610 ;
        RECT 283.035 309.440 283.205 309.610 ;
        RECT 286.145 309.440 286.315 309.610 ;
        RECT 286.505 309.440 286.675 309.610 ;
        RECT 98.025 308.190 98.195 308.360 ;
        RECT 98.385 308.190 98.555 308.360 ;
        RECT 101.495 308.190 101.665 308.360 ;
        RECT 101.855 308.190 102.025 308.360 ;
        RECT 98.025 304.900 98.195 305.070 ;
        RECT 98.385 304.900 98.555 305.070 ;
        RECT 101.495 304.900 101.665 305.070 ;
        RECT 101.855 304.900 102.025 305.070 ;
        RECT 215.250 303.100 225.860 303.990 ;
        RECT 235.220 303.100 245.830 303.990 ;
        RECT 255.330 303.100 265.940 303.990 ;
        RECT 275.440 303.100 286.050 303.990 ;
        RECT 98.025 301.610 98.195 301.780 ;
        RECT 98.385 301.610 98.555 301.780 ;
        RECT 101.495 301.610 101.665 301.780 ;
        RECT 101.855 301.610 102.025 301.780 ;
        RECT 212.075 301.620 212.245 301.790 ;
        RECT 212.435 301.620 212.605 301.790 ;
        RECT 215.545 301.620 215.715 301.790 ;
        RECT 215.905 301.620 216.075 301.790 ;
        RECT 219.015 301.620 219.185 301.790 ;
        RECT 219.375 301.620 219.545 301.790 ;
        RECT 222.485 301.620 222.655 301.790 ;
        RECT 222.845 301.620 223.015 301.790 ;
        RECT 225.955 301.620 226.125 301.790 ;
        RECT 226.315 301.620 226.485 301.790 ;
        RECT 232.045 301.620 232.215 301.790 ;
        RECT 232.405 301.620 232.575 301.790 ;
        RECT 235.515 301.620 235.685 301.790 ;
        RECT 235.875 301.620 236.045 301.790 ;
        RECT 238.985 301.620 239.155 301.790 ;
        RECT 239.345 301.620 239.515 301.790 ;
        RECT 242.455 301.620 242.625 301.790 ;
        RECT 242.815 301.620 242.985 301.790 ;
        RECT 245.925 301.620 246.095 301.790 ;
        RECT 246.285 301.620 246.455 301.790 ;
        RECT 252.155 301.620 252.325 301.790 ;
        RECT 252.515 301.620 252.685 301.790 ;
        RECT 255.625 301.620 255.795 301.790 ;
        RECT 255.985 301.620 256.155 301.790 ;
        RECT 259.095 301.620 259.265 301.790 ;
        RECT 259.455 301.620 259.625 301.790 ;
        RECT 262.565 301.620 262.735 301.790 ;
        RECT 262.925 301.620 263.095 301.790 ;
        RECT 266.035 301.620 266.205 301.790 ;
        RECT 266.395 301.620 266.565 301.790 ;
        RECT 272.265 301.620 272.435 301.790 ;
        RECT 272.625 301.620 272.795 301.790 ;
        RECT 275.735 301.620 275.905 301.790 ;
        RECT 276.095 301.620 276.265 301.790 ;
        RECT 279.205 301.620 279.375 301.790 ;
        RECT 279.565 301.620 279.735 301.790 ;
        RECT 282.675 301.620 282.845 301.790 ;
        RECT 283.035 301.620 283.205 301.790 ;
        RECT 286.145 301.620 286.315 301.790 ;
        RECT 286.505 301.620 286.675 301.790 ;
        RECT 4.995 301.360 5.165 301.530 ;
        RECT 5.355 301.360 5.525 301.530 ;
        RECT 8.465 301.360 8.635 301.530 ;
        RECT 8.825 301.360 8.995 301.530 ;
        RECT 11.935 301.360 12.105 301.530 ;
        RECT 12.295 301.360 12.465 301.530 ;
        RECT 18.335 301.340 18.505 301.510 ;
        RECT 18.695 301.340 18.865 301.510 ;
        RECT 21.805 301.340 21.975 301.510 ;
        RECT 22.165 301.340 22.335 301.510 ;
        RECT 25.275 301.340 25.445 301.510 ;
        RECT 25.635 301.340 25.805 301.510 ;
        RECT 31.705 301.370 31.875 301.540 ;
        RECT 32.065 301.370 32.235 301.540 ;
        RECT 35.175 301.370 35.345 301.540 ;
        RECT 35.535 301.370 35.705 301.540 ;
        RECT 38.645 301.370 38.815 301.540 ;
        RECT 39.005 301.370 39.175 301.540 ;
        RECT 44.935 301.370 45.105 301.540 ;
        RECT 45.295 301.370 45.465 301.540 ;
        RECT 48.405 301.370 48.575 301.540 ;
        RECT 48.765 301.370 48.935 301.540 ;
        RECT 51.875 301.370 52.045 301.540 ;
        RECT 52.235 301.370 52.405 301.540 ;
        RECT 58.205 301.340 58.375 301.510 ;
        RECT 58.565 301.340 58.735 301.510 ;
        RECT 61.675 301.340 61.845 301.510 ;
        RECT 62.035 301.340 62.205 301.510 ;
        RECT 65.145 301.340 65.315 301.510 ;
        RECT 65.505 301.340 65.675 301.510 ;
        RECT 71.475 301.370 71.645 301.540 ;
        RECT 71.835 301.370 72.005 301.540 ;
        RECT 74.945 301.370 75.115 301.540 ;
        RECT 75.305 301.370 75.475 301.540 ;
        RECT 78.415 301.370 78.585 301.540 ;
        RECT 78.775 301.370 78.945 301.540 ;
        RECT 84.605 301.390 84.775 301.560 ;
        RECT 84.965 301.390 85.135 301.560 ;
        RECT 88.075 301.390 88.245 301.560 ;
        RECT 88.435 301.390 88.605 301.560 ;
        RECT 91.545 301.390 91.715 301.560 ;
        RECT 91.905 301.390 92.075 301.560 ;
        RECT 355.435 308.145 355.605 308.315 ;
        RECT 355.435 307.785 355.605 307.955 ;
        RECT 355.435 307.425 355.605 307.595 ;
        RECT 355.435 307.065 355.605 307.235 ;
        RECT 355.435 306.705 355.605 306.875 ;
        RECT 355.435 306.345 355.605 306.515 ;
        RECT 355.435 305.985 355.605 306.155 ;
        RECT 355.435 305.625 355.605 305.795 ;
        RECT 355.435 305.265 355.605 305.435 ;
        RECT 355.435 304.905 355.605 305.075 ;
        RECT 355.435 304.545 355.605 304.715 ;
        RECT 355.435 304.185 355.605 304.355 ;
        RECT 355.435 303.825 355.605 303.995 ;
        RECT 355.435 303.465 355.605 303.635 ;
        RECT 355.435 303.105 355.605 303.275 ;
        RECT 355.435 302.745 355.605 302.915 ;
        RECT 355.435 302.385 355.605 302.555 ;
        RECT 355.435 302.025 355.605 302.195 ;
        RECT 355.435 301.665 355.605 301.835 ;
        RECT 5.295 297.920 5.465 298.090 ;
        RECT 5.655 297.920 5.825 298.090 ;
        RECT 6.015 297.920 6.185 298.090 ;
        RECT 6.375 297.920 6.545 298.090 ;
        RECT 6.735 297.920 6.905 298.090 ;
        RECT 7.095 297.920 7.265 298.090 ;
        RECT 7.455 297.920 7.625 298.090 ;
        RECT 7.815 297.920 7.985 298.090 ;
        RECT 8.175 297.920 8.345 298.090 ;
        RECT 8.535 297.920 8.705 298.090 ;
        RECT 8.895 297.920 9.065 298.090 ;
        RECT 9.255 297.920 9.425 298.090 ;
        RECT 9.615 297.920 9.785 298.090 ;
        RECT 9.975 297.920 10.145 298.090 ;
        RECT 10.335 297.920 10.505 298.090 ;
        RECT 10.695 297.920 10.865 298.090 ;
        RECT 11.055 297.920 11.225 298.090 ;
        RECT 11.415 297.920 11.585 298.090 ;
        RECT 11.775 297.920 11.945 298.090 ;
        RECT 12.135 297.920 12.305 298.090 ;
        RECT 18.635 297.900 18.805 298.070 ;
        RECT 18.995 297.900 19.165 298.070 ;
        RECT 19.355 297.900 19.525 298.070 ;
        RECT 19.715 297.900 19.885 298.070 ;
        RECT 20.075 297.900 20.245 298.070 ;
        RECT 20.435 297.900 20.605 298.070 ;
        RECT 20.795 297.900 20.965 298.070 ;
        RECT 21.155 297.900 21.325 298.070 ;
        RECT 21.515 297.900 21.685 298.070 ;
        RECT 21.875 297.900 22.045 298.070 ;
        RECT 22.235 297.900 22.405 298.070 ;
        RECT 22.595 297.900 22.765 298.070 ;
        RECT 22.955 297.900 23.125 298.070 ;
        RECT 23.315 297.900 23.485 298.070 ;
        RECT 23.675 297.900 23.845 298.070 ;
        RECT 24.035 297.900 24.205 298.070 ;
        RECT 24.395 297.900 24.565 298.070 ;
        RECT 24.755 297.900 24.925 298.070 ;
        RECT 25.115 297.900 25.285 298.070 ;
        RECT 25.475 297.900 25.645 298.070 ;
        RECT 32.005 297.930 32.175 298.100 ;
        RECT 32.365 297.930 32.535 298.100 ;
        RECT 32.725 297.930 32.895 298.100 ;
        RECT 33.085 297.930 33.255 298.100 ;
        RECT 33.445 297.930 33.615 298.100 ;
        RECT 33.805 297.930 33.975 298.100 ;
        RECT 34.165 297.930 34.335 298.100 ;
        RECT 34.525 297.930 34.695 298.100 ;
        RECT 34.885 297.930 35.055 298.100 ;
        RECT 35.245 297.930 35.415 298.100 ;
        RECT 35.605 297.930 35.775 298.100 ;
        RECT 35.965 297.930 36.135 298.100 ;
        RECT 36.325 297.930 36.495 298.100 ;
        RECT 36.685 297.930 36.855 298.100 ;
        RECT 37.045 297.930 37.215 298.100 ;
        RECT 37.405 297.930 37.575 298.100 ;
        RECT 37.765 297.930 37.935 298.100 ;
        RECT 38.125 297.930 38.295 298.100 ;
        RECT 38.485 297.930 38.655 298.100 ;
        RECT 38.845 297.930 39.015 298.100 ;
        RECT 45.235 297.930 45.405 298.100 ;
        RECT 45.595 297.930 45.765 298.100 ;
        RECT 45.955 297.930 46.125 298.100 ;
        RECT 46.315 297.930 46.485 298.100 ;
        RECT 46.675 297.930 46.845 298.100 ;
        RECT 47.035 297.930 47.205 298.100 ;
        RECT 47.395 297.930 47.565 298.100 ;
        RECT 47.755 297.930 47.925 298.100 ;
        RECT 48.115 297.930 48.285 298.100 ;
        RECT 48.475 297.930 48.645 298.100 ;
        RECT 48.835 297.930 49.005 298.100 ;
        RECT 49.195 297.930 49.365 298.100 ;
        RECT 49.555 297.930 49.725 298.100 ;
        RECT 49.915 297.930 50.085 298.100 ;
        RECT 50.275 297.930 50.445 298.100 ;
        RECT 50.635 297.930 50.805 298.100 ;
        RECT 50.995 297.930 51.165 298.100 ;
        RECT 51.355 297.930 51.525 298.100 ;
        RECT 51.715 297.930 51.885 298.100 ;
        RECT 52.075 297.930 52.245 298.100 ;
        RECT 58.505 297.900 58.675 298.070 ;
        RECT 58.865 297.900 59.035 298.070 ;
        RECT 59.225 297.900 59.395 298.070 ;
        RECT 59.585 297.900 59.755 298.070 ;
        RECT 59.945 297.900 60.115 298.070 ;
        RECT 60.305 297.900 60.475 298.070 ;
        RECT 60.665 297.900 60.835 298.070 ;
        RECT 61.025 297.900 61.195 298.070 ;
        RECT 61.385 297.900 61.555 298.070 ;
        RECT 61.745 297.900 61.915 298.070 ;
        RECT 62.105 297.900 62.275 298.070 ;
        RECT 62.465 297.900 62.635 298.070 ;
        RECT 62.825 297.900 62.995 298.070 ;
        RECT 63.185 297.900 63.355 298.070 ;
        RECT 63.545 297.900 63.715 298.070 ;
        RECT 63.905 297.900 64.075 298.070 ;
        RECT 64.265 297.900 64.435 298.070 ;
        RECT 64.625 297.900 64.795 298.070 ;
        RECT 64.985 297.900 65.155 298.070 ;
        RECT 65.345 297.900 65.515 298.070 ;
        RECT 71.775 297.930 71.945 298.100 ;
        RECT 72.135 297.930 72.305 298.100 ;
        RECT 72.495 297.930 72.665 298.100 ;
        RECT 72.855 297.930 73.025 298.100 ;
        RECT 73.215 297.930 73.385 298.100 ;
        RECT 73.575 297.930 73.745 298.100 ;
        RECT 73.935 297.930 74.105 298.100 ;
        RECT 74.295 297.930 74.465 298.100 ;
        RECT 74.655 297.930 74.825 298.100 ;
        RECT 75.015 297.930 75.185 298.100 ;
        RECT 75.375 297.930 75.545 298.100 ;
        RECT 75.735 297.930 75.905 298.100 ;
        RECT 76.095 297.930 76.265 298.100 ;
        RECT 76.455 297.930 76.625 298.100 ;
        RECT 76.815 297.930 76.985 298.100 ;
        RECT 77.175 297.930 77.345 298.100 ;
        RECT 77.535 297.930 77.705 298.100 ;
        RECT 77.895 297.930 78.065 298.100 ;
        RECT 78.255 297.930 78.425 298.100 ;
        RECT 78.615 297.930 78.785 298.100 ;
        RECT 84.905 297.950 85.075 298.120 ;
        RECT 85.265 297.950 85.435 298.120 ;
        RECT 85.625 297.950 85.795 298.120 ;
        RECT 85.985 297.950 86.155 298.120 ;
        RECT 86.345 297.950 86.515 298.120 ;
        RECT 86.705 297.950 86.875 298.120 ;
        RECT 87.065 297.950 87.235 298.120 ;
        RECT 87.425 297.950 87.595 298.120 ;
        RECT 87.785 297.950 87.955 298.120 ;
        RECT 88.145 297.950 88.315 298.120 ;
        RECT 88.505 297.950 88.675 298.120 ;
        RECT 88.865 297.950 89.035 298.120 ;
        RECT 89.225 297.950 89.395 298.120 ;
        RECT 89.585 297.950 89.755 298.120 ;
        RECT 89.945 297.950 90.115 298.120 ;
        RECT 90.305 297.950 90.475 298.120 ;
        RECT 90.665 297.950 90.835 298.120 ;
        RECT 91.025 297.950 91.195 298.120 ;
        RECT 91.385 297.950 91.555 298.120 ;
        RECT 91.745 297.950 91.915 298.120 ;
        RECT 97.820 297.745 102.310 298.275 ;
        RECT 355.435 301.305 355.605 301.475 ;
        RECT 355.435 300.945 355.605 301.115 ;
        RECT 355.435 300.585 355.605 300.755 ;
        RECT 355.435 300.225 355.605 300.395 ;
        RECT 355.435 299.865 355.605 300.035 ;
        RECT 355.435 299.505 355.605 299.675 ;
        RECT 355.435 299.145 355.605 299.315 ;
        RECT 355.435 298.785 355.605 298.955 ;
        RECT 355.435 298.425 355.605 298.595 ;
        RECT 355.435 298.065 355.605 298.235 ;
        RECT 355.435 297.705 355.605 297.875 ;
        RECT 355.435 297.345 355.605 297.515 ;
        RECT 355.435 296.985 355.605 297.155 ;
        RECT 355.435 296.625 355.605 296.795 ;
        RECT 355.435 296.265 355.605 296.435 ;
        RECT 355.435 295.905 355.605 296.075 ;
        RECT 356.530 308.745 356.700 308.915 ;
        RECT 356.530 308.385 356.700 308.555 ;
        RECT 356.530 305.275 356.700 305.445 ;
        RECT 356.530 304.915 356.700 305.085 ;
        RECT 356.530 301.805 356.700 301.975 ;
        RECT 356.530 301.445 356.700 301.615 ;
        RECT 356.530 298.335 356.700 298.505 ;
        RECT 356.530 297.975 356.700 298.145 ;
        RECT 382.430 313.225 382.600 313.395 ;
        RECT 394.005 326.935 394.175 327.105 ;
        RECT 394.005 326.575 394.175 326.745 ;
        RECT 394.005 326.215 394.175 326.385 ;
        RECT 394.005 325.855 394.175 326.025 ;
        RECT 394.005 325.495 394.175 325.665 ;
        RECT 394.005 325.135 394.175 325.305 ;
        RECT 394.005 324.775 394.175 324.945 ;
        RECT 394.005 324.415 394.175 324.585 ;
        RECT 394.005 324.055 394.175 324.225 ;
        RECT 394.005 323.695 394.175 323.865 ;
        RECT 394.005 323.335 394.175 323.505 ;
        RECT 394.005 322.975 394.175 323.145 ;
        RECT 394.005 322.615 394.175 322.785 ;
        RECT 394.005 322.255 394.175 322.425 ;
        RECT 394.005 321.895 394.175 322.065 ;
        RECT 394.005 321.535 394.175 321.705 ;
        RECT 394.005 321.175 394.175 321.345 ;
        RECT 394.005 320.815 394.175 320.985 ;
        RECT 394.005 320.455 394.175 320.625 ;
        RECT 394.005 320.095 394.175 320.265 ;
        RECT 394.005 319.735 394.175 319.905 ;
        RECT 394.005 319.375 394.175 319.545 ;
        RECT 394.005 319.015 394.175 319.185 ;
        RECT 394.005 318.655 394.175 318.825 ;
        RECT 394.005 318.295 394.175 318.465 ;
        RECT 394.005 317.935 394.175 318.105 ;
        RECT 394.005 317.575 394.175 317.745 ;
        RECT 394.005 317.215 394.175 317.385 ;
        RECT 394.005 316.855 394.175 317.025 ;
        RECT 394.005 316.495 394.175 316.665 ;
        RECT 394.005 316.135 394.175 316.305 ;
        RECT 394.005 315.775 394.175 315.945 ;
        RECT 394.005 315.415 394.175 315.585 ;
        RECT 394.005 315.055 394.175 315.225 ;
        RECT 394.005 314.695 394.175 314.865 ;
        RECT 394.005 314.335 394.175 314.505 ;
        RECT 395.100 327.535 395.270 327.705 ;
        RECT 395.100 327.175 395.270 327.345 ;
        RECT 395.100 324.065 395.270 324.235 ;
        RECT 395.100 323.705 395.270 323.875 ;
        RECT 395.100 320.595 395.270 320.765 ;
        RECT 395.100 320.235 395.270 320.405 ;
        RECT 395.100 317.125 395.270 317.295 ;
        RECT 395.100 316.765 395.270 316.935 ;
        RECT 395.100 313.655 395.270 313.825 ;
        RECT 398.390 327.535 398.560 327.705 ;
        RECT 398.390 327.175 398.560 327.345 ;
        RECT 398.390 324.065 398.560 324.235 ;
        RECT 398.390 323.705 398.560 323.875 ;
        RECT 398.390 320.595 398.560 320.765 ;
        RECT 398.390 320.235 398.560 320.405 ;
        RECT 398.390 317.125 398.560 317.295 ;
        RECT 398.390 316.765 398.560 316.935 ;
        RECT 389.010 313.225 389.180 313.395 ;
        RECT 395.100 313.295 395.270 313.465 ;
        RECT 359.820 308.745 359.990 308.915 ;
        RECT 359.820 308.385 359.990 308.555 ;
        RECT 359.820 305.275 359.990 305.445 ;
        RECT 359.820 304.915 359.990 305.085 ;
        RECT 359.820 301.805 359.990 301.975 ;
        RECT 359.820 301.445 359.990 301.615 ;
        RECT 359.820 298.335 359.990 298.505 ;
        RECT 359.820 297.975 359.990 298.145 ;
        RECT 355.435 295.545 355.605 295.715 ;
        RECT 212.075 295.040 212.245 295.210 ;
        RECT 212.435 295.040 212.605 295.210 ;
        RECT 215.545 295.040 215.715 295.210 ;
        RECT 215.905 295.040 216.075 295.210 ;
        RECT 219.015 295.040 219.185 295.210 ;
        RECT 219.375 295.040 219.545 295.210 ;
        RECT 222.485 295.040 222.655 295.210 ;
        RECT 222.845 295.040 223.015 295.210 ;
        RECT 225.955 295.040 226.125 295.210 ;
        RECT 226.315 295.040 226.485 295.210 ;
        RECT 232.045 295.040 232.215 295.210 ;
        RECT 232.405 295.040 232.575 295.210 ;
        RECT 235.515 295.040 235.685 295.210 ;
        RECT 235.875 295.040 236.045 295.210 ;
        RECT 238.985 295.040 239.155 295.210 ;
        RECT 239.345 295.040 239.515 295.210 ;
        RECT 242.455 295.040 242.625 295.210 ;
        RECT 242.815 295.040 242.985 295.210 ;
        RECT 245.925 295.040 246.095 295.210 ;
        RECT 246.285 295.040 246.455 295.210 ;
        RECT 252.155 295.040 252.325 295.210 ;
        RECT 252.515 295.040 252.685 295.210 ;
        RECT 255.625 295.040 255.795 295.210 ;
        RECT 255.985 295.040 256.155 295.210 ;
        RECT 259.095 295.040 259.265 295.210 ;
        RECT 259.455 295.040 259.625 295.210 ;
        RECT 262.565 295.040 262.735 295.210 ;
        RECT 262.925 295.040 263.095 295.210 ;
        RECT 266.035 295.040 266.205 295.210 ;
        RECT 266.395 295.040 266.565 295.210 ;
        RECT 272.265 295.040 272.435 295.210 ;
        RECT 272.625 295.040 272.795 295.210 ;
        RECT 275.735 295.040 275.905 295.210 ;
        RECT 276.095 295.040 276.265 295.210 ;
        RECT 279.205 295.040 279.375 295.210 ;
        RECT 279.565 295.040 279.735 295.210 ;
        RECT 282.675 295.040 282.845 295.210 ;
        RECT 283.035 295.040 283.205 295.210 ;
        RECT 286.145 295.040 286.315 295.210 ;
        RECT 286.505 295.040 286.675 295.210 ;
        RECT 4.855 293.050 5.025 293.220 ;
        RECT 5.215 293.050 5.385 293.220 ;
        RECT 8.325 293.050 8.495 293.220 ;
        RECT 8.685 293.050 8.855 293.220 ;
        RECT 11.795 293.050 11.965 293.220 ;
        RECT 12.155 293.050 12.325 293.220 ;
        RECT 18.195 293.030 18.365 293.200 ;
        RECT 18.555 293.030 18.725 293.200 ;
        RECT 21.665 293.030 21.835 293.200 ;
        RECT 22.025 293.030 22.195 293.200 ;
        RECT 25.135 293.030 25.305 293.200 ;
        RECT 25.495 293.030 25.665 293.200 ;
        RECT 31.565 293.060 31.735 293.230 ;
        RECT 31.925 293.060 32.095 293.230 ;
        RECT 35.035 293.060 35.205 293.230 ;
        RECT 35.395 293.060 35.565 293.230 ;
        RECT 38.505 293.060 38.675 293.230 ;
        RECT 38.865 293.060 39.035 293.230 ;
        RECT 44.795 293.060 44.965 293.230 ;
        RECT 45.155 293.060 45.325 293.230 ;
        RECT 48.265 293.060 48.435 293.230 ;
        RECT 48.625 293.060 48.795 293.230 ;
        RECT 51.735 293.060 51.905 293.230 ;
        RECT 52.095 293.060 52.265 293.230 ;
        RECT 97.885 293.300 98.055 293.470 ;
        RECT 98.245 293.300 98.415 293.470 ;
        RECT 101.355 293.300 101.525 293.470 ;
        RECT 101.715 293.300 101.885 293.470 ;
        RECT 58.065 293.030 58.235 293.200 ;
        RECT 58.425 293.030 58.595 293.200 ;
        RECT 61.535 293.030 61.705 293.200 ;
        RECT 61.895 293.030 62.065 293.200 ;
        RECT 65.005 293.030 65.175 293.200 ;
        RECT 65.365 293.030 65.535 293.200 ;
        RECT 71.335 293.060 71.505 293.230 ;
        RECT 71.695 293.060 71.865 293.230 ;
        RECT 74.805 293.060 74.975 293.230 ;
        RECT 75.165 293.060 75.335 293.230 ;
        RECT 78.275 293.060 78.445 293.230 ;
        RECT 78.635 293.060 78.805 293.230 ;
        RECT 84.465 293.080 84.635 293.250 ;
        RECT 84.825 293.080 84.995 293.250 ;
        RECT 87.935 293.080 88.105 293.250 ;
        RECT 88.295 293.080 88.465 293.250 ;
        RECT 91.405 293.080 91.575 293.250 ;
        RECT 91.765 293.080 91.935 293.250 ;
        RECT 1.855 288.280 2.025 288.450 ;
        RECT 1.855 287.920 2.025 288.090 ;
        RECT 1.855 287.560 2.025 287.730 ;
        RECT 1.855 287.200 2.025 287.370 ;
        RECT 1.855 286.840 2.025 287.010 ;
        RECT 1.855 286.480 2.025 286.650 ;
        RECT 356.530 294.865 356.700 295.035 ;
        RECT 356.530 294.505 356.700 294.675 ;
        RECT 359.820 294.865 359.990 295.035 ;
        RECT 363.110 308.745 363.280 308.915 ;
        RECT 363.110 308.385 363.280 308.555 ;
        RECT 363.110 305.275 363.280 305.445 ;
        RECT 363.110 304.915 363.280 305.085 ;
        RECT 363.110 301.805 363.280 301.975 ;
        RECT 363.110 301.445 363.280 301.615 ;
        RECT 363.110 298.335 363.280 298.505 ;
        RECT 363.110 297.975 363.280 298.145 ;
        RECT 363.110 294.865 363.280 295.035 ;
        RECT 366.400 308.745 366.570 308.915 ;
        RECT 398.390 313.655 398.560 313.825 ;
        RECT 401.680 327.535 401.850 327.705 ;
        RECT 401.680 327.175 401.850 327.345 ;
        RECT 401.680 324.065 401.850 324.235 ;
        RECT 401.680 323.705 401.850 323.875 ;
        RECT 401.680 320.595 401.850 320.765 ;
        RECT 401.680 320.235 401.850 320.405 ;
        RECT 401.680 317.125 401.850 317.295 ;
        RECT 401.680 316.765 401.850 316.935 ;
        RECT 401.680 313.655 401.850 313.825 ;
        RECT 404.970 327.535 405.140 327.705 ;
        RECT 408.260 327.535 408.430 327.705 ;
        RECT 858.170 327.545 858.340 327.715 ;
        RECT 404.970 327.175 405.140 327.345 ;
        RECT 404.970 324.065 405.140 324.235 ;
        RECT 404.970 323.705 405.140 323.875 ;
        RECT 404.970 320.595 405.140 320.765 ;
        RECT 404.970 320.235 405.140 320.405 ;
        RECT 404.970 317.125 405.140 317.295 ;
        RECT 404.970 316.765 405.140 316.935 ;
        RECT 404.970 313.655 405.140 313.825 ;
        RECT 860.750 327.545 860.920 327.715 ;
        RECT 408.260 327.175 408.430 327.345 ;
        RECT 658.915 326.185 659.085 326.355 ;
        RECT 659.395 326.185 659.565 326.355 ;
        RECT 659.875 326.185 660.045 326.355 ;
        RECT 663.815 326.145 663.985 326.315 ;
        RECT 664.295 326.145 664.465 326.315 ;
        RECT 664.775 326.145 664.945 326.315 ;
        RECT 668.405 326.175 668.575 326.345 ;
        RECT 668.885 326.175 669.055 326.345 ;
        RECT 669.365 326.175 669.535 326.345 ;
        RECT 672.945 326.155 673.115 326.325 ;
        RECT 673.425 326.155 673.595 326.325 ;
        RECT 673.905 326.155 674.075 326.325 ;
        RECT 676.375 326.165 676.545 326.335 ;
        RECT 676.855 326.165 677.025 326.335 ;
        RECT 677.335 326.165 677.505 326.335 ;
        RECT 677.815 326.165 677.985 326.335 ;
        RECT 678.295 326.165 678.465 326.335 ;
        RECT 678.775 326.165 678.945 326.335 ;
        RECT 679.255 326.165 679.425 326.335 ;
        RECT 679.735 326.165 679.905 326.335 ;
        RECT 682.145 326.165 682.315 326.335 ;
        RECT 682.625 326.165 682.795 326.335 ;
        RECT 683.105 326.165 683.275 326.335 ;
        RECT 683.585 326.165 683.755 326.335 ;
        RECT 684.065 326.165 684.235 326.335 ;
        RECT 684.545 326.165 684.715 326.335 ;
        RECT 685.025 326.165 685.195 326.335 ;
        RECT 687.595 326.165 687.765 326.335 ;
        RECT 688.075 326.165 688.245 326.335 ;
        RECT 688.555 326.165 688.725 326.335 ;
        RECT 689.035 326.165 689.205 326.335 ;
        RECT 689.515 326.165 689.685 326.335 ;
        RECT 689.995 326.165 690.165 326.335 ;
        RECT 690.475 326.165 690.645 326.335 ;
        RECT 692.905 326.185 693.075 326.355 ;
        RECT 693.385 326.185 693.555 326.355 ;
        RECT 693.865 326.185 694.035 326.355 ;
        RECT 694.345 326.185 694.515 326.355 ;
        RECT 694.825 326.185 694.995 326.355 ;
        RECT 695.305 326.185 695.475 326.355 ;
        RECT 695.785 326.185 695.955 326.355 ;
        RECT 858.170 326.075 858.340 326.245 ;
        RECT 658.880 325.705 659.050 325.875 ;
        RECT 659.240 325.705 659.410 325.875 ;
        RECT 408.260 324.065 408.430 324.235 ;
        RECT 408.260 323.705 408.430 323.875 ;
        RECT 591.920 325.360 592.090 325.530 ;
        RECT 591.920 325.000 592.090 325.170 ;
        RECT 591.920 324.640 592.090 324.810 ;
        RECT 591.920 324.280 592.090 324.450 ;
        RECT 663.780 325.665 663.950 325.835 ;
        RECT 664.140 325.665 664.310 325.835 ;
        RECT 668.370 325.695 668.540 325.865 ;
        RECT 668.730 325.695 668.900 325.865 ;
        RECT 672.910 325.675 673.080 325.845 ;
        RECT 673.270 325.675 673.440 325.845 ;
        RECT 676.810 325.685 676.980 325.855 ;
        RECT 677.170 325.685 677.340 325.855 ;
        RECT 677.530 325.685 677.700 325.855 ;
        RECT 678.450 325.685 678.620 325.855 ;
        RECT 678.810 325.685 678.980 325.855 ;
        RECT 679.170 325.685 679.340 325.855 ;
        RECT 682.100 325.685 682.270 325.855 ;
        RECT 682.460 325.685 682.630 325.855 ;
        RECT 682.820 325.685 682.990 325.855 ;
        RECT 683.540 325.685 683.710 325.855 ;
        RECT 683.900 325.685 684.070 325.855 ;
        RECT 684.260 325.685 684.430 325.855 ;
        RECT 684.620 325.685 684.790 325.855 ;
        RECT 687.550 325.685 687.720 325.855 ;
        RECT 687.910 325.685 688.080 325.855 ;
        RECT 688.270 325.685 688.440 325.855 ;
        RECT 688.990 325.685 689.160 325.855 ;
        RECT 689.350 325.685 689.520 325.855 ;
        RECT 689.710 325.685 689.880 325.855 ;
        RECT 690.070 325.685 690.240 325.855 ;
        RECT 860.750 326.075 860.920 326.245 ;
        RECT 693.580 325.705 693.750 325.875 ;
        RECT 693.940 325.705 694.110 325.875 ;
        RECT 694.300 325.705 694.470 325.875 ;
        RECT 694.660 325.705 694.830 325.875 ;
        RECT 695.020 325.705 695.190 325.875 ;
        RECT 695.380 325.705 695.550 325.875 ;
        RECT 858.170 324.605 858.340 324.775 ;
        RECT 860.750 324.605 860.920 324.775 ;
        RECT 591.920 323.920 592.090 324.090 ;
        RECT 591.920 323.560 592.090 323.730 ;
        RECT 858.170 323.135 858.340 323.305 ;
        RECT 860.750 323.135 860.920 323.305 ;
        RECT 858.170 321.665 858.340 321.835 ;
        RECT 860.750 321.665 860.920 321.835 ;
        RECT 408.260 320.595 408.430 320.765 ;
        RECT 864.740 320.575 864.910 320.745 ;
        RECT 408.260 320.235 408.430 320.405 ;
        RECT 661.555 320.305 661.725 320.475 ;
        RECT 662.035 320.305 662.205 320.475 ;
        RECT 662.515 320.305 662.685 320.475 ;
        RECT 662.995 320.305 663.165 320.475 ;
        RECT 663.475 320.305 663.645 320.475 ;
        RECT 663.955 320.305 664.125 320.475 ;
        RECT 664.435 320.305 664.605 320.475 ;
        RECT 664.915 320.305 665.085 320.475 ;
        RECT 667.375 320.315 667.545 320.485 ;
        RECT 667.855 320.315 668.025 320.485 ;
        RECT 668.335 320.315 668.505 320.485 ;
        RECT 668.815 320.315 668.985 320.485 ;
        RECT 669.295 320.315 669.465 320.485 ;
        RECT 669.775 320.315 669.945 320.485 ;
        RECT 670.255 320.315 670.425 320.485 ;
        RECT 672.815 320.325 672.985 320.495 ;
        RECT 673.295 320.325 673.465 320.495 ;
        RECT 673.775 320.325 673.945 320.495 ;
        RECT 674.255 320.325 674.425 320.495 ;
        RECT 674.735 320.325 674.905 320.495 ;
        RECT 675.215 320.325 675.385 320.495 ;
        RECT 675.695 320.325 675.865 320.495 ;
        RECT 678.135 320.325 678.305 320.495 ;
        RECT 678.615 320.325 678.785 320.495 ;
        RECT 679.095 320.325 679.265 320.495 ;
        RECT 679.575 320.325 679.745 320.495 ;
        RECT 680.055 320.325 680.225 320.495 ;
        RECT 680.535 320.325 680.705 320.495 ;
        RECT 681.015 320.325 681.185 320.495 ;
        RECT 683.485 320.325 683.655 320.495 ;
        RECT 683.965 320.325 684.135 320.495 ;
        RECT 684.445 320.325 684.615 320.495 ;
        RECT 684.925 320.325 685.095 320.495 ;
        RECT 685.405 320.325 685.575 320.495 ;
        RECT 685.885 320.325 686.055 320.495 ;
        RECT 686.365 320.325 686.535 320.495 ;
        RECT 689.305 320.305 689.475 320.475 ;
        RECT 689.785 320.305 689.955 320.475 ;
        RECT 690.265 320.305 690.435 320.475 ;
        RECT 690.745 320.305 690.915 320.475 ;
        RECT 691.225 320.305 691.395 320.475 ;
        RECT 661.990 319.825 662.160 319.995 ;
        RECT 662.350 319.825 662.520 319.995 ;
        RECT 662.710 319.825 662.880 319.995 ;
        RECT 663.630 319.825 663.800 319.995 ;
        RECT 663.990 319.825 664.160 319.995 ;
        RECT 664.350 319.825 664.520 319.995 ;
        RECT 667.330 319.835 667.500 320.005 ;
        RECT 667.690 319.835 667.860 320.005 ;
        RECT 668.050 319.835 668.220 320.005 ;
        RECT 668.770 319.835 668.940 320.005 ;
        RECT 669.130 319.835 669.300 320.005 ;
        RECT 669.490 319.835 669.660 320.005 ;
        RECT 669.850 319.835 670.020 320.005 ;
        RECT 672.770 319.845 672.940 320.015 ;
        RECT 673.130 319.845 673.300 320.015 ;
        RECT 673.490 319.845 673.660 320.015 ;
        RECT 674.210 319.845 674.380 320.015 ;
        RECT 674.570 319.845 674.740 320.015 ;
        RECT 674.930 319.845 675.100 320.015 ;
        RECT 675.290 319.845 675.460 320.015 ;
        RECT 678.810 319.845 678.980 320.015 ;
        RECT 679.170 319.845 679.340 320.015 ;
        RECT 679.530 319.845 679.700 320.015 ;
        RECT 679.890 319.845 680.060 320.015 ;
        RECT 680.250 319.845 680.420 320.015 ;
        RECT 680.610 319.845 680.780 320.015 ;
        RECT 683.440 319.845 683.610 320.015 ;
        RECT 683.800 319.845 683.970 320.015 ;
        RECT 684.160 319.845 684.330 320.015 ;
        RECT 684.880 319.845 685.050 320.015 ;
        RECT 685.240 319.845 685.410 320.015 ;
        RECT 685.600 319.845 685.770 320.015 ;
        RECT 685.960 319.845 686.130 320.015 ;
        RECT 690.280 319.825 690.450 319.995 ;
        RECT 690.640 319.825 690.810 319.995 ;
        RECT 693.705 320.305 693.875 320.475 ;
        RECT 694.185 320.305 694.355 320.475 ;
        RECT 694.665 320.305 694.835 320.475 ;
        RECT 695.145 320.305 695.315 320.475 ;
        RECT 695.625 320.305 695.795 320.475 ;
        RECT 858.170 320.195 858.340 320.365 ;
        RECT 867.320 320.575 867.490 320.745 ;
        RECT 868.680 320.565 868.850 320.735 ;
        RECT 871.260 320.565 871.430 320.735 ;
        RECT 860.750 320.195 860.920 320.365 ;
        RECT 694.680 319.825 694.850 319.995 ;
        RECT 695.040 319.825 695.210 319.995 ;
        RECT 864.740 319.105 864.910 319.275 ;
        RECT 858.170 318.725 858.340 318.895 ;
        RECT 867.320 319.105 867.490 319.275 ;
        RECT 868.680 319.095 868.850 319.265 ;
        RECT 871.260 319.095 871.430 319.265 ;
        RECT 860.750 318.725 860.920 318.895 ;
        RECT 871.970 318.370 872.140 318.540 ;
        RECT 871.970 318.010 872.140 318.180 ;
        RECT 864.740 317.635 864.910 317.805 ;
        RECT 408.260 317.125 408.430 317.295 ;
        RECT 858.170 317.255 858.340 317.425 ;
        RECT 867.320 317.635 867.490 317.805 ;
        RECT 868.680 317.625 868.850 317.795 ;
        RECT 871.260 317.625 871.430 317.795 ;
        RECT 871.970 317.650 872.140 317.820 ;
        RECT 860.750 317.255 860.920 317.425 ;
        RECT 871.970 317.290 872.140 317.460 ;
        RECT 408.260 316.765 408.430 316.935 ;
        RECT 871.970 316.930 872.140 317.100 ;
        RECT 871.970 316.570 872.140 316.740 ;
        RECT 864.740 316.165 864.910 316.335 ;
        RECT 858.170 315.785 858.340 315.955 ;
        RECT 867.320 316.165 867.490 316.335 ;
        RECT 868.680 316.155 868.850 316.325 ;
        RECT 871.260 316.155 871.430 316.325 ;
        RECT 871.970 316.210 872.140 316.380 ;
        RECT 860.750 315.785 860.920 315.955 ;
        RECT 871.970 315.850 872.140 316.020 ;
        RECT 871.970 315.490 872.140 315.660 ;
        RECT 398.390 313.295 398.560 313.465 ;
        RECT 401.680 313.295 401.850 313.465 ;
        RECT 404.970 313.295 405.140 313.465 ;
        RECT 408.260 313.655 408.430 313.825 ;
        RECT 408.260 313.295 408.430 313.465 ;
        RECT 864.740 314.695 864.910 314.865 ;
        RECT 601.300 313.995 601.470 314.165 ;
        RECT 602.480 314.005 602.650 314.175 ;
        RECT 604.060 314.005 604.230 314.175 ;
        RECT 605.640 314.005 605.810 314.175 ;
        RECT 607.000 314.015 607.170 314.185 ;
        RECT 608.580 314.015 608.750 314.185 ;
        RECT 610.160 314.015 610.330 314.185 ;
        RECT 611.520 314.015 611.690 314.185 ;
        RECT 613.100 314.015 613.270 314.185 ;
        RECT 614.680 314.015 614.850 314.185 ;
        RECT 615.950 313.995 616.120 314.165 ;
        RECT 617.530 313.995 617.700 314.165 ;
        RECT 619.110 313.995 619.280 314.165 ;
        RECT 620.330 314.005 620.500 314.175 ;
        RECT 621.910 314.005 622.080 314.175 ;
        RECT 623.490 314.005 623.660 314.175 ;
        RECT 624.650 313.995 624.820 314.165 ;
        RECT 626.230 313.995 626.400 314.165 ;
        RECT 627.810 313.995 627.980 314.165 ;
        RECT 629.030 314.225 629.200 314.395 ;
        RECT 858.170 314.315 858.340 314.485 ;
        RECT 867.320 314.695 867.490 314.865 ;
        RECT 868.680 314.685 868.850 314.855 ;
        RECT 871.260 314.685 871.430 314.855 ;
        RECT 860.750 314.315 860.920 314.485 ;
        RECT 601.300 313.635 601.470 313.805 ;
        RECT 601.300 313.275 601.470 313.445 ;
        RECT 601.300 312.915 601.470 313.085 ;
        RECT 629.030 313.865 629.200 314.035 ;
        RECT 629.030 313.505 629.200 313.675 ;
        RECT 629.030 313.145 629.200 313.315 ;
        RECT 635.265 312.975 635.435 313.145 ;
        RECT 635.745 312.975 635.915 313.145 ;
        RECT 636.225 312.975 636.395 313.145 ;
        RECT 639.455 313.065 639.625 313.235 ;
        RECT 639.935 313.065 640.105 313.235 ;
        RECT 640.415 313.065 640.585 313.235 ;
        RECT 643.555 313.045 643.725 313.215 ;
        RECT 644.035 313.045 644.205 313.215 ;
        RECT 644.515 313.045 644.685 313.215 ;
        RECT 595.375 312.525 595.545 312.695 ;
        RECT 595.855 312.525 596.025 312.695 ;
        RECT 596.335 312.525 596.505 312.695 ;
        RECT 601.300 312.555 601.470 312.725 ;
        RECT 596.010 312.045 596.180 312.215 ;
        RECT 596.370 312.045 596.540 312.215 ;
        RECT 602.480 312.535 602.650 312.705 ;
        RECT 604.060 312.535 604.230 312.705 ;
        RECT 605.640 312.535 605.810 312.705 ;
        RECT 607.000 312.545 607.170 312.715 ;
        RECT 608.580 312.545 608.750 312.715 ;
        RECT 610.160 312.545 610.330 312.715 ;
        RECT 611.520 312.545 611.690 312.715 ;
        RECT 613.100 312.545 613.270 312.715 ;
        RECT 614.680 312.545 614.850 312.715 ;
        RECT 615.950 312.525 616.120 312.695 ;
        RECT 617.530 312.525 617.700 312.695 ;
        RECT 619.110 312.525 619.280 312.695 ;
        RECT 620.330 312.535 620.500 312.705 ;
        RECT 621.910 312.535 622.080 312.705 ;
        RECT 623.490 312.535 623.660 312.705 ;
        RECT 624.650 312.525 624.820 312.695 ;
        RECT 626.230 312.525 626.400 312.695 ;
        RECT 627.810 312.525 627.980 312.695 ;
        RECT 629.030 312.785 629.200 312.955 ;
        RECT 629.030 312.425 629.200 312.595 ;
        RECT 635.230 312.495 635.400 312.665 ;
        RECT 635.590 312.495 635.760 312.665 ;
        RECT 639.420 312.585 639.590 312.755 ;
        RECT 639.780 312.585 639.950 312.755 ;
        RECT 643.520 312.565 643.690 312.735 ;
        RECT 643.880 312.565 644.050 312.735 ;
        RECT 369.690 308.745 369.860 308.915 ;
        RECT 366.400 308.385 366.570 308.555 ;
        RECT 366.400 305.275 366.570 305.445 ;
        RECT 366.400 304.915 366.570 305.085 ;
        RECT 366.400 301.805 366.570 301.975 ;
        RECT 366.400 301.445 366.570 301.615 ;
        RECT 366.400 298.335 366.570 298.505 ;
        RECT 366.400 297.975 366.570 298.145 ;
        RECT 366.400 294.865 366.570 295.035 ;
        RECT 369.690 308.385 369.860 308.555 ;
        RECT 369.690 305.275 369.860 305.445 ;
        RECT 369.690 304.915 369.860 305.085 ;
        RECT 369.690 301.805 369.860 301.975 ;
        RECT 369.690 301.445 369.860 301.615 ;
        RECT 369.690 298.335 369.860 298.505 ;
        RECT 369.690 297.975 369.860 298.145 ;
        RECT 359.820 294.505 359.990 294.675 ;
        RECT 363.110 294.505 363.280 294.675 ;
        RECT 366.400 294.505 366.570 294.675 ;
        RECT 369.690 294.865 369.860 295.035 ;
        RECT 374.755 308.045 374.925 308.215 ;
        RECT 374.755 307.685 374.925 307.855 ;
        RECT 374.755 307.325 374.925 307.495 ;
        RECT 374.755 306.965 374.925 307.135 ;
        RECT 374.755 306.605 374.925 306.775 ;
        RECT 374.755 306.245 374.925 306.415 ;
        RECT 374.755 305.885 374.925 306.055 ;
        RECT 374.755 305.525 374.925 305.695 ;
        RECT 374.755 305.165 374.925 305.335 ;
        RECT 374.755 304.805 374.925 304.975 ;
        RECT 374.755 304.445 374.925 304.615 ;
        RECT 374.755 304.085 374.925 304.255 ;
        RECT 374.755 303.725 374.925 303.895 ;
        RECT 374.755 303.365 374.925 303.535 ;
        RECT 374.755 303.005 374.925 303.175 ;
        RECT 374.755 302.645 374.925 302.815 ;
        RECT 374.755 302.285 374.925 302.455 ;
        RECT 374.755 301.925 374.925 302.095 ;
        RECT 374.755 301.565 374.925 301.735 ;
        RECT 374.755 301.205 374.925 301.375 ;
        RECT 374.755 300.845 374.925 301.015 ;
        RECT 374.755 300.485 374.925 300.655 ;
        RECT 374.755 300.125 374.925 300.295 ;
        RECT 374.755 299.765 374.925 299.935 ;
        RECT 374.755 299.405 374.925 299.575 ;
        RECT 374.755 299.045 374.925 299.215 ;
        RECT 374.755 298.685 374.925 298.855 ;
        RECT 374.755 298.325 374.925 298.495 ;
        RECT 374.755 297.965 374.925 298.135 ;
        RECT 374.755 297.605 374.925 297.775 ;
        RECT 374.755 297.245 374.925 297.415 ;
        RECT 374.755 296.885 374.925 297.055 ;
        RECT 374.755 296.525 374.925 296.695 ;
        RECT 374.755 296.165 374.925 296.335 ;
        RECT 374.755 295.805 374.925 295.975 ;
        RECT 375.850 308.645 376.020 308.815 ;
        RECT 375.850 308.285 376.020 308.455 ;
        RECT 375.850 305.175 376.020 305.345 ;
        RECT 375.850 304.815 376.020 304.985 ;
        RECT 375.850 301.705 376.020 301.875 ;
        RECT 375.850 301.345 376.020 301.515 ;
        RECT 375.850 298.235 376.020 298.405 ;
        RECT 375.850 297.875 376.020 298.045 ;
        RECT 382.430 308.645 382.600 308.815 ;
        RECT 389.010 308.645 389.180 308.815 ;
        RECT 382.430 308.285 382.600 308.455 ;
        RECT 382.430 305.175 382.600 305.345 ;
        RECT 382.430 304.815 382.600 304.985 ;
        RECT 382.430 301.705 382.600 301.875 ;
        RECT 382.430 301.345 382.600 301.515 ;
        RECT 382.430 298.235 382.600 298.405 ;
        RECT 382.430 297.875 382.600 298.045 ;
        RECT 374.755 295.445 374.925 295.615 ;
        RECT 375.850 294.765 376.020 294.935 ;
        RECT 369.690 294.505 369.860 294.675 ;
        RECT 382.430 294.765 382.600 294.935 ;
        RECT 389.010 308.285 389.180 308.455 ;
        RECT 389.010 305.175 389.180 305.345 ;
        RECT 389.010 304.815 389.180 304.985 ;
        RECT 389.010 301.705 389.180 301.875 ;
        RECT 389.010 301.345 389.180 301.515 ;
        RECT 389.010 298.235 389.180 298.405 ;
        RECT 389.010 297.875 389.180 298.045 ;
        RECT 389.010 294.765 389.180 294.935 ;
        RECT 375.850 294.405 376.020 294.575 ;
        RECT 355.435 289.265 355.605 289.435 ;
        RECT 355.435 288.905 355.605 289.075 ;
        RECT 212.075 288.460 212.245 288.630 ;
        RECT 212.435 288.460 212.605 288.630 ;
        RECT 215.545 288.460 215.715 288.630 ;
        RECT 215.905 288.460 216.075 288.630 ;
        RECT 219.015 288.460 219.185 288.630 ;
        RECT 219.375 288.460 219.545 288.630 ;
        RECT 222.485 288.460 222.655 288.630 ;
        RECT 222.845 288.460 223.015 288.630 ;
        RECT 225.955 288.460 226.125 288.630 ;
        RECT 226.315 288.460 226.485 288.630 ;
        RECT 232.045 288.460 232.215 288.630 ;
        RECT 232.405 288.460 232.575 288.630 ;
        RECT 235.515 288.460 235.685 288.630 ;
        RECT 235.875 288.460 236.045 288.630 ;
        RECT 238.985 288.460 239.155 288.630 ;
        RECT 239.345 288.460 239.515 288.630 ;
        RECT 242.455 288.460 242.625 288.630 ;
        RECT 242.815 288.460 242.985 288.630 ;
        RECT 245.925 288.460 246.095 288.630 ;
        RECT 246.285 288.460 246.455 288.630 ;
        RECT 252.155 288.460 252.325 288.630 ;
        RECT 252.515 288.460 252.685 288.630 ;
        RECT 255.625 288.460 255.795 288.630 ;
        RECT 255.985 288.460 256.155 288.630 ;
        RECT 259.095 288.460 259.265 288.630 ;
        RECT 259.455 288.460 259.625 288.630 ;
        RECT 262.565 288.460 262.735 288.630 ;
        RECT 262.925 288.460 263.095 288.630 ;
        RECT 266.035 288.460 266.205 288.630 ;
        RECT 266.395 288.460 266.565 288.630 ;
        RECT 272.265 288.460 272.435 288.630 ;
        RECT 272.625 288.460 272.795 288.630 ;
        RECT 275.735 288.460 275.905 288.630 ;
        RECT 276.095 288.460 276.265 288.630 ;
        RECT 279.205 288.460 279.375 288.630 ;
        RECT 279.565 288.460 279.735 288.630 ;
        RECT 282.675 288.460 282.845 288.630 ;
        RECT 283.035 288.460 283.205 288.630 ;
        RECT 286.145 288.460 286.315 288.630 ;
        RECT 286.505 288.460 286.675 288.630 ;
        RECT 355.435 288.545 355.605 288.715 ;
        RECT 355.435 288.185 355.605 288.355 ;
        RECT 355.435 287.825 355.605 287.995 ;
        RECT 355.435 287.465 355.605 287.635 ;
        RECT 355.435 287.105 355.605 287.275 ;
        RECT 97.885 286.720 98.055 286.890 ;
        RECT 98.245 286.720 98.415 286.890 ;
        RECT 101.355 286.720 101.525 286.890 ;
        RECT 101.715 286.720 101.885 286.890 ;
        RECT 355.435 286.745 355.605 286.915 ;
        RECT 4.855 286.470 5.025 286.640 ;
        RECT 5.215 286.470 5.385 286.640 ;
        RECT 8.325 286.470 8.495 286.640 ;
        RECT 8.685 286.470 8.855 286.640 ;
        RECT 11.795 286.470 11.965 286.640 ;
        RECT 12.155 286.470 12.325 286.640 ;
        RECT 18.195 286.450 18.365 286.620 ;
        RECT 18.555 286.450 18.725 286.620 ;
        RECT 21.665 286.450 21.835 286.620 ;
        RECT 22.025 286.450 22.195 286.620 ;
        RECT 25.135 286.450 25.305 286.620 ;
        RECT 25.495 286.450 25.665 286.620 ;
        RECT 31.565 286.480 31.735 286.650 ;
        RECT 31.925 286.480 32.095 286.650 ;
        RECT 35.035 286.480 35.205 286.650 ;
        RECT 35.395 286.480 35.565 286.650 ;
        RECT 38.505 286.480 38.675 286.650 ;
        RECT 38.865 286.480 39.035 286.650 ;
        RECT 44.795 286.480 44.965 286.650 ;
        RECT 45.155 286.480 45.325 286.650 ;
        RECT 48.265 286.480 48.435 286.650 ;
        RECT 48.625 286.480 48.795 286.650 ;
        RECT 51.735 286.480 51.905 286.650 ;
        RECT 52.095 286.480 52.265 286.650 ;
        RECT 1.855 286.120 2.025 286.290 ;
        RECT 58.065 286.450 58.235 286.620 ;
        RECT 58.425 286.450 58.595 286.620 ;
        RECT 61.535 286.450 61.705 286.620 ;
        RECT 61.895 286.450 62.065 286.620 ;
        RECT 65.005 286.450 65.175 286.620 ;
        RECT 65.365 286.450 65.535 286.620 ;
        RECT 71.335 286.480 71.505 286.650 ;
        RECT 71.695 286.480 71.865 286.650 ;
        RECT 74.805 286.480 74.975 286.650 ;
        RECT 75.165 286.480 75.335 286.650 ;
        RECT 78.275 286.480 78.445 286.650 ;
        RECT 78.635 286.480 78.805 286.650 ;
        RECT 84.465 286.500 84.635 286.670 ;
        RECT 84.825 286.500 84.995 286.670 ;
        RECT 87.935 286.500 88.105 286.670 ;
        RECT 88.295 286.500 88.465 286.670 ;
        RECT 91.405 286.500 91.575 286.670 ;
        RECT 91.765 286.500 91.935 286.670 ;
        RECT 1.855 285.760 2.025 285.930 ;
        RECT 1.855 285.400 2.025 285.570 ;
        RECT 1.855 285.040 2.025 285.210 ;
        RECT 1.855 284.680 2.025 284.850 ;
        RECT 1.855 284.320 2.025 284.490 ;
        RECT 1.855 283.960 2.025 284.130 ;
        RECT 355.435 286.385 355.605 286.555 ;
        RECT 355.435 286.025 355.605 286.195 ;
        RECT 355.435 285.665 355.605 285.835 ;
        RECT 355.435 285.305 355.605 285.475 ;
        RECT 355.435 284.945 355.605 285.115 ;
        RECT 355.435 284.585 355.605 284.755 ;
        RECT 355.435 284.225 355.605 284.395 ;
        RECT 355.435 283.865 355.605 284.035 ;
        RECT 355.435 283.505 355.605 283.675 ;
        RECT 355.435 283.145 355.605 283.315 ;
        RECT 355.435 282.785 355.605 282.955 ;
        RECT 215.010 281.150 225.620 282.040 ;
        RECT 235.050 281.140 245.660 282.030 ;
        RECT 255.110 281.140 265.720 282.030 ;
        RECT 275.160 281.140 285.770 282.030 ;
        RECT 355.435 282.425 355.605 282.595 ;
        RECT 355.435 282.065 355.605 282.235 ;
        RECT 355.435 281.705 355.605 281.875 ;
        RECT 355.435 281.345 355.605 281.515 ;
        RECT 355.435 280.985 355.605 281.155 ;
        RECT 355.435 280.625 355.605 280.795 ;
        RECT 4.855 279.890 5.025 280.060 ;
        RECT 5.215 279.890 5.385 280.060 ;
        RECT 8.325 279.890 8.495 280.060 ;
        RECT 8.685 279.890 8.855 280.060 ;
        RECT 11.795 279.890 11.965 280.060 ;
        RECT 12.155 279.890 12.325 280.060 ;
        RECT 97.885 280.140 98.055 280.310 ;
        RECT 98.245 280.140 98.415 280.310 ;
        RECT 101.355 280.140 101.525 280.310 ;
        RECT 101.715 280.140 101.885 280.310 ;
        RECT 355.435 280.265 355.605 280.435 ;
        RECT 18.195 279.870 18.365 280.040 ;
        RECT 18.555 279.870 18.725 280.040 ;
        RECT 21.665 279.870 21.835 280.040 ;
        RECT 22.025 279.870 22.195 280.040 ;
        RECT 25.135 279.870 25.305 280.040 ;
        RECT 25.495 279.870 25.665 280.040 ;
        RECT 31.565 279.900 31.735 280.070 ;
        RECT 31.925 279.900 32.095 280.070 ;
        RECT 35.035 279.900 35.205 280.070 ;
        RECT 35.395 279.900 35.565 280.070 ;
        RECT 38.505 279.900 38.675 280.070 ;
        RECT 38.865 279.900 39.035 280.070 ;
        RECT 44.795 279.900 44.965 280.070 ;
        RECT 45.155 279.900 45.325 280.070 ;
        RECT 48.265 279.900 48.435 280.070 ;
        RECT 48.625 279.900 48.795 280.070 ;
        RECT 51.735 279.900 51.905 280.070 ;
        RECT 52.095 279.900 52.265 280.070 ;
        RECT 58.065 279.870 58.235 280.040 ;
        RECT 58.425 279.870 58.595 280.040 ;
        RECT 61.535 279.870 61.705 280.040 ;
        RECT 61.895 279.870 62.065 280.040 ;
        RECT 65.005 279.870 65.175 280.040 ;
        RECT 65.365 279.870 65.535 280.040 ;
        RECT 71.335 279.900 71.505 280.070 ;
        RECT 71.695 279.900 71.865 280.070 ;
        RECT 74.805 279.900 74.975 280.070 ;
        RECT 75.165 279.900 75.335 280.070 ;
        RECT 78.275 279.900 78.445 280.070 ;
        RECT 78.635 279.900 78.805 280.070 ;
        RECT 84.465 279.920 84.635 280.090 ;
        RECT 84.825 279.920 84.995 280.090 ;
        RECT 87.935 279.920 88.105 280.090 ;
        RECT 88.295 279.920 88.465 280.090 ;
        RECT 91.405 279.920 91.575 280.090 ;
        RECT 91.765 279.920 91.935 280.090 ;
        RECT 4.855 273.310 5.025 273.480 ;
        RECT 5.215 273.310 5.385 273.480 ;
        RECT 8.325 273.310 8.495 273.480 ;
        RECT 8.685 273.310 8.855 273.480 ;
        RECT 11.795 273.310 11.965 273.480 ;
        RECT 12.155 273.310 12.325 273.480 ;
        RECT 15.390 272.320 16.280 273.930 ;
        RECT 18.195 273.290 18.365 273.460 ;
        RECT 18.555 273.290 18.725 273.460 ;
        RECT 21.665 273.290 21.835 273.460 ;
        RECT 22.025 273.290 22.195 273.460 ;
        RECT 25.135 273.290 25.305 273.460 ;
        RECT 25.495 273.290 25.665 273.460 ;
        RECT 28.605 272.470 29.495 274.080 ;
        RECT 31.565 273.320 31.735 273.490 ;
        RECT 31.925 273.320 32.095 273.490 ;
        RECT 35.035 273.320 35.205 273.490 ;
        RECT 35.395 273.320 35.565 273.490 ;
        RECT 38.505 273.320 38.675 273.490 ;
        RECT 38.865 273.320 39.035 273.490 ;
        RECT 41.820 272.175 42.710 274.505 ;
        RECT 44.795 273.320 44.965 273.490 ;
        RECT 45.155 273.320 45.325 273.490 ;
        RECT 48.265 273.320 48.435 273.490 ;
        RECT 48.625 273.320 48.795 273.490 ;
        RECT 51.735 273.320 51.905 273.490 ;
        RECT 52.095 273.320 52.265 273.490 ;
        RECT 55.240 272.060 56.130 274.030 ;
        RECT 58.065 273.290 58.235 273.460 ;
        RECT 58.425 273.290 58.595 273.460 ;
        RECT 61.535 273.290 61.705 273.460 ;
        RECT 61.895 273.290 62.065 273.460 ;
        RECT 65.005 273.290 65.175 273.460 ;
        RECT 65.365 273.290 65.535 273.460 ;
        RECT 68.545 272.245 69.075 274.215 ;
        RECT 71.335 273.320 71.505 273.490 ;
        RECT 71.695 273.320 71.865 273.490 ;
        RECT 74.805 273.320 74.975 273.490 ;
        RECT 75.165 273.320 75.335 273.490 ;
        RECT 78.275 273.320 78.445 273.490 ;
        RECT 78.635 273.320 78.805 273.490 ;
        RECT 81.480 272.710 82.730 273.960 ;
        RECT 84.465 273.340 84.635 273.510 ;
        RECT 84.825 273.340 84.995 273.510 ;
        RECT 87.935 273.340 88.105 273.510 ;
        RECT 88.295 273.340 88.465 273.510 ;
        RECT 91.405 273.340 91.575 273.510 ;
        RECT 91.765 273.340 91.935 273.510 ;
        RECT 94.300 272.800 95.190 274.410 ;
        RECT 211.835 279.670 212.005 279.840 ;
        RECT 212.195 279.670 212.365 279.840 ;
        RECT 215.305 279.670 215.475 279.840 ;
        RECT 215.665 279.670 215.835 279.840 ;
        RECT 218.775 279.670 218.945 279.840 ;
        RECT 219.135 279.670 219.305 279.840 ;
        RECT 222.245 279.670 222.415 279.840 ;
        RECT 222.605 279.670 222.775 279.840 ;
        RECT 225.715 279.670 225.885 279.840 ;
        RECT 226.075 279.670 226.245 279.840 ;
        RECT 231.875 279.660 232.045 279.830 ;
        RECT 232.235 279.660 232.405 279.830 ;
        RECT 235.345 279.660 235.515 279.830 ;
        RECT 235.705 279.660 235.875 279.830 ;
        RECT 238.815 279.660 238.985 279.830 ;
        RECT 239.175 279.660 239.345 279.830 ;
        RECT 242.285 279.660 242.455 279.830 ;
        RECT 242.645 279.660 242.815 279.830 ;
        RECT 245.755 279.660 245.925 279.830 ;
        RECT 246.115 279.660 246.285 279.830 ;
        RECT 251.935 279.660 252.105 279.830 ;
        RECT 252.295 279.660 252.465 279.830 ;
        RECT 255.405 279.660 255.575 279.830 ;
        RECT 255.765 279.660 255.935 279.830 ;
        RECT 258.875 279.660 259.045 279.830 ;
        RECT 259.235 279.660 259.405 279.830 ;
        RECT 262.345 279.660 262.515 279.830 ;
        RECT 262.705 279.660 262.875 279.830 ;
        RECT 265.815 279.660 265.985 279.830 ;
        RECT 266.175 279.660 266.345 279.830 ;
        RECT 271.985 279.660 272.155 279.830 ;
        RECT 272.345 279.660 272.515 279.830 ;
        RECT 275.455 279.660 275.625 279.830 ;
        RECT 275.815 279.660 275.985 279.830 ;
        RECT 278.925 279.660 279.095 279.830 ;
        RECT 279.285 279.660 279.455 279.830 ;
        RECT 282.395 279.660 282.565 279.830 ;
        RECT 282.755 279.660 282.925 279.830 ;
        RECT 285.865 279.660 286.035 279.830 ;
        RECT 286.225 279.660 286.395 279.830 ;
        RECT 211.835 276.380 212.005 276.550 ;
        RECT 212.195 276.380 212.365 276.550 ;
        RECT 215.305 276.380 215.475 276.550 ;
        RECT 215.665 276.380 215.835 276.550 ;
        RECT 218.775 276.380 218.945 276.550 ;
        RECT 219.135 276.380 219.305 276.550 ;
        RECT 222.245 276.380 222.415 276.550 ;
        RECT 222.605 276.380 222.775 276.550 ;
        RECT 225.715 276.380 225.885 276.550 ;
        RECT 226.075 276.380 226.245 276.550 ;
        RECT 97.885 273.560 98.055 273.730 ;
        RECT 98.245 273.560 98.415 273.730 ;
        RECT 101.355 273.560 101.525 273.730 ;
        RECT 101.715 273.560 101.885 273.730 ;
        RECT 355.435 279.905 355.605 280.075 ;
        RECT 231.875 276.370 232.045 276.540 ;
        RECT 232.235 276.370 232.405 276.540 ;
        RECT 235.345 276.370 235.515 276.540 ;
        RECT 235.705 276.370 235.875 276.540 ;
        RECT 238.815 276.370 238.985 276.540 ;
        RECT 239.175 276.370 239.345 276.540 ;
        RECT 242.285 276.370 242.455 276.540 ;
        RECT 242.645 276.370 242.815 276.540 ;
        RECT 245.755 276.370 245.925 276.540 ;
        RECT 246.115 276.370 246.285 276.540 ;
        RECT 211.835 273.090 212.005 273.260 ;
        RECT 212.195 273.090 212.365 273.260 ;
        RECT 215.305 273.090 215.475 273.260 ;
        RECT 215.665 273.090 215.835 273.260 ;
        RECT 218.775 273.090 218.945 273.260 ;
        RECT 219.135 273.090 219.305 273.260 ;
        RECT 222.245 273.090 222.415 273.260 ;
        RECT 222.605 273.090 222.775 273.260 ;
        RECT 225.715 273.090 225.885 273.260 ;
        RECT 226.075 273.090 226.245 273.260 ;
        RECT 211.835 269.800 212.005 269.970 ;
        RECT 212.195 269.800 212.365 269.970 ;
        RECT 215.305 269.800 215.475 269.970 ;
        RECT 215.665 269.800 215.835 269.970 ;
        RECT 218.775 269.800 218.945 269.970 ;
        RECT 219.135 269.800 219.305 269.970 ;
        RECT 222.245 269.800 222.415 269.970 ;
        RECT 222.605 269.800 222.775 269.970 ;
        RECT 225.715 269.800 225.885 269.970 ;
        RECT 226.075 269.800 226.245 269.970 ;
        RECT 5.295 266.090 5.465 266.260 ;
        RECT 5.655 266.090 5.825 266.260 ;
        RECT 6.015 266.090 6.185 266.260 ;
        RECT 6.375 266.090 6.545 266.260 ;
        RECT 6.735 266.090 6.905 266.260 ;
        RECT 7.095 266.090 7.265 266.260 ;
        RECT 7.455 266.090 7.625 266.260 ;
        RECT 7.815 266.090 7.985 266.260 ;
        RECT 8.175 266.090 8.345 266.260 ;
        RECT 8.535 266.090 8.705 266.260 ;
        RECT 8.895 266.090 9.065 266.260 ;
        RECT 9.255 266.090 9.425 266.260 ;
        RECT 9.615 266.090 9.785 266.260 ;
        RECT 9.975 266.090 10.145 266.260 ;
        RECT 10.335 266.090 10.505 266.260 ;
        RECT 10.695 266.090 10.865 266.260 ;
        RECT 11.055 266.090 11.225 266.260 ;
        RECT 11.415 266.090 11.585 266.260 ;
        RECT 11.775 266.090 11.945 266.260 ;
        RECT 12.135 266.090 12.305 266.260 ;
        RECT 18.635 266.070 18.805 266.240 ;
        RECT 18.995 266.070 19.165 266.240 ;
        RECT 19.355 266.070 19.525 266.240 ;
        RECT 19.715 266.070 19.885 266.240 ;
        RECT 20.075 266.070 20.245 266.240 ;
        RECT 20.435 266.070 20.605 266.240 ;
        RECT 20.795 266.070 20.965 266.240 ;
        RECT 21.155 266.070 21.325 266.240 ;
        RECT 21.515 266.070 21.685 266.240 ;
        RECT 21.875 266.070 22.045 266.240 ;
        RECT 22.235 266.070 22.405 266.240 ;
        RECT 22.595 266.070 22.765 266.240 ;
        RECT 22.955 266.070 23.125 266.240 ;
        RECT 23.315 266.070 23.485 266.240 ;
        RECT 23.675 266.070 23.845 266.240 ;
        RECT 24.035 266.070 24.205 266.240 ;
        RECT 24.395 266.070 24.565 266.240 ;
        RECT 24.755 266.070 24.925 266.240 ;
        RECT 25.115 266.070 25.285 266.240 ;
        RECT 25.475 266.070 25.645 266.240 ;
        RECT 32.005 266.100 32.175 266.270 ;
        RECT 32.365 266.100 32.535 266.270 ;
        RECT 32.725 266.100 32.895 266.270 ;
        RECT 33.085 266.100 33.255 266.270 ;
        RECT 33.445 266.100 33.615 266.270 ;
        RECT 33.805 266.100 33.975 266.270 ;
        RECT 34.165 266.100 34.335 266.270 ;
        RECT 34.525 266.100 34.695 266.270 ;
        RECT 34.885 266.100 35.055 266.270 ;
        RECT 35.245 266.100 35.415 266.270 ;
        RECT 35.605 266.100 35.775 266.270 ;
        RECT 35.965 266.100 36.135 266.270 ;
        RECT 36.325 266.100 36.495 266.270 ;
        RECT 36.685 266.100 36.855 266.270 ;
        RECT 37.045 266.100 37.215 266.270 ;
        RECT 37.405 266.100 37.575 266.270 ;
        RECT 37.765 266.100 37.935 266.270 ;
        RECT 38.125 266.100 38.295 266.270 ;
        RECT 38.485 266.100 38.655 266.270 ;
        RECT 38.845 266.100 39.015 266.270 ;
        RECT 45.235 266.100 45.405 266.270 ;
        RECT 45.595 266.100 45.765 266.270 ;
        RECT 45.955 266.100 46.125 266.270 ;
        RECT 46.315 266.100 46.485 266.270 ;
        RECT 46.675 266.100 46.845 266.270 ;
        RECT 47.035 266.100 47.205 266.270 ;
        RECT 47.395 266.100 47.565 266.270 ;
        RECT 47.755 266.100 47.925 266.270 ;
        RECT 48.115 266.100 48.285 266.270 ;
        RECT 48.475 266.100 48.645 266.270 ;
        RECT 48.835 266.100 49.005 266.270 ;
        RECT 49.195 266.100 49.365 266.270 ;
        RECT 49.555 266.100 49.725 266.270 ;
        RECT 49.915 266.100 50.085 266.270 ;
        RECT 50.275 266.100 50.445 266.270 ;
        RECT 50.635 266.100 50.805 266.270 ;
        RECT 50.995 266.100 51.165 266.270 ;
        RECT 51.355 266.100 51.525 266.270 ;
        RECT 51.715 266.100 51.885 266.270 ;
        RECT 52.075 266.100 52.245 266.270 ;
        RECT 58.505 266.070 58.675 266.240 ;
        RECT 58.865 266.070 59.035 266.240 ;
        RECT 59.225 266.070 59.395 266.240 ;
        RECT 59.585 266.070 59.755 266.240 ;
        RECT 59.945 266.070 60.115 266.240 ;
        RECT 60.305 266.070 60.475 266.240 ;
        RECT 60.665 266.070 60.835 266.240 ;
        RECT 61.025 266.070 61.195 266.240 ;
        RECT 61.385 266.070 61.555 266.240 ;
        RECT 61.745 266.070 61.915 266.240 ;
        RECT 62.105 266.070 62.275 266.240 ;
        RECT 62.465 266.070 62.635 266.240 ;
        RECT 62.825 266.070 62.995 266.240 ;
        RECT 63.185 266.070 63.355 266.240 ;
        RECT 63.545 266.070 63.715 266.240 ;
        RECT 63.905 266.070 64.075 266.240 ;
        RECT 64.265 266.070 64.435 266.240 ;
        RECT 64.625 266.070 64.795 266.240 ;
        RECT 64.985 266.070 65.155 266.240 ;
        RECT 65.345 266.070 65.515 266.240 ;
        RECT 71.775 266.100 71.945 266.270 ;
        RECT 72.135 266.100 72.305 266.270 ;
        RECT 72.495 266.100 72.665 266.270 ;
        RECT 72.855 266.100 73.025 266.270 ;
        RECT 73.215 266.100 73.385 266.270 ;
        RECT 73.575 266.100 73.745 266.270 ;
        RECT 73.935 266.100 74.105 266.270 ;
        RECT 74.295 266.100 74.465 266.270 ;
        RECT 74.655 266.100 74.825 266.270 ;
        RECT 75.015 266.100 75.185 266.270 ;
        RECT 75.375 266.100 75.545 266.270 ;
        RECT 75.735 266.100 75.905 266.270 ;
        RECT 76.095 266.100 76.265 266.270 ;
        RECT 76.455 266.100 76.625 266.270 ;
        RECT 76.815 266.100 76.985 266.270 ;
        RECT 77.175 266.100 77.345 266.270 ;
        RECT 77.535 266.100 77.705 266.270 ;
        RECT 77.895 266.100 78.065 266.270 ;
        RECT 78.255 266.100 78.425 266.270 ;
        RECT 78.615 266.100 78.785 266.270 ;
        RECT 84.905 266.120 85.075 266.290 ;
        RECT 85.265 266.120 85.435 266.290 ;
        RECT 85.625 266.120 85.795 266.290 ;
        RECT 85.985 266.120 86.155 266.290 ;
        RECT 86.345 266.120 86.515 266.290 ;
        RECT 86.705 266.120 86.875 266.290 ;
        RECT 87.065 266.120 87.235 266.290 ;
        RECT 87.425 266.120 87.595 266.290 ;
        RECT 87.785 266.120 87.955 266.290 ;
        RECT 88.145 266.120 88.315 266.290 ;
        RECT 88.505 266.120 88.675 266.290 ;
        RECT 88.865 266.120 89.035 266.290 ;
        RECT 89.225 266.120 89.395 266.290 ;
        RECT 89.585 266.120 89.755 266.290 ;
        RECT 89.945 266.120 90.115 266.290 ;
        RECT 90.305 266.120 90.475 266.290 ;
        RECT 90.665 266.120 90.835 266.290 ;
        RECT 91.025 266.120 91.195 266.290 ;
        RECT 91.385 266.120 91.555 266.290 ;
        RECT 91.745 266.120 91.915 266.290 ;
        RECT 97.820 265.915 102.310 266.445 ;
        RECT 97.885 264.760 98.055 264.930 ;
        RECT 98.245 264.760 98.415 264.930 ;
        RECT 101.355 264.760 101.525 264.930 ;
        RECT 101.715 264.760 101.885 264.930 ;
        RECT 4.855 264.510 5.025 264.680 ;
        RECT 5.215 264.510 5.385 264.680 ;
        RECT 8.325 264.510 8.495 264.680 ;
        RECT 8.685 264.510 8.855 264.680 ;
        RECT 11.795 264.510 11.965 264.680 ;
        RECT 12.155 264.510 12.325 264.680 ;
        RECT 18.195 264.490 18.365 264.660 ;
        RECT 18.555 264.490 18.725 264.660 ;
        RECT 21.665 264.490 21.835 264.660 ;
        RECT 22.025 264.490 22.195 264.660 ;
        RECT 25.135 264.490 25.305 264.660 ;
        RECT 25.495 264.490 25.665 264.660 ;
        RECT 31.565 264.520 31.735 264.690 ;
        RECT 31.925 264.520 32.095 264.690 ;
        RECT 35.035 264.520 35.205 264.690 ;
        RECT 35.395 264.520 35.565 264.690 ;
        RECT 38.505 264.520 38.675 264.690 ;
        RECT 38.865 264.520 39.035 264.690 ;
        RECT 44.795 264.520 44.965 264.690 ;
        RECT 45.155 264.520 45.325 264.690 ;
        RECT 48.265 264.520 48.435 264.690 ;
        RECT 48.625 264.520 48.795 264.690 ;
        RECT 51.735 264.520 51.905 264.690 ;
        RECT 52.095 264.520 52.265 264.690 ;
        RECT 58.065 264.490 58.235 264.660 ;
        RECT 58.425 264.490 58.595 264.660 ;
        RECT 61.535 264.490 61.705 264.660 ;
        RECT 61.895 264.490 62.065 264.660 ;
        RECT 65.005 264.490 65.175 264.660 ;
        RECT 65.365 264.490 65.535 264.660 ;
        RECT 71.335 264.520 71.505 264.690 ;
        RECT 71.695 264.520 71.865 264.690 ;
        RECT 74.805 264.520 74.975 264.690 ;
        RECT 75.165 264.520 75.335 264.690 ;
        RECT 78.275 264.520 78.445 264.690 ;
        RECT 78.635 264.520 78.805 264.690 ;
        RECT 84.465 264.540 84.635 264.710 ;
        RECT 84.825 264.540 84.995 264.710 ;
        RECT 87.935 264.540 88.105 264.710 ;
        RECT 88.295 264.540 88.465 264.710 ;
        RECT 91.405 264.540 91.575 264.710 ;
        RECT 91.765 264.540 91.935 264.710 ;
        RECT 4.855 261.220 5.025 261.390 ;
        RECT 5.215 261.220 5.385 261.390 ;
        RECT 8.325 261.220 8.495 261.390 ;
        RECT 8.685 261.220 8.855 261.390 ;
        RECT 11.795 261.220 11.965 261.390 ;
        RECT 12.155 261.220 12.325 261.390 ;
        RECT 4.855 257.930 5.025 258.100 ;
        RECT 5.215 257.930 5.385 258.100 ;
        RECT 8.325 257.930 8.495 258.100 ;
        RECT 8.685 257.930 8.855 258.100 ;
        RECT 11.795 257.930 11.965 258.100 ;
        RECT 12.155 257.930 12.325 258.100 ;
        RECT 4.855 254.640 5.025 254.810 ;
        RECT 5.215 254.640 5.385 254.810 ;
        RECT 8.325 254.640 8.495 254.810 ;
        RECT 8.685 254.640 8.855 254.810 ;
        RECT 11.795 254.640 11.965 254.810 ;
        RECT 12.155 254.640 12.325 254.810 ;
        RECT 4.855 251.350 5.025 251.520 ;
        RECT 5.215 251.350 5.385 251.520 ;
        RECT 8.325 251.350 8.495 251.520 ;
        RECT 8.685 251.350 8.855 251.520 ;
        RECT 11.795 251.350 11.965 251.520 ;
        RECT 12.155 251.350 12.325 251.520 ;
        RECT 4.855 248.060 5.025 248.230 ;
        RECT 5.215 248.060 5.385 248.230 ;
        RECT 8.325 248.060 8.495 248.230 ;
        RECT 8.685 248.060 8.855 248.230 ;
        RECT 11.795 248.060 11.965 248.230 ;
        RECT 12.155 248.060 12.325 248.230 ;
        RECT 18.195 261.200 18.365 261.370 ;
        RECT 18.555 261.200 18.725 261.370 ;
        RECT 21.665 261.200 21.835 261.370 ;
        RECT 22.025 261.200 22.195 261.370 ;
        RECT 25.135 261.200 25.305 261.370 ;
        RECT 25.495 261.200 25.665 261.370 ;
        RECT 18.195 257.910 18.365 258.080 ;
        RECT 18.555 257.910 18.725 258.080 ;
        RECT 21.665 257.910 21.835 258.080 ;
        RECT 22.025 257.910 22.195 258.080 ;
        RECT 25.135 257.910 25.305 258.080 ;
        RECT 25.495 257.910 25.665 258.080 ;
        RECT 18.195 254.620 18.365 254.790 ;
        RECT 18.555 254.620 18.725 254.790 ;
        RECT 21.665 254.620 21.835 254.790 ;
        RECT 22.025 254.620 22.195 254.790 ;
        RECT 25.135 254.620 25.305 254.790 ;
        RECT 25.495 254.620 25.665 254.790 ;
        RECT 18.195 251.330 18.365 251.500 ;
        RECT 18.555 251.330 18.725 251.500 ;
        RECT 21.665 251.330 21.835 251.500 ;
        RECT 22.025 251.330 22.195 251.500 ;
        RECT 25.135 251.330 25.305 251.500 ;
        RECT 25.495 251.330 25.665 251.500 ;
        RECT 18.195 248.040 18.365 248.210 ;
        RECT 18.555 248.040 18.725 248.210 ;
        RECT 21.665 248.040 21.835 248.210 ;
        RECT 22.025 248.040 22.195 248.210 ;
        RECT 25.135 248.040 25.305 248.210 ;
        RECT 25.495 248.040 25.665 248.210 ;
        RECT 4.855 244.770 5.025 244.940 ;
        RECT 5.215 244.770 5.385 244.940 ;
        RECT 8.325 244.770 8.495 244.940 ;
        RECT 8.685 244.770 8.855 244.940 ;
        RECT 11.795 244.770 11.965 244.940 ;
        RECT 12.155 244.770 12.325 244.940 ;
        RECT 4.855 241.480 5.025 241.650 ;
        RECT 5.215 241.480 5.385 241.650 ;
        RECT 8.325 241.480 8.495 241.650 ;
        RECT 8.685 241.480 8.855 241.650 ;
        RECT 11.795 241.480 11.965 241.650 ;
        RECT 12.155 241.480 12.325 241.650 ;
        RECT -46.120 236.805 -32.630 239.135 ;
        RECT 15.390 240.490 16.280 242.100 ;
        RECT 31.565 261.230 31.735 261.400 ;
        RECT 31.925 261.230 32.095 261.400 ;
        RECT 35.035 261.230 35.205 261.400 ;
        RECT 35.395 261.230 35.565 261.400 ;
        RECT 38.505 261.230 38.675 261.400 ;
        RECT 38.865 261.230 39.035 261.400 ;
        RECT 31.565 257.940 31.735 258.110 ;
        RECT 31.925 257.940 32.095 258.110 ;
        RECT 35.035 257.940 35.205 258.110 ;
        RECT 35.395 257.940 35.565 258.110 ;
        RECT 38.505 257.940 38.675 258.110 ;
        RECT 38.865 257.940 39.035 258.110 ;
        RECT 31.565 254.650 31.735 254.820 ;
        RECT 31.925 254.650 32.095 254.820 ;
        RECT 35.035 254.650 35.205 254.820 ;
        RECT 35.395 254.650 35.565 254.820 ;
        RECT 38.505 254.650 38.675 254.820 ;
        RECT 38.865 254.650 39.035 254.820 ;
        RECT 31.565 251.360 31.735 251.530 ;
        RECT 31.925 251.360 32.095 251.530 ;
        RECT 35.035 251.360 35.205 251.530 ;
        RECT 35.395 251.360 35.565 251.530 ;
        RECT 38.505 251.360 38.675 251.530 ;
        RECT 38.865 251.360 39.035 251.530 ;
        RECT 31.565 248.070 31.735 248.240 ;
        RECT 31.925 248.070 32.095 248.240 ;
        RECT 35.035 248.070 35.205 248.240 ;
        RECT 35.395 248.070 35.565 248.240 ;
        RECT 38.505 248.070 38.675 248.240 ;
        RECT 38.865 248.070 39.035 248.240 ;
        RECT 18.195 244.750 18.365 244.920 ;
        RECT 18.555 244.750 18.725 244.920 ;
        RECT 21.665 244.750 21.835 244.920 ;
        RECT 22.025 244.750 22.195 244.920 ;
        RECT 25.135 244.750 25.305 244.920 ;
        RECT 25.495 244.750 25.665 244.920 ;
        RECT 18.195 241.460 18.365 241.630 ;
        RECT 18.555 241.460 18.725 241.630 ;
        RECT 21.665 241.460 21.835 241.630 ;
        RECT 22.025 241.460 22.195 241.630 ;
        RECT 25.135 241.460 25.305 241.630 ;
        RECT 25.495 241.460 25.665 241.630 ;
        RECT 28.605 240.640 29.495 242.250 ;
        RECT 44.795 261.230 44.965 261.400 ;
        RECT 45.155 261.230 45.325 261.400 ;
        RECT 48.265 261.230 48.435 261.400 ;
        RECT 48.625 261.230 48.795 261.400 ;
        RECT 51.735 261.230 51.905 261.400 ;
        RECT 52.095 261.230 52.265 261.400 ;
        RECT 44.795 257.940 44.965 258.110 ;
        RECT 45.155 257.940 45.325 258.110 ;
        RECT 48.265 257.940 48.435 258.110 ;
        RECT 48.625 257.940 48.795 258.110 ;
        RECT 51.735 257.940 51.905 258.110 ;
        RECT 52.095 257.940 52.265 258.110 ;
        RECT 44.795 254.650 44.965 254.820 ;
        RECT 45.155 254.650 45.325 254.820 ;
        RECT 48.265 254.650 48.435 254.820 ;
        RECT 48.625 254.650 48.795 254.820 ;
        RECT 51.735 254.650 51.905 254.820 ;
        RECT 52.095 254.650 52.265 254.820 ;
        RECT 44.795 251.360 44.965 251.530 ;
        RECT 45.155 251.360 45.325 251.530 ;
        RECT 48.265 251.360 48.435 251.530 ;
        RECT 48.625 251.360 48.795 251.530 ;
        RECT 51.735 251.360 51.905 251.530 ;
        RECT 52.095 251.360 52.265 251.530 ;
        RECT 44.795 248.070 44.965 248.240 ;
        RECT 45.155 248.070 45.325 248.240 ;
        RECT 48.265 248.070 48.435 248.240 ;
        RECT 48.625 248.070 48.795 248.240 ;
        RECT 51.735 248.070 51.905 248.240 ;
        RECT 52.095 248.070 52.265 248.240 ;
        RECT 31.565 244.780 31.735 244.950 ;
        RECT 31.925 244.780 32.095 244.950 ;
        RECT 35.035 244.780 35.205 244.950 ;
        RECT 35.395 244.780 35.565 244.950 ;
        RECT 38.505 244.780 38.675 244.950 ;
        RECT 38.865 244.780 39.035 244.950 ;
        RECT 31.565 241.490 31.735 241.660 ;
        RECT 31.925 241.490 32.095 241.660 ;
        RECT 35.035 241.490 35.205 241.660 ;
        RECT 35.395 241.490 35.565 241.660 ;
        RECT 38.505 241.490 38.675 241.660 ;
        RECT 38.865 241.490 39.035 241.660 ;
        RECT 41.820 240.345 42.710 242.675 ;
        RECT 58.065 261.200 58.235 261.370 ;
        RECT 58.425 261.200 58.595 261.370 ;
        RECT 61.535 261.200 61.705 261.370 ;
        RECT 61.895 261.200 62.065 261.370 ;
        RECT 65.005 261.200 65.175 261.370 ;
        RECT 65.365 261.200 65.535 261.370 ;
        RECT 58.065 257.910 58.235 258.080 ;
        RECT 58.425 257.910 58.595 258.080 ;
        RECT 61.535 257.910 61.705 258.080 ;
        RECT 61.895 257.910 62.065 258.080 ;
        RECT 65.005 257.910 65.175 258.080 ;
        RECT 65.365 257.910 65.535 258.080 ;
        RECT 58.065 254.620 58.235 254.790 ;
        RECT 58.425 254.620 58.595 254.790 ;
        RECT 61.535 254.620 61.705 254.790 ;
        RECT 61.895 254.620 62.065 254.790 ;
        RECT 65.005 254.620 65.175 254.790 ;
        RECT 65.365 254.620 65.535 254.790 ;
        RECT 58.065 251.330 58.235 251.500 ;
        RECT 58.425 251.330 58.595 251.500 ;
        RECT 61.535 251.330 61.705 251.500 ;
        RECT 61.895 251.330 62.065 251.500 ;
        RECT 65.005 251.330 65.175 251.500 ;
        RECT 65.365 251.330 65.535 251.500 ;
        RECT 58.065 248.040 58.235 248.210 ;
        RECT 58.425 248.040 58.595 248.210 ;
        RECT 61.535 248.040 61.705 248.210 ;
        RECT 61.895 248.040 62.065 248.210 ;
        RECT 65.005 248.040 65.175 248.210 ;
        RECT 65.365 248.040 65.535 248.210 ;
        RECT 44.795 244.780 44.965 244.950 ;
        RECT 45.155 244.780 45.325 244.950 ;
        RECT 48.265 244.780 48.435 244.950 ;
        RECT 48.625 244.780 48.795 244.950 ;
        RECT 51.735 244.780 51.905 244.950 ;
        RECT 52.095 244.780 52.265 244.950 ;
        RECT 44.795 241.490 44.965 241.660 ;
        RECT 45.155 241.490 45.325 241.660 ;
        RECT 48.265 241.490 48.435 241.660 ;
        RECT 48.625 241.490 48.795 241.660 ;
        RECT 51.735 241.490 51.905 241.660 ;
        RECT 52.095 241.490 52.265 241.660 ;
        RECT 55.240 240.230 56.130 242.200 ;
        RECT 71.335 261.230 71.505 261.400 ;
        RECT 71.695 261.230 71.865 261.400 ;
        RECT 74.805 261.230 74.975 261.400 ;
        RECT 75.165 261.230 75.335 261.400 ;
        RECT 78.275 261.230 78.445 261.400 ;
        RECT 78.635 261.230 78.805 261.400 ;
        RECT 71.335 257.940 71.505 258.110 ;
        RECT 71.695 257.940 71.865 258.110 ;
        RECT 74.805 257.940 74.975 258.110 ;
        RECT 75.165 257.940 75.335 258.110 ;
        RECT 78.275 257.940 78.445 258.110 ;
        RECT 78.635 257.940 78.805 258.110 ;
        RECT 71.335 254.650 71.505 254.820 ;
        RECT 71.695 254.650 71.865 254.820 ;
        RECT 74.805 254.650 74.975 254.820 ;
        RECT 75.165 254.650 75.335 254.820 ;
        RECT 78.275 254.650 78.445 254.820 ;
        RECT 78.635 254.650 78.805 254.820 ;
        RECT 71.335 251.360 71.505 251.530 ;
        RECT 71.695 251.360 71.865 251.530 ;
        RECT 74.805 251.360 74.975 251.530 ;
        RECT 75.165 251.360 75.335 251.530 ;
        RECT 78.275 251.360 78.445 251.530 ;
        RECT 78.635 251.360 78.805 251.530 ;
        RECT 71.335 248.070 71.505 248.240 ;
        RECT 71.695 248.070 71.865 248.240 ;
        RECT 74.805 248.070 74.975 248.240 ;
        RECT 75.165 248.070 75.335 248.240 ;
        RECT 78.275 248.070 78.445 248.240 ;
        RECT 78.635 248.070 78.805 248.240 ;
        RECT 58.065 244.750 58.235 244.920 ;
        RECT 58.425 244.750 58.595 244.920 ;
        RECT 61.535 244.750 61.705 244.920 ;
        RECT 61.895 244.750 62.065 244.920 ;
        RECT 65.005 244.750 65.175 244.920 ;
        RECT 65.365 244.750 65.535 244.920 ;
        RECT 58.065 241.460 58.235 241.630 ;
        RECT 58.425 241.460 58.595 241.630 ;
        RECT 61.535 241.460 61.705 241.630 ;
        RECT 61.895 241.460 62.065 241.630 ;
        RECT 65.005 241.460 65.175 241.630 ;
        RECT 65.365 241.460 65.535 241.630 ;
        RECT 68.545 240.415 69.075 242.385 ;
        RECT 84.465 261.250 84.635 261.420 ;
        RECT 84.825 261.250 84.995 261.420 ;
        RECT 87.935 261.250 88.105 261.420 ;
        RECT 88.295 261.250 88.465 261.420 ;
        RECT 91.405 261.250 91.575 261.420 ;
        RECT 91.765 261.250 91.935 261.420 ;
        RECT 97.885 261.470 98.055 261.640 ;
        RECT 98.245 261.470 98.415 261.640 ;
        RECT 101.355 261.470 101.525 261.640 ;
        RECT 101.715 261.470 101.885 261.640 ;
        RECT 84.465 257.960 84.635 258.130 ;
        RECT 84.825 257.960 84.995 258.130 ;
        RECT 87.935 257.960 88.105 258.130 ;
        RECT 88.295 257.960 88.465 258.130 ;
        RECT 91.405 257.960 91.575 258.130 ;
        RECT 91.765 257.960 91.935 258.130 ;
        RECT 84.465 254.670 84.635 254.840 ;
        RECT 84.825 254.670 84.995 254.840 ;
        RECT 87.935 254.670 88.105 254.840 ;
        RECT 88.295 254.670 88.465 254.840 ;
        RECT 91.405 254.670 91.575 254.840 ;
        RECT 91.765 254.670 91.935 254.840 ;
        RECT 84.465 251.380 84.635 251.550 ;
        RECT 84.825 251.380 84.995 251.550 ;
        RECT 87.935 251.380 88.105 251.550 ;
        RECT 88.295 251.380 88.465 251.550 ;
        RECT 91.405 251.380 91.575 251.550 ;
        RECT 91.765 251.380 91.935 251.550 ;
        RECT 84.465 248.090 84.635 248.260 ;
        RECT 84.825 248.090 84.995 248.260 ;
        RECT 87.935 248.090 88.105 248.260 ;
        RECT 88.295 248.090 88.465 248.260 ;
        RECT 91.405 248.090 91.575 248.260 ;
        RECT 91.765 248.090 91.935 248.260 ;
        RECT 71.335 244.780 71.505 244.950 ;
        RECT 71.695 244.780 71.865 244.950 ;
        RECT 74.805 244.780 74.975 244.950 ;
        RECT 75.165 244.780 75.335 244.950 ;
        RECT 78.275 244.780 78.445 244.950 ;
        RECT 78.635 244.780 78.805 244.950 ;
        RECT 71.335 241.490 71.505 241.660 ;
        RECT 71.695 241.490 71.865 241.660 ;
        RECT 74.805 241.490 74.975 241.660 ;
        RECT 75.165 241.490 75.335 241.660 ;
        RECT 78.275 241.490 78.445 241.660 ;
        RECT 78.635 241.490 78.805 241.660 ;
        RECT 81.480 240.880 82.730 242.130 ;
        RECT 251.935 276.370 252.105 276.540 ;
        RECT 252.295 276.370 252.465 276.540 ;
        RECT 255.405 276.370 255.575 276.540 ;
        RECT 255.765 276.370 255.935 276.540 ;
        RECT 258.875 276.370 259.045 276.540 ;
        RECT 259.235 276.370 259.405 276.540 ;
        RECT 262.345 276.370 262.515 276.540 ;
        RECT 262.705 276.370 262.875 276.540 ;
        RECT 265.815 276.370 265.985 276.540 ;
        RECT 266.175 276.370 266.345 276.540 ;
        RECT 231.875 273.080 232.045 273.250 ;
        RECT 232.235 273.080 232.405 273.250 ;
        RECT 235.345 273.080 235.515 273.250 ;
        RECT 235.705 273.080 235.875 273.250 ;
        RECT 238.815 273.080 238.985 273.250 ;
        RECT 239.175 273.080 239.345 273.250 ;
        RECT 242.285 273.080 242.455 273.250 ;
        RECT 242.645 273.080 242.815 273.250 ;
        RECT 245.755 273.080 245.925 273.250 ;
        RECT 246.115 273.080 246.285 273.250 ;
        RECT 231.875 269.790 232.045 269.960 ;
        RECT 232.235 269.790 232.405 269.960 ;
        RECT 235.345 269.790 235.515 269.960 ;
        RECT 235.705 269.790 235.875 269.960 ;
        RECT 238.815 269.790 238.985 269.960 ;
        RECT 239.175 269.790 239.345 269.960 ;
        RECT 242.285 269.790 242.455 269.960 ;
        RECT 242.645 269.790 242.815 269.960 ;
        RECT 245.755 269.790 245.925 269.960 ;
        RECT 246.115 269.790 246.285 269.960 ;
        RECT 211.835 266.510 212.005 266.680 ;
        RECT 212.195 266.510 212.365 266.680 ;
        RECT 215.305 266.510 215.475 266.680 ;
        RECT 215.665 266.510 215.835 266.680 ;
        RECT 218.775 266.510 218.945 266.680 ;
        RECT 219.135 266.510 219.305 266.680 ;
        RECT 222.245 266.510 222.415 266.680 ;
        RECT 222.605 266.510 222.775 266.680 ;
        RECT 225.715 266.510 225.885 266.680 ;
        RECT 226.075 266.510 226.245 266.680 ;
        RECT 97.885 258.180 98.055 258.350 ;
        RECT 98.245 258.180 98.415 258.350 ;
        RECT 101.355 258.180 101.525 258.350 ;
        RECT 101.715 258.180 101.885 258.350 ;
        RECT 97.885 254.890 98.055 255.060 ;
        RECT 98.245 254.890 98.415 255.060 ;
        RECT 101.355 254.890 101.525 255.060 ;
        RECT 101.715 254.890 101.885 255.060 ;
        RECT 271.985 276.370 272.155 276.540 ;
        RECT 272.345 276.370 272.515 276.540 ;
        RECT 275.455 276.370 275.625 276.540 ;
        RECT 275.815 276.370 275.985 276.540 ;
        RECT 278.925 276.370 279.095 276.540 ;
        RECT 279.285 276.370 279.455 276.540 ;
        RECT 282.395 276.370 282.565 276.540 ;
        RECT 282.755 276.370 282.925 276.540 ;
        RECT 285.865 276.370 286.035 276.540 ;
        RECT 286.225 276.370 286.395 276.540 ;
        RECT 251.935 273.080 252.105 273.250 ;
        RECT 252.295 273.080 252.465 273.250 ;
        RECT 255.405 273.080 255.575 273.250 ;
        RECT 255.765 273.080 255.935 273.250 ;
        RECT 258.875 273.080 259.045 273.250 ;
        RECT 259.235 273.080 259.405 273.250 ;
        RECT 262.345 273.080 262.515 273.250 ;
        RECT 262.705 273.080 262.875 273.250 ;
        RECT 265.815 273.080 265.985 273.250 ;
        RECT 266.175 273.080 266.345 273.250 ;
        RECT 251.935 269.790 252.105 269.960 ;
        RECT 252.295 269.790 252.465 269.960 ;
        RECT 255.405 269.790 255.575 269.960 ;
        RECT 255.765 269.790 255.935 269.960 ;
        RECT 258.875 269.790 259.045 269.960 ;
        RECT 259.235 269.790 259.405 269.960 ;
        RECT 262.345 269.790 262.515 269.960 ;
        RECT 262.705 269.790 262.875 269.960 ;
        RECT 265.815 269.790 265.985 269.960 ;
        RECT 266.175 269.790 266.345 269.960 ;
        RECT 231.875 266.500 232.045 266.670 ;
        RECT 232.235 266.500 232.405 266.670 ;
        RECT 235.345 266.500 235.515 266.670 ;
        RECT 235.705 266.500 235.875 266.670 ;
        RECT 238.815 266.500 238.985 266.670 ;
        RECT 239.175 266.500 239.345 266.670 ;
        RECT 242.285 266.500 242.455 266.670 ;
        RECT 242.645 266.500 242.815 266.670 ;
        RECT 245.755 266.500 245.925 266.670 ;
        RECT 246.115 266.500 246.285 266.670 ;
        RECT 355.435 279.545 355.605 279.715 ;
        RECT 355.435 279.185 355.605 279.355 ;
        RECT 355.435 278.825 355.605 278.995 ;
        RECT 355.435 278.465 355.605 278.635 ;
        RECT 355.435 278.105 355.605 278.275 ;
        RECT 355.435 277.745 355.605 277.915 ;
        RECT 355.435 277.385 355.605 277.555 ;
        RECT 355.435 277.025 355.605 277.195 ;
        RECT 355.435 276.665 355.605 276.835 ;
        RECT 356.530 289.865 356.700 290.035 ;
        RECT 356.530 289.505 356.700 289.675 ;
        RECT 356.530 286.395 356.700 286.565 ;
        RECT 356.530 286.035 356.700 286.205 ;
        RECT 356.530 282.925 356.700 283.095 ;
        RECT 356.530 282.565 356.700 282.735 ;
        RECT 356.530 279.455 356.700 279.625 ;
        RECT 356.530 279.095 356.700 279.265 ;
        RECT 382.430 294.405 382.600 294.575 ;
        RECT 394.005 308.115 394.175 308.285 ;
        RECT 394.005 307.755 394.175 307.925 ;
        RECT 394.005 307.395 394.175 307.565 ;
        RECT 394.005 307.035 394.175 307.205 ;
        RECT 394.005 306.675 394.175 306.845 ;
        RECT 394.005 306.315 394.175 306.485 ;
        RECT 394.005 305.955 394.175 306.125 ;
        RECT 394.005 305.595 394.175 305.765 ;
        RECT 394.005 305.235 394.175 305.405 ;
        RECT 394.005 304.875 394.175 305.045 ;
        RECT 394.005 304.515 394.175 304.685 ;
        RECT 394.005 304.155 394.175 304.325 ;
        RECT 394.005 303.795 394.175 303.965 ;
        RECT 394.005 303.435 394.175 303.605 ;
        RECT 394.005 303.075 394.175 303.245 ;
        RECT 394.005 302.715 394.175 302.885 ;
        RECT 394.005 302.355 394.175 302.525 ;
        RECT 394.005 301.995 394.175 302.165 ;
        RECT 394.005 301.635 394.175 301.805 ;
        RECT 394.005 301.275 394.175 301.445 ;
        RECT 394.005 300.915 394.175 301.085 ;
        RECT 394.005 300.555 394.175 300.725 ;
        RECT 394.005 300.195 394.175 300.365 ;
        RECT 394.005 299.835 394.175 300.005 ;
        RECT 394.005 299.475 394.175 299.645 ;
        RECT 394.005 299.115 394.175 299.285 ;
        RECT 394.005 298.755 394.175 298.925 ;
        RECT 394.005 298.395 394.175 298.565 ;
        RECT 394.005 298.035 394.175 298.205 ;
        RECT 394.005 297.675 394.175 297.845 ;
        RECT 394.005 297.315 394.175 297.485 ;
        RECT 394.005 296.955 394.175 297.125 ;
        RECT 394.005 296.595 394.175 296.765 ;
        RECT 394.005 296.235 394.175 296.405 ;
        RECT 394.005 295.875 394.175 296.045 ;
        RECT 395.100 308.715 395.270 308.885 ;
        RECT 395.100 308.355 395.270 308.525 ;
        RECT 395.100 305.245 395.270 305.415 ;
        RECT 395.100 304.885 395.270 305.055 ;
        RECT 395.100 301.775 395.270 301.945 ;
        RECT 395.100 301.415 395.270 301.585 ;
        RECT 395.100 298.305 395.270 298.475 ;
        RECT 395.100 297.945 395.270 298.115 ;
        RECT 398.390 308.715 398.560 308.885 ;
        RECT 398.390 308.355 398.560 308.525 ;
        RECT 398.390 305.245 398.560 305.415 ;
        RECT 398.390 304.885 398.560 305.055 ;
        RECT 398.390 301.775 398.560 301.945 ;
        RECT 398.390 301.415 398.560 301.585 ;
        RECT 398.390 298.305 398.560 298.475 ;
        RECT 398.390 297.945 398.560 298.115 ;
        RECT 394.005 295.515 394.175 295.685 ;
        RECT 395.100 294.835 395.270 295.005 ;
        RECT 389.010 294.405 389.180 294.575 ;
        RECT 395.100 294.475 395.270 294.645 ;
        RECT 359.820 289.865 359.990 290.035 ;
        RECT 359.820 289.505 359.990 289.675 ;
        RECT 359.820 286.395 359.990 286.565 ;
        RECT 359.820 286.035 359.990 286.205 ;
        RECT 359.820 282.925 359.990 283.095 ;
        RECT 359.820 282.565 359.990 282.735 ;
        RECT 359.820 279.455 359.990 279.625 ;
        RECT 359.820 279.095 359.990 279.265 ;
        RECT 356.530 275.985 356.700 276.155 ;
        RECT 356.530 275.625 356.700 275.795 ;
        RECT 271.985 273.080 272.155 273.250 ;
        RECT 272.345 273.080 272.515 273.250 ;
        RECT 275.455 273.080 275.625 273.250 ;
        RECT 275.815 273.080 275.985 273.250 ;
        RECT 278.925 273.080 279.095 273.250 ;
        RECT 279.285 273.080 279.455 273.250 ;
        RECT 282.395 273.080 282.565 273.250 ;
        RECT 282.755 273.080 282.925 273.250 ;
        RECT 285.865 273.080 286.035 273.250 ;
        RECT 286.225 273.080 286.395 273.250 ;
        RECT 271.985 269.790 272.155 269.960 ;
        RECT 272.345 269.790 272.515 269.960 ;
        RECT 275.455 269.790 275.625 269.960 ;
        RECT 275.815 269.790 275.985 269.960 ;
        RECT 278.925 269.790 279.095 269.960 ;
        RECT 279.285 269.790 279.455 269.960 ;
        RECT 282.395 269.790 282.565 269.960 ;
        RECT 282.755 269.790 282.925 269.960 ;
        RECT 285.865 269.790 286.035 269.960 ;
        RECT 286.225 269.790 286.395 269.960 ;
        RECT 251.935 266.500 252.105 266.670 ;
        RECT 252.295 266.500 252.465 266.670 ;
        RECT 255.405 266.500 255.575 266.670 ;
        RECT 255.765 266.500 255.935 266.670 ;
        RECT 258.875 266.500 259.045 266.670 ;
        RECT 259.235 266.500 259.405 266.670 ;
        RECT 262.345 266.500 262.515 266.670 ;
        RECT 262.705 266.500 262.875 266.670 ;
        RECT 265.815 266.500 265.985 266.670 ;
        RECT 266.175 266.500 266.345 266.670 ;
        RECT 359.820 275.985 359.990 276.155 ;
        RECT 363.110 289.865 363.280 290.035 ;
        RECT 363.110 289.505 363.280 289.675 ;
        RECT 363.110 286.395 363.280 286.565 ;
        RECT 363.110 286.035 363.280 286.205 ;
        RECT 363.110 282.925 363.280 283.095 ;
        RECT 363.110 282.565 363.280 282.735 ;
        RECT 363.110 279.455 363.280 279.625 ;
        RECT 363.110 279.095 363.280 279.265 ;
        RECT 363.110 275.985 363.280 276.155 ;
        RECT 366.400 289.865 366.570 290.035 ;
        RECT 369.690 289.865 369.860 290.035 ;
        RECT 366.400 289.505 366.570 289.675 ;
        RECT 366.400 286.395 366.570 286.565 ;
        RECT 366.400 286.035 366.570 286.205 ;
        RECT 366.400 282.925 366.570 283.095 ;
        RECT 366.400 282.565 366.570 282.735 ;
        RECT 366.400 279.455 366.570 279.625 ;
        RECT 366.400 279.095 366.570 279.265 ;
        RECT 366.400 275.985 366.570 276.155 ;
        RECT 369.690 289.505 369.860 289.675 ;
        RECT 369.690 286.395 369.860 286.565 ;
        RECT 369.690 286.035 369.860 286.205 ;
        RECT 369.690 282.925 369.860 283.095 ;
        RECT 369.690 282.565 369.860 282.735 ;
        RECT 369.690 279.455 369.860 279.625 ;
        RECT 369.690 279.095 369.860 279.265 ;
        RECT 359.820 275.625 359.990 275.795 ;
        RECT 363.110 275.625 363.280 275.795 ;
        RECT 366.400 275.625 366.570 275.795 ;
        RECT 369.690 275.985 369.860 276.155 ;
        RECT 374.755 289.165 374.925 289.335 ;
        RECT 374.755 288.805 374.925 288.975 ;
        RECT 374.755 288.445 374.925 288.615 ;
        RECT 374.755 288.085 374.925 288.255 ;
        RECT 374.755 287.725 374.925 287.895 ;
        RECT 374.755 287.365 374.925 287.535 ;
        RECT 374.755 287.005 374.925 287.175 ;
        RECT 374.755 286.645 374.925 286.815 ;
        RECT 374.755 286.285 374.925 286.455 ;
        RECT 374.755 285.925 374.925 286.095 ;
        RECT 374.755 285.565 374.925 285.735 ;
        RECT 374.755 285.205 374.925 285.375 ;
        RECT 374.755 284.845 374.925 285.015 ;
        RECT 374.755 284.485 374.925 284.655 ;
        RECT 374.755 284.125 374.925 284.295 ;
        RECT 374.755 283.765 374.925 283.935 ;
        RECT 374.755 283.405 374.925 283.575 ;
        RECT 374.755 283.045 374.925 283.215 ;
        RECT 374.755 282.685 374.925 282.855 ;
        RECT 374.755 282.325 374.925 282.495 ;
        RECT 374.755 281.965 374.925 282.135 ;
        RECT 374.755 281.605 374.925 281.775 ;
        RECT 374.755 281.245 374.925 281.415 ;
        RECT 374.755 280.885 374.925 281.055 ;
        RECT 374.755 280.525 374.925 280.695 ;
        RECT 374.755 280.165 374.925 280.335 ;
        RECT 374.755 279.805 374.925 279.975 ;
        RECT 374.755 279.445 374.925 279.615 ;
        RECT 374.755 279.085 374.925 279.255 ;
        RECT 374.755 278.725 374.925 278.895 ;
        RECT 374.755 278.365 374.925 278.535 ;
        RECT 374.755 278.005 374.925 278.175 ;
        RECT 374.755 277.645 374.925 277.815 ;
        RECT 374.755 277.285 374.925 277.455 ;
        RECT 374.755 276.925 374.925 277.095 ;
        RECT 374.755 276.565 374.925 276.735 ;
        RECT 375.850 289.765 376.020 289.935 ;
        RECT 375.850 289.405 376.020 289.575 ;
        RECT 375.850 286.295 376.020 286.465 ;
        RECT 375.850 285.935 376.020 286.105 ;
        RECT 375.850 282.825 376.020 282.995 ;
        RECT 375.850 282.465 376.020 282.635 ;
        RECT 375.850 279.355 376.020 279.525 ;
        RECT 375.850 278.995 376.020 279.165 ;
        RECT 382.430 289.765 382.600 289.935 ;
        RECT 398.390 294.835 398.560 295.005 ;
        RECT 401.680 308.715 401.850 308.885 ;
        RECT 401.680 308.355 401.850 308.525 ;
        RECT 401.680 305.245 401.850 305.415 ;
        RECT 401.680 304.885 401.850 305.055 ;
        RECT 401.680 301.775 401.850 301.945 ;
        RECT 401.680 301.415 401.850 301.585 ;
        RECT 401.680 298.305 401.850 298.475 ;
        RECT 401.680 297.945 401.850 298.115 ;
        RECT 401.680 294.835 401.850 295.005 ;
        RECT 404.970 308.715 405.140 308.885 ;
        RECT 408.260 308.715 408.430 308.885 ;
        RECT 404.970 308.355 405.140 308.525 ;
        RECT 404.970 305.245 405.140 305.415 ;
        RECT 404.970 304.885 405.140 305.055 ;
        RECT 404.970 301.775 405.140 301.945 ;
        RECT 404.970 301.415 405.140 301.585 ;
        RECT 404.970 298.305 405.140 298.475 ;
        RECT 404.970 297.945 405.140 298.115 ;
        RECT 404.970 294.835 405.140 295.005 ;
        RECT 408.260 308.355 408.430 308.525 ;
        RECT 796.635 308.015 796.805 308.185 ;
        RECT 797.115 308.015 797.285 308.185 ;
        RECT 797.595 308.015 797.765 308.185 ;
        RECT 798.075 308.015 798.245 308.185 ;
        RECT 798.555 308.015 798.725 308.185 ;
        RECT 799.035 308.015 799.205 308.185 ;
        RECT 799.515 308.015 799.685 308.185 ;
        RECT 799.995 308.015 800.165 308.185 ;
        RECT 800.475 308.015 800.645 308.185 ;
        RECT 800.955 308.015 801.125 308.185 ;
        RECT 801.435 308.015 801.605 308.185 ;
        RECT 801.915 308.015 802.085 308.185 ;
        RECT 802.395 308.015 802.565 308.185 ;
        RECT 802.875 308.015 803.045 308.185 ;
        RECT 803.355 308.015 803.525 308.185 ;
        RECT 803.835 308.015 804.005 308.185 ;
        RECT 804.315 308.015 804.485 308.185 ;
        RECT 804.795 308.015 804.965 308.185 ;
        RECT 805.275 308.015 805.445 308.185 ;
        RECT 805.755 308.015 805.925 308.185 ;
        RECT 806.235 308.015 806.405 308.185 ;
        RECT 806.715 308.015 806.885 308.185 ;
        RECT 807.195 308.015 807.365 308.185 ;
        RECT 807.675 308.015 807.845 308.185 ;
        RECT 808.155 308.015 808.325 308.185 ;
        RECT 808.635 308.015 808.805 308.185 ;
        RECT 809.115 308.015 809.285 308.185 ;
        RECT 809.595 308.015 809.765 308.185 ;
        RECT 810.075 308.015 810.245 308.185 ;
        RECT 810.555 308.015 810.725 308.185 ;
        RECT 811.035 308.015 811.205 308.185 ;
        RECT 811.515 308.015 811.685 308.185 ;
        RECT 797.140 307.535 797.310 307.705 ;
        RECT 797.500 307.535 797.670 307.705 ;
        RECT 799.530 307.535 799.700 307.705 ;
        RECT 801.960 307.535 802.130 307.705 ;
        RECT 802.320 307.535 802.490 307.705 ;
        RECT 802.680 307.535 802.850 307.705 ;
        RECT 804.300 307.535 804.470 307.705 ;
        RECT 804.660 307.535 804.830 307.705 ;
        RECT 805.020 307.535 805.190 307.705 ;
        RECT 806.995 307.535 807.165 307.705 ;
        RECT 807.355 307.535 807.525 307.705 ;
        RECT 807.715 307.535 807.885 307.705 ;
        RECT 808.750 307.535 808.920 307.705 ;
        RECT 809.110 307.535 809.280 307.705 ;
        RECT 809.470 307.535 809.640 307.705 ;
        RECT 810.280 307.535 810.450 307.705 ;
        RECT 810.640 307.535 810.810 307.705 ;
        RECT 811.000 307.535 811.170 307.705 ;
        RECT 814.395 308.015 814.565 308.185 ;
        RECT 814.875 308.015 815.045 308.185 ;
        RECT 815.355 308.015 815.525 308.185 ;
        RECT 815.835 308.015 816.005 308.185 ;
        RECT 816.315 308.015 816.485 308.185 ;
        RECT 816.795 308.015 816.965 308.185 ;
        RECT 817.275 308.015 817.445 308.185 ;
        RECT 817.755 308.015 817.925 308.185 ;
        RECT 818.235 308.015 818.405 308.185 ;
        RECT 818.715 308.015 818.885 308.185 ;
        RECT 819.195 308.015 819.365 308.185 ;
        RECT 819.675 308.015 819.845 308.185 ;
        RECT 820.155 308.015 820.325 308.185 ;
        RECT 820.635 308.015 820.805 308.185 ;
        RECT 821.115 308.015 821.285 308.185 ;
        RECT 821.595 308.015 821.765 308.185 ;
        RECT 822.075 308.015 822.245 308.185 ;
        RECT 822.555 308.015 822.725 308.185 ;
        RECT 823.035 308.015 823.205 308.185 ;
        RECT 823.515 308.015 823.685 308.185 ;
        RECT 823.995 308.015 824.165 308.185 ;
        RECT 824.475 308.015 824.645 308.185 ;
        RECT 824.955 308.015 825.125 308.185 ;
        RECT 825.435 308.015 825.605 308.185 ;
        RECT 825.915 308.015 826.085 308.185 ;
        RECT 826.395 308.015 826.565 308.185 ;
        RECT 826.875 308.015 827.045 308.185 ;
        RECT 827.355 308.015 827.525 308.185 ;
        RECT 827.835 308.015 828.005 308.185 ;
        RECT 828.315 308.015 828.485 308.185 ;
        RECT 828.795 308.015 828.965 308.185 ;
        RECT 829.275 308.015 829.445 308.185 ;
        RECT 814.900 307.535 815.070 307.705 ;
        RECT 815.260 307.535 815.430 307.705 ;
        RECT 817.290 307.535 817.460 307.705 ;
        RECT 819.720 307.535 819.890 307.705 ;
        RECT 820.080 307.535 820.250 307.705 ;
        RECT 820.440 307.535 820.610 307.705 ;
        RECT 822.060 307.535 822.230 307.705 ;
        RECT 822.420 307.535 822.590 307.705 ;
        RECT 822.780 307.535 822.950 307.705 ;
        RECT 824.755 307.535 824.925 307.705 ;
        RECT 825.115 307.535 825.285 307.705 ;
        RECT 825.475 307.535 825.645 307.705 ;
        RECT 826.510 307.535 826.680 307.705 ;
        RECT 826.870 307.535 827.040 307.705 ;
        RECT 827.230 307.535 827.400 307.705 ;
        RECT 828.040 307.535 828.210 307.705 ;
        RECT 828.400 307.535 828.570 307.705 ;
        RECT 828.760 307.535 828.930 307.705 ;
        RECT 831.935 307.985 832.105 308.155 ;
        RECT 832.415 307.985 832.585 308.155 ;
        RECT 832.895 307.985 833.065 308.155 ;
        RECT 835.575 308.045 835.745 308.215 ;
        RECT 836.055 308.045 836.225 308.215 ;
        RECT 836.535 308.045 836.705 308.215 ;
        RECT 837.015 308.045 837.185 308.215 ;
        RECT 837.495 308.045 837.665 308.215 ;
        RECT 837.975 308.045 838.145 308.215 ;
        RECT 838.455 308.045 838.625 308.215 ;
        RECT 838.935 308.045 839.105 308.215 ;
        RECT 839.415 308.045 839.585 308.215 ;
        RECT 839.895 308.045 840.065 308.215 ;
        RECT 840.375 308.045 840.545 308.215 ;
        RECT 831.900 307.505 832.070 307.675 ;
        RECT 832.260 307.505 832.430 307.675 ;
        RECT 835.980 307.565 836.150 307.735 ;
        RECT 836.340 307.565 836.510 307.735 ;
        RECT 836.700 307.565 836.870 307.735 ;
        RECT 837.060 307.565 837.230 307.735 ;
        RECT 837.420 307.565 837.590 307.735 ;
        RECT 837.780 307.565 837.950 307.735 ;
        RECT 838.505 307.565 838.675 307.735 ;
        RECT 838.865 307.565 839.035 307.735 ;
        RECT 839.225 307.565 839.395 307.735 ;
        RECT 839.585 307.565 839.755 307.735 ;
        RECT 839.945 307.565 840.115 307.735 ;
        RECT 842.845 308.045 843.015 308.215 ;
        RECT 843.325 308.045 843.495 308.215 ;
        RECT 843.805 308.045 843.975 308.215 ;
        RECT 842.810 307.565 842.980 307.735 ;
        RECT 843.170 307.565 843.340 307.735 ;
        RECT 408.260 305.245 408.430 305.415 ;
        RECT 408.260 304.885 408.430 305.055 ;
        RECT 408.260 301.775 408.430 301.945 ;
        RECT 408.260 301.415 408.430 301.585 ;
        RECT 680.215 298.955 680.385 299.125 ;
        RECT 680.695 298.955 680.865 299.125 ;
        RECT 681.175 298.955 681.345 299.125 ;
        RECT 681.655 298.955 681.825 299.125 ;
        RECT 682.135 298.955 682.305 299.125 ;
        RECT 682.615 298.955 682.785 299.125 ;
        RECT 683.095 298.955 683.265 299.125 ;
        RECT 683.575 298.955 683.745 299.125 ;
        RECT 684.055 298.955 684.225 299.125 ;
        RECT 684.535 298.955 684.705 299.125 ;
        RECT 685.015 298.955 685.185 299.125 ;
        RECT 685.495 298.955 685.665 299.125 ;
        RECT 685.975 298.955 686.145 299.125 ;
        RECT 686.455 298.955 686.625 299.125 ;
        RECT 686.935 298.955 687.105 299.125 ;
        RECT 687.415 298.955 687.585 299.125 ;
        RECT 687.895 298.955 688.065 299.125 ;
        RECT 688.375 298.955 688.545 299.125 ;
        RECT 688.855 298.955 689.025 299.125 ;
        RECT 689.335 298.955 689.505 299.125 ;
        RECT 689.815 298.955 689.985 299.125 ;
        RECT 690.295 298.955 690.465 299.125 ;
        RECT 690.775 298.955 690.945 299.125 ;
        RECT 691.255 298.955 691.425 299.125 ;
        RECT 691.735 298.955 691.905 299.125 ;
        RECT 692.215 298.955 692.385 299.125 ;
        RECT 692.695 298.955 692.865 299.125 ;
        RECT 693.175 298.955 693.345 299.125 ;
        RECT 693.655 298.955 693.825 299.125 ;
        RECT 694.135 298.955 694.305 299.125 ;
        RECT 694.615 298.955 694.785 299.125 ;
        RECT 695.095 298.955 695.265 299.125 ;
        RECT 408.260 298.305 408.430 298.475 ;
        RECT 408.260 297.945 408.430 298.115 ;
        RECT 680.720 298.475 680.890 298.645 ;
        RECT 681.080 298.475 681.250 298.645 ;
        RECT 683.110 298.475 683.280 298.645 ;
        RECT 685.540 298.475 685.710 298.645 ;
        RECT 685.900 298.475 686.070 298.645 ;
        RECT 686.260 298.475 686.430 298.645 ;
        RECT 687.880 298.475 688.050 298.645 ;
        RECT 688.240 298.475 688.410 298.645 ;
        RECT 688.600 298.475 688.770 298.645 ;
        RECT 690.575 298.475 690.745 298.645 ;
        RECT 690.935 298.475 691.105 298.645 ;
        RECT 691.295 298.475 691.465 298.645 ;
        RECT 692.330 298.475 692.500 298.645 ;
        RECT 692.690 298.475 692.860 298.645 ;
        RECT 693.050 298.475 693.220 298.645 ;
        RECT 693.860 298.475 694.030 298.645 ;
        RECT 694.220 298.475 694.390 298.645 ;
        RECT 694.580 298.475 694.750 298.645 ;
        RECT 697.705 298.915 697.875 299.085 ;
        RECT 698.185 298.915 698.355 299.085 ;
        RECT 698.665 298.915 698.835 299.085 ;
        RECT 699.145 298.915 699.315 299.085 ;
        RECT 699.625 298.915 699.795 299.085 ;
        RECT 700.105 298.915 700.275 299.085 ;
        RECT 700.585 298.915 700.755 299.085 ;
        RECT 701.065 298.915 701.235 299.085 ;
        RECT 701.545 298.915 701.715 299.085 ;
        RECT 702.025 298.915 702.195 299.085 ;
        RECT 702.505 298.915 702.675 299.085 ;
        RECT 702.985 298.915 703.155 299.085 ;
        RECT 703.465 298.915 703.635 299.085 ;
        RECT 703.945 298.915 704.115 299.085 ;
        RECT 704.425 298.915 704.595 299.085 ;
        RECT 704.905 298.915 705.075 299.085 ;
        RECT 705.385 298.915 705.555 299.085 ;
        RECT 705.865 298.915 706.035 299.085 ;
        RECT 706.345 298.915 706.515 299.085 ;
        RECT 706.825 298.915 706.995 299.085 ;
        RECT 707.305 298.915 707.475 299.085 ;
        RECT 707.785 298.915 707.955 299.085 ;
        RECT 708.265 298.915 708.435 299.085 ;
        RECT 708.745 298.915 708.915 299.085 ;
        RECT 709.225 298.915 709.395 299.085 ;
        RECT 709.705 298.915 709.875 299.085 ;
        RECT 710.185 298.915 710.355 299.085 ;
        RECT 710.665 298.915 710.835 299.085 ;
        RECT 711.145 298.915 711.315 299.085 ;
        RECT 711.625 298.915 711.795 299.085 ;
        RECT 712.105 298.915 712.275 299.085 ;
        RECT 712.585 298.915 712.755 299.085 ;
        RECT 698.210 298.435 698.380 298.605 ;
        RECT 698.570 298.435 698.740 298.605 ;
        RECT 700.600 298.435 700.770 298.605 ;
        RECT 703.030 298.435 703.200 298.605 ;
        RECT 703.390 298.435 703.560 298.605 ;
        RECT 703.750 298.435 703.920 298.605 ;
        RECT 705.370 298.435 705.540 298.605 ;
        RECT 705.730 298.435 705.900 298.605 ;
        RECT 706.090 298.435 706.260 298.605 ;
        RECT 708.065 298.435 708.235 298.605 ;
        RECT 708.425 298.435 708.595 298.605 ;
        RECT 708.785 298.435 708.955 298.605 ;
        RECT 709.820 298.435 709.990 298.605 ;
        RECT 710.180 298.435 710.350 298.605 ;
        RECT 710.540 298.435 710.710 298.605 ;
        RECT 711.350 298.435 711.520 298.605 ;
        RECT 711.710 298.435 711.880 298.605 ;
        RECT 712.070 298.435 712.240 298.605 ;
        RECT 715.315 298.975 715.485 299.145 ;
        RECT 715.795 298.975 715.965 299.145 ;
        RECT 716.275 298.975 716.445 299.145 ;
        RECT 716.755 298.975 716.925 299.145 ;
        RECT 717.235 298.975 717.405 299.145 ;
        RECT 717.715 298.975 717.885 299.145 ;
        RECT 718.195 298.975 718.365 299.145 ;
        RECT 718.675 298.975 718.845 299.145 ;
        RECT 719.155 298.975 719.325 299.145 ;
        RECT 719.635 298.975 719.805 299.145 ;
        RECT 720.115 298.975 720.285 299.145 ;
        RECT 720.595 298.975 720.765 299.145 ;
        RECT 721.075 298.975 721.245 299.145 ;
        RECT 721.555 298.975 721.725 299.145 ;
        RECT 722.035 298.975 722.205 299.145 ;
        RECT 722.515 298.975 722.685 299.145 ;
        RECT 722.995 298.975 723.165 299.145 ;
        RECT 723.475 298.975 723.645 299.145 ;
        RECT 723.955 298.975 724.125 299.145 ;
        RECT 724.435 298.975 724.605 299.145 ;
        RECT 724.915 298.975 725.085 299.145 ;
        RECT 725.395 298.975 725.565 299.145 ;
        RECT 725.875 298.975 726.045 299.145 ;
        RECT 726.355 298.975 726.525 299.145 ;
        RECT 726.835 298.975 727.005 299.145 ;
        RECT 727.315 298.975 727.485 299.145 ;
        RECT 727.795 298.975 727.965 299.145 ;
        RECT 728.275 298.975 728.445 299.145 ;
        RECT 728.755 298.975 728.925 299.145 ;
        RECT 729.235 298.975 729.405 299.145 ;
        RECT 729.715 298.975 729.885 299.145 ;
        RECT 730.195 298.975 730.365 299.145 ;
        RECT 715.820 298.495 715.990 298.665 ;
        RECT 716.180 298.495 716.350 298.665 ;
        RECT 718.210 298.495 718.380 298.665 ;
        RECT 720.640 298.495 720.810 298.665 ;
        RECT 721.000 298.495 721.170 298.665 ;
        RECT 721.360 298.495 721.530 298.665 ;
        RECT 722.980 298.495 723.150 298.665 ;
        RECT 723.340 298.495 723.510 298.665 ;
        RECT 723.700 298.495 723.870 298.665 ;
        RECT 725.675 298.495 725.845 298.665 ;
        RECT 726.035 298.495 726.205 298.665 ;
        RECT 726.395 298.495 726.565 298.665 ;
        RECT 727.430 298.495 727.600 298.665 ;
        RECT 727.790 298.495 727.960 298.665 ;
        RECT 728.150 298.495 728.320 298.665 ;
        RECT 728.960 298.495 729.130 298.665 ;
        RECT 729.320 298.495 729.490 298.665 ;
        RECT 729.680 298.495 729.850 298.665 ;
        RECT 733.015 298.925 733.185 299.095 ;
        RECT 733.495 298.925 733.665 299.095 ;
        RECT 733.975 298.925 734.145 299.095 ;
        RECT 734.455 298.925 734.625 299.095 ;
        RECT 734.935 298.925 735.105 299.095 ;
        RECT 735.415 298.925 735.585 299.095 ;
        RECT 735.895 298.925 736.065 299.095 ;
        RECT 736.375 298.925 736.545 299.095 ;
        RECT 736.855 298.925 737.025 299.095 ;
        RECT 737.335 298.925 737.505 299.095 ;
        RECT 737.815 298.925 737.985 299.095 ;
        RECT 738.295 298.925 738.465 299.095 ;
        RECT 738.775 298.925 738.945 299.095 ;
        RECT 739.255 298.925 739.425 299.095 ;
        RECT 739.735 298.925 739.905 299.095 ;
        RECT 740.215 298.925 740.385 299.095 ;
        RECT 740.695 298.925 740.865 299.095 ;
        RECT 741.175 298.925 741.345 299.095 ;
        RECT 741.655 298.925 741.825 299.095 ;
        RECT 742.135 298.925 742.305 299.095 ;
        RECT 742.615 298.925 742.785 299.095 ;
        RECT 743.095 298.925 743.265 299.095 ;
        RECT 743.575 298.925 743.745 299.095 ;
        RECT 744.055 298.925 744.225 299.095 ;
        RECT 744.535 298.925 744.705 299.095 ;
        RECT 745.015 298.925 745.185 299.095 ;
        RECT 745.495 298.925 745.665 299.095 ;
        RECT 745.975 298.925 746.145 299.095 ;
        RECT 746.455 298.925 746.625 299.095 ;
        RECT 746.935 298.925 747.105 299.095 ;
        RECT 747.415 298.925 747.585 299.095 ;
        RECT 747.895 298.925 748.065 299.095 ;
        RECT 733.520 298.445 733.690 298.615 ;
        RECT 733.880 298.445 734.050 298.615 ;
        RECT 735.910 298.445 736.080 298.615 ;
        RECT 738.340 298.445 738.510 298.615 ;
        RECT 738.700 298.445 738.870 298.615 ;
        RECT 739.060 298.445 739.230 298.615 ;
        RECT 740.680 298.445 740.850 298.615 ;
        RECT 741.040 298.445 741.210 298.615 ;
        RECT 741.400 298.445 741.570 298.615 ;
        RECT 743.375 298.445 743.545 298.615 ;
        RECT 743.735 298.445 743.905 298.615 ;
        RECT 744.095 298.445 744.265 298.615 ;
        RECT 745.130 298.445 745.300 298.615 ;
        RECT 745.490 298.445 745.660 298.615 ;
        RECT 745.850 298.445 746.020 298.615 ;
        RECT 746.660 298.445 746.830 298.615 ;
        RECT 747.020 298.445 747.190 298.615 ;
        RECT 747.380 298.445 747.550 298.615 ;
        RECT 750.755 298.915 750.925 299.085 ;
        RECT 751.235 298.915 751.405 299.085 ;
        RECT 751.715 298.915 751.885 299.085 ;
        RECT 752.195 298.915 752.365 299.085 ;
        RECT 752.675 298.915 752.845 299.085 ;
        RECT 753.155 298.915 753.325 299.085 ;
        RECT 753.635 298.915 753.805 299.085 ;
        RECT 754.115 298.915 754.285 299.085 ;
        RECT 754.595 298.915 754.765 299.085 ;
        RECT 755.075 298.915 755.245 299.085 ;
        RECT 755.555 298.915 755.725 299.085 ;
        RECT 756.035 298.915 756.205 299.085 ;
        RECT 756.515 298.915 756.685 299.085 ;
        RECT 756.995 298.915 757.165 299.085 ;
        RECT 757.475 298.915 757.645 299.085 ;
        RECT 757.955 298.915 758.125 299.085 ;
        RECT 758.435 298.915 758.605 299.085 ;
        RECT 758.915 298.915 759.085 299.085 ;
        RECT 759.395 298.915 759.565 299.085 ;
        RECT 759.875 298.915 760.045 299.085 ;
        RECT 760.355 298.915 760.525 299.085 ;
        RECT 760.835 298.915 761.005 299.085 ;
        RECT 761.315 298.915 761.485 299.085 ;
        RECT 761.795 298.915 761.965 299.085 ;
        RECT 762.275 298.915 762.445 299.085 ;
        RECT 762.755 298.915 762.925 299.085 ;
        RECT 763.235 298.915 763.405 299.085 ;
        RECT 763.715 298.915 763.885 299.085 ;
        RECT 764.195 298.915 764.365 299.085 ;
        RECT 764.675 298.915 764.845 299.085 ;
        RECT 765.155 298.915 765.325 299.085 ;
        RECT 765.635 298.915 765.805 299.085 ;
        RECT 751.260 298.435 751.430 298.605 ;
        RECT 751.620 298.435 751.790 298.605 ;
        RECT 753.650 298.435 753.820 298.605 ;
        RECT 756.080 298.435 756.250 298.605 ;
        RECT 756.440 298.435 756.610 298.605 ;
        RECT 756.800 298.435 756.970 298.605 ;
        RECT 758.420 298.435 758.590 298.605 ;
        RECT 758.780 298.435 758.950 298.605 ;
        RECT 759.140 298.435 759.310 298.605 ;
        RECT 761.115 298.435 761.285 298.605 ;
        RECT 761.475 298.435 761.645 298.605 ;
        RECT 761.835 298.435 762.005 298.605 ;
        RECT 762.870 298.435 763.040 298.605 ;
        RECT 763.230 298.435 763.400 298.605 ;
        RECT 763.590 298.435 763.760 298.605 ;
        RECT 764.400 298.435 764.570 298.605 ;
        RECT 764.760 298.435 764.930 298.605 ;
        RECT 765.120 298.435 765.290 298.605 ;
        RECT 855.955 298.275 856.125 298.445 ;
        RECT 856.435 298.275 856.605 298.445 ;
        RECT 856.915 298.275 857.085 298.445 ;
        RECT 857.395 298.275 857.565 298.445 ;
        RECT 857.875 298.275 858.045 298.445 ;
        RECT 858.355 298.275 858.525 298.445 ;
        RECT 858.835 298.275 859.005 298.445 ;
        RECT 855.910 297.795 856.080 297.965 ;
        RECT 856.270 297.795 856.440 297.965 ;
        RECT 856.630 297.795 856.800 297.965 ;
        RECT 857.350 297.795 857.520 297.965 ;
        RECT 857.710 297.795 857.880 297.965 ;
        RECT 858.070 297.795 858.240 297.965 ;
        RECT 858.430 297.795 858.600 297.965 ;
        RECT 839.545 296.295 839.715 296.465 ;
        RECT 840.025 296.295 840.195 296.465 ;
        RECT 840.505 296.295 840.675 296.465 ;
        RECT 840.985 296.295 841.155 296.465 ;
        RECT 841.465 296.295 841.635 296.465 ;
        RECT 841.945 296.295 842.115 296.465 ;
        RECT 842.425 296.295 842.595 296.465 ;
        RECT 839.500 295.815 839.670 295.985 ;
        RECT 839.860 295.815 840.030 295.985 ;
        RECT 840.220 295.815 840.390 295.985 ;
        RECT 398.390 294.475 398.560 294.645 ;
        RECT 401.680 294.475 401.850 294.645 ;
        RECT 404.970 294.475 405.140 294.645 ;
        RECT 408.260 294.835 408.430 295.005 ;
        RECT 408.260 294.475 408.430 294.645 ;
        RECT 601.250 294.815 601.420 294.985 ;
        RECT 602.430 294.825 602.600 294.995 ;
        RECT 604.010 294.825 604.180 294.995 ;
        RECT 605.590 294.825 605.760 294.995 ;
        RECT 606.950 294.835 607.120 295.005 ;
        RECT 608.530 294.835 608.700 295.005 ;
        RECT 610.110 294.835 610.280 295.005 ;
        RECT 611.470 294.835 611.640 295.005 ;
        RECT 613.050 294.835 613.220 295.005 ;
        RECT 614.630 294.835 614.800 295.005 ;
        RECT 615.900 294.815 616.070 294.985 ;
        RECT 617.480 294.815 617.650 294.985 ;
        RECT 619.060 294.815 619.230 294.985 ;
        RECT 620.280 294.825 620.450 294.995 ;
        RECT 621.860 294.825 622.030 294.995 ;
        RECT 623.440 294.825 623.610 294.995 ;
        RECT 624.600 294.815 624.770 294.985 ;
        RECT 626.180 294.815 626.350 294.985 ;
        RECT 627.760 294.815 627.930 294.985 ;
        RECT 628.980 295.045 629.150 295.215 ;
        RECT 601.250 294.455 601.420 294.625 ;
        RECT 601.250 294.095 601.420 294.265 ;
        RECT 601.250 293.735 601.420 293.905 ;
        RECT 628.980 294.685 629.150 294.855 ;
        RECT 840.940 295.815 841.110 295.985 ;
        RECT 841.300 295.815 841.470 295.985 ;
        RECT 841.660 295.815 841.830 295.985 ;
        RECT 842.020 295.815 842.190 295.985 ;
        RECT 845.245 294.645 845.415 294.815 ;
        RECT 845.725 294.645 845.895 294.815 ;
        RECT 846.205 294.645 846.375 294.815 ;
        RECT 846.685 294.645 846.855 294.815 ;
        RECT 847.165 294.645 847.335 294.815 ;
        RECT 847.645 294.645 847.815 294.815 ;
        RECT 848.125 294.645 848.295 294.815 ;
        RECT 628.980 294.325 629.150 294.495 ;
        RECT 628.980 293.965 629.150 294.135 ;
        RECT 861.335 294.375 861.505 294.545 ;
        RECT 861.815 294.375 861.985 294.545 ;
        RECT 862.295 294.375 862.465 294.545 ;
        RECT 862.775 294.375 862.945 294.545 ;
        RECT 863.255 294.375 863.425 294.545 ;
        RECT 863.735 294.375 863.905 294.545 ;
        RECT 864.215 294.375 864.385 294.545 ;
        RECT 845.920 294.165 846.090 294.335 ;
        RECT 846.280 294.165 846.450 294.335 ;
        RECT 846.640 294.165 846.810 294.335 ;
        RECT 847.000 294.165 847.170 294.335 ;
        RECT 847.360 294.165 847.530 294.335 ;
        RECT 847.720 294.165 847.890 294.335 ;
        RECT 635.215 293.795 635.385 293.965 ;
        RECT 635.695 293.795 635.865 293.965 ;
        RECT 636.175 293.795 636.345 293.965 ;
        RECT 639.405 293.885 639.575 294.055 ;
        RECT 639.885 293.885 640.055 294.055 ;
        RECT 640.365 293.885 640.535 294.055 ;
        RECT 643.505 293.865 643.675 294.035 ;
        RECT 643.985 293.865 644.155 294.035 ;
        RECT 644.465 293.865 644.635 294.035 ;
        RECT 595.325 293.345 595.495 293.515 ;
        RECT 595.805 293.345 595.975 293.515 ;
        RECT 596.285 293.345 596.455 293.515 ;
        RECT 601.250 293.375 601.420 293.545 ;
        RECT 595.960 292.865 596.130 293.035 ;
        RECT 596.320 292.865 596.490 293.035 ;
        RECT 602.430 293.355 602.600 293.525 ;
        RECT 604.010 293.355 604.180 293.525 ;
        RECT 605.590 293.355 605.760 293.525 ;
        RECT 606.950 293.365 607.120 293.535 ;
        RECT 608.530 293.365 608.700 293.535 ;
        RECT 610.110 293.365 610.280 293.535 ;
        RECT 611.470 293.365 611.640 293.535 ;
        RECT 613.050 293.365 613.220 293.535 ;
        RECT 614.630 293.365 614.800 293.535 ;
        RECT 615.900 293.345 616.070 293.515 ;
        RECT 617.480 293.345 617.650 293.515 ;
        RECT 619.060 293.345 619.230 293.515 ;
        RECT 620.280 293.355 620.450 293.525 ;
        RECT 621.860 293.355 622.030 293.525 ;
        RECT 623.440 293.355 623.610 293.525 ;
        RECT 624.600 293.345 624.770 293.515 ;
        RECT 626.180 293.345 626.350 293.515 ;
        RECT 627.760 293.345 627.930 293.515 ;
        RECT 628.980 293.605 629.150 293.775 ;
        RECT 628.980 293.245 629.150 293.415 ;
        RECT 635.180 293.315 635.350 293.485 ;
        RECT 635.540 293.315 635.710 293.485 ;
        RECT 639.370 293.405 639.540 293.575 ;
        RECT 639.730 293.405 639.900 293.575 ;
        RECT 643.470 293.385 643.640 293.555 ;
        RECT 643.830 293.385 644.000 293.555 ;
        RECT 819.095 293.285 819.265 293.455 ;
        RECT 819.575 293.285 819.745 293.455 ;
        RECT 820.055 293.285 820.225 293.455 ;
        RECT 820.535 293.285 820.705 293.455 ;
        RECT 821.015 293.285 821.185 293.455 ;
        RECT 821.495 293.285 821.665 293.455 ;
        RECT 821.975 293.285 822.145 293.455 ;
        RECT 819.050 292.805 819.220 292.975 ;
        RECT 819.410 292.805 819.580 292.975 ;
        RECT 819.770 292.805 819.940 292.975 ;
        RECT 820.490 292.805 820.660 292.975 ;
        RECT 820.850 292.805 821.020 292.975 ;
        RECT 821.210 292.805 821.380 292.975 ;
        RECT 821.570 292.805 821.740 292.975 ;
        RECT 862.010 293.895 862.180 294.065 ;
        RECT 862.370 293.895 862.540 294.065 ;
        RECT 862.730 293.895 862.900 294.065 ;
        RECT 863.090 293.895 863.260 294.065 ;
        RECT 863.450 293.895 863.620 294.065 ;
        RECT 863.810 293.895 863.980 294.065 ;
        RECT 855.995 292.745 856.165 292.915 ;
        RECT 856.475 292.745 856.645 292.915 ;
        RECT 856.955 292.745 857.125 292.915 ;
        RECT 857.435 292.745 857.605 292.915 ;
        RECT 857.915 292.745 858.085 292.915 ;
        RECT 858.395 292.745 858.565 292.915 ;
        RECT 858.875 292.745 859.045 292.915 ;
        RECT 855.950 292.265 856.120 292.435 ;
        RECT 856.310 292.265 856.480 292.435 ;
        RECT 856.670 292.265 856.840 292.435 ;
        RECT 824.545 291.115 824.715 291.285 ;
        RECT 825.025 291.115 825.195 291.285 ;
        RECT 825.505 291.115 825.675 291.285 ;
        RECT 825.985 291.115 826.155 291.285 ;
        RECT 826.465 291.115 826.635 291.285 ;
        RECT 826.945 291.115 827.115 291.285 ;
        RECT 827.425 291.115 827.595 291.285 ;
        RECT 389.010 289.765 389.180 289.935 ;
        RECT 382.430 289.405 382.600 289.575 ;
        RECT 382.430 286.295 382.600 286.465 ;
        RECT 382.430 285.935 382.600 286.105 ;
        RECT 382.430 282.825 382.600 282.995 ;
        RECT 382.430 282.465 382.600 282.635 ;
        RECT 382.430 279.355 382.600 279.525 ;
        RECT 382.430 278.995 382.600 279.165 ;
        RECT 375.850 275.885 376.020 276.055 ;
        RECT 369.690 275.625 369.860 275.795 ;
        RECT 382.430 275.885 382.600 276.055 ;
        RECT 389.010 289.405 389.180 289.575 ;
        RECT 389.010 286.295 389.180 286.465 ;
        RECT 389.010 285.935 389.180 286.105 ;
        RECT 389.010 282.825 389.180 282.995 ;
        RECT 389.010 282.465 389.180 282.635 ;
        RECT 389.010 279.355 389.180 279.525 ;
        RECT 389.010 278.995 389.180 279.165 ;
        RECT 389.010 275.885 389.180 276.055 ;
        RECT 375.850 275.525 376.020 275.695 ;
        RECT 382.430 275.525 382.600 275.695 ;
        RECT 394.005 289.235 394.175 289.405 ;
        RECT 394.005 288.875 394.175 289.045 ;
        RECT 394.005 288.515 394.175 288.685 ;
        RECT 394.005 288.155 394.175 288.325 ;
        RECT 394.005 287.795 394.175 287.965 ;
        RECT 394.005 287.435 394.175 287.605 ;
        RECT 394.005 287.075 394.175 287.245 ;
        RECT 394.005 286.715 394.175 286.885 ;
        RECT 394.005 286.355 394.175 286.525 ;
        RECT 394.005 285.995 394.175 286.165 ;
        RECT 394.005 285.635 394.175 285.805 ;
        RECT 394.005 285.275 394.175 285.445 ;
        RECT 394.005 284.915 394.175 285.085 ;
        RECT 394.005 284.555 394.175 284.725 ;
        RECT 394.005 284.195 394.175 284.365 ;
        RECT 394.005 283.835 394.175 284.005 ;
        RECT 394.005 283.475 394.175 283.645 ;
        RECT 394.005 283.115 394.175 283.285 ;
        RECT 394.005 282.755 394.175 282.925 ;
        RECT 394.005 282.395 394.175 282.565 ;
        RECT 394.005 282.035 394.175 282.205 ;
        RECT 394.005 281.675 394.175 281.845 ;
        RECT 394.005 281.315 394.175 281.485 ;
        RECT 394.005 280.955 394.175 281.125 ;
        RECT 394.005 280.595 394.175 280.765 ;
        RECT 394.005 280.235 394.175 280.405 ;
        RECT 394.005 279.875 394.175 280.045 ;
        RECT 394.005 279.515 394.175 279.685 ;
        RECT 394.005 279.155 394.175 279.325 ;
        RECT 394.005 278.795 394.175 278.965 ;
        RECT 394.005 278.435 394.175 278.605 ;
        RECT 394.005 278.075 394.175 278.245 ;
        RECT 394.005 277.715 394.175 277.885 ;
        RECT 394.005 277.355 394.175 277.525 ;
        RECT 394.005 276.995 394.175 277.165 ;
        RECT 394.005 276.635 394.175 276.805 ;
        RECT 395.100 289.835 395.270 290.005 ;
        RECT 395.100 289.475 395.270 289.645 ;
        RECT 395.100 286.365 395.270 286.535 ;
        RECT 395.100 286.005 395.270 286.175 ;
        RECT 395.100 282.895 395.270 283.065 ;
        RECT 395.100 282.535 395.270 282.705 ;
        RECT 395.100 279.425 395.270 279.595 ;
        RECT 395.100 279.065 395.270 279.235 ;
        RECT 398.390 289.835 398.560 290.005 ;
        RECT 398.390 289.475 398.560 289.645 ;
        RECT 398.390 286.365 398.560 286.535 ;
        RECT 398.390 286.005 398.560 286.175 ;
        RECT 398.390 282.895 398.560 283.065 ;
        RECT 398.390 282.535 398.560 282.705 ;
        RECT 398.390 279.425 398.560 279.595 ;
        RECT 398.390 279.065 398.560 279.235 ;
        RECT 395.100 275.955 395.270 276.125 ;
        RECT 389.010 275.525 389.180 275.695 ;
        RECT 395.100 275.595 395.270 275.765 ;
        RECT 398.390 275.955 398.560 276.125 ;
        RECT 401.680 289.835 401.850 290.005 ;
        RECT 401.680 289.475 401.850 289.645 ;
        RECT 401.680 286.365 401.850 286.535 ;
        RECT 401.680 286.005 401.850 286.175 ;
        RECT 401.680 282.895 401.850 283.065 ;
        RECT 401.680 282.535 401.850 282.705 ;
        RECT 401.680 279.425 401.850 279.595 ;
        RECT 401.680 279.065 401.850 279.235 ;
        RECT 401.680 275.955 401.850 276.125 ;
        RECT 404.970 289.835 405.140 290.005 ;
        RECT 408.260 289.835 408.430 290.005 ;
        RECT 824.500 290.635 824.670 290.805 ;
        RECT 824.860 290.635 825.030 290.805 ;
        RECT 825.220 290.635 825.390 290.805 ;
        RECT 404.970 289.475 405.140 289.645 ;
        RECT 404.970 286.365 405.140 286.535 ;
        RECT 404.970 286.005 405.140 286.175 ;
        RECT 404.970 282.895 405.140 283.065 ;
        RECT 404.970 282.535 405.140 282.705 ;
        RECT 404.970 279.425 405.140 279.595 ;
        RECT 404.970 279.065 405.140 279.235 ;
        RECT 404.970 275.955 405.140 276.125 ;
        RECT 408.260 289.475 408.430 289.645 ;
        RECT 825.940 290.635 826.110 290.805 ;
        RECT 826.300 290.635 826.470 290.805 ;
        RECT 826.660 290.635 826.830 290.805 ;
        RECT 827.020 290.635 827.190 290.805 ;
        RECT 830.085 291.135 830.255 291.305 ;
        RECT 830.565 291.135 830.735 291.305 ;
        RECT 831.045 291.135 831.215 291.305 ;
        RECT 831.525 291.135 831.695 291.305 ;
        RECT 832.005 291.135 832.175 291.305 ;
        RECT 832.485 291.135 832.655 291.305 ;
        RECT 832.965 291.135 833.135 291.305 ;
        RECT 833.445 291.135 833.615 291.305 ;
        RECT 833.925 291.135 834.095 291.305 ;
        RECT 834.405 291.135 834.575 291.305 ;
        RECT 834.885 291.135 835.055 291.305 ;
        RECT 839.555 291.175 839.725 291.345 ;
        RECT 840.035 291.175 840.205 291.345 ;
        RECT 840.515 291.175 840.685 291.345 ;
        RECT 840.995 291.175 841.165 291.345 ;
        RECT 841.475 291.175 841.645 291.345 ;
        RECT 841.955 291.175 842.125 291.345 ;
        RECT 842.435 291.175 842.605 291.345 ;
        RECT 857.390 292.265 857.560 292.435 ;
        RECT 857.750 292.265 857.920 292.435 ;
        RECT 858.110 292.265 858.280 292.435 ;
        RECT 858.470 292.265 858.640 292.435 ;
        RECT 830.490 290.655 830.660 290.825 ;
        RECT 830.850 290.655 831.020 290.825 ;
        RECT 831.210 290.655 831.380 290.825 ;
        RECT 831.570 290.655 831.740 290.825 ;
        RECT 831.930 290.655 832.100 290.825 ;
        RECT 832.290 290.655 832.460 290.825 ;
        RECT 833.015 290.655 833.185 290.825 ;
        RECT 833.375 290.655 833.545 290.825 ;
        RECT 833.735 290.655 833.905 290.825 ;
        RECT 834.095 290.655 834.265 290.825 ;
        RECT 834.455 290.655 834.625 290.825 ;
        RECT 839.510 290.695 839.680 290.865 ;
        RECT 839.870 290.695 840.040 290.865 ;
        RECT 840.230 290.695 840.400 290.865 ;
        RECT 840.950 290.695 841.120 290.865 ;
        RECT 841.310 290.695 841.480 290.865 ;
        RECT 841.670 290.695 841.840 290.865 ;
        RECT 842.030 290.695 842.200 290.865 ;
        RECT 819.065 288.125 819.235 288.295 ;
        RECT 819.545 288.125 819.715 288.295 ;
        RECT 820.025 288.125 820.195 288.295 ;
        RECT 820.505 288.125 820.675 288.295 ;
        RECT 820.985 288.125 821.155 288.295 ;
        RECT 821.465 288.125 821.635 288.295 ;
        RECT 821.945 288.125 822.115 288.295 ;
        RECT 408.260 286.365 408.430 286.535 ;
        RECT 819.020 287.645 819.190 287.815 ;
        RECT 819.380 287.645 819.550 287.815 ;
        RECT 819.740 287.645 819.910 287.815 ;
        RECT 820.460 287.645 820.630 287.815 ;
        RECT 820.820 287.645 820.990 287.815 ;
        RECT 821.180 287.645 821.350 287.815 ;
        RECT 821.540 287.645 821.710 287.815 ;
        RECT 856.065 287.345 856.235 287.515 ;
        RECT 856.545 287.345 856.715 287.515 ;
        RECT 857.025 287.345 857.195 287.515 ;
        RECT 857.505 287.345 857.675 287.515 ;
        RECT 857.985 287.345 858.155 287.515 ;
        RECT 858.465 287.345 858.635 287.515 ;
        RECT 858.945 287.345 859.115 287.515 ;
        RECT 856.020 286.865 856.190 287.035 ;
        RECT 856.380 286.865 856.550 287.035 ;
        RECT 856.740 286.865 856.910 287.035 ;
        RECT 408.260 286.005 408.430 286.175 ;
        RECT 857.460 286.865 857.630 287.035 ;
        RECT 857.820 286.865 857.990 287.035 ;
        RECT 858.180 286.865 858.350 287.035 ;
        RECT 858.540 286.865 858.710 287.035 ;
        RECT 861.415 285.325 861.585 285.495 ;
        RECT 861.895 285.325 862.065 285.495 ;
        RECT 862.375 285.325 862.545 285.495 ;
        RECT 862.855 285.325 863.025 285.495 ;
        RECT 863.335 285.325 863.505 285.495 ;
        RECT 863.815 285.325 863.985 285.495 ;
        RECT 864.295 285.325 864.465 285.495 ;
        RECT 862.090 284.845 862.260 285.015 ;
        RECT 862.450 284.845 862.620 285.015 ;
        RECT 862.810 284.845 862.980 285.015 ;
        RECT 863.170 284.845 863.340 285.015 ;
        RECT 863.530 284.845 863.700 285.015 ;
        RECT 863.890 284.845 864.060 285.015 ;
        RECT 799.685 283.435 799.855 283.605 ;
        RECT 800.165 283.435 800.335 283.605 ;
        RECT 800.645 283.435 800.815 283.605 ;
        RECT 408.260 282.895 408.430 283.065 ;
        RECT 408.260 282.535 408.430 282.705 ;
        RECT 799.650 282.955 799.820 283.125 ;
        RECT 800.010 282.955 800.180 283.125 ;
        RECT 819.505 283.095 819.675 283.265 ;
        RECT 819.985 283.095 820.155 283.265 ;
        RECT 820.465 283.095 820.635 283.265 ;
        RECT 820.945 283.095 821.115 283.265 ;
        RECT 821.425 283.095 821.595 283.265 ;
        RECT 821.905 283.095 822.075 283.265 ;
        RECT 822.385 283.095 822.555 283.265 ;
        RECT 822.865 283.095 823.035 283.265 ;
        RECT 823.345 283.095 823.515 283.265 ;
        RECT 823.825 283.095 823.995 283.265 ;
        RECT 824.305 283.095 824.475 283.265 ;
        RECT 828.115 283.005 828.285 283.175 ;
        RECT 828.595 283.005 828.765 283.175 ;
        RECT 829.075 283.005 829.245 283.175 ;
        RECT 829.555 283.005 829.725 283.175 ;
        RECT 830.035 283.005 830.205 283.175 ;
        RECT 830.515 283.005 830.685 283.175 ;
        RECT 830.995 283.005 831.165 283.175 ;
        RECT 679.545 282.215 679.715 282.385 ;
        RECT 680.025 282.215 680.195 282.385 ;
        RECT 680.505 282.215 680.675 282.385 ;
        RECT 680.985 282.215 681.155 282.385 ;
        RECT 681.465 282.215 681.635 282.385 ;
        RECT 681.945 282.215 682.115 282.385 ;
        RECT 682.425 282.215 682.595 282.385 ;
        RECT 682.905 282.215 683.075 282.385 ;
        RECT 683.385 282.215 683.555 282.385 ;
        RECT 683.865 282.215 684.035 282.385 ;
        RECT 684.345 282.215 684.515 282.385 ;
        RECT 679.950 281.735 680.120 281.905 ;
        RECT 680.310 281.735 680.480 281.905 ;
        RECT 680.670 281.735 680.840 281.905 ;
        RECT 681.030 281.735 681.200 281.905 ;
        RECT 681.390 281.735 681.560 281.905 ;
        RECT 681.750 281.735 681.920 281.905 ;
        RECT 682.475 281.735 682.645 281.905 ;
        RECT 682.835 281.735 683.005 281.905 ;
        RECT 683.195 281.735 683.365 281.905 ;
        RECT 683.555 281.735 683.725 281.905 ;
        RECT 683.915 281.735 684.085 281.905 ;
        RECT 696.825 282.225 696.995 282.395 ;
        RECT 697.305 282.225 697.475 282.395 ;
        RECT 697.785 282.225 697.955 282.395 ;
        RECT 698.265 282.225 698.435 282.395 ;
        RECT 698.745 282.225 698.915 282.395 ;
        RECT 699.225 282.225 699.395 282.395 ;
        RECT 699.705 282.225 699.875 282.395 ;
        RECT 700.185 282.225 700.355 282.395 ;
        RECT 700.665 282.225 700.835 282.395 ;
        RECT 701.145 282.225 701.315 282.395 ;
        RECT 701.625 282.225 701.795 282.395 ;
        RECT 697.230 281.745 697.400 281.915 ;
        RECT 697.590 281.745 697.760 281.915 ;
        RECT 697.950 281.745 698.120 281.915 ;
        RECT 698.310 281.745 698.480 281.915 ;
        RECT 698.670 281.745 698.840 281.915 ;
        RECT 699.030 281.745 699.200 281.915 ;
        RECT 699.755 281.745 699.925 281.915 ;
        RECT 700.115 281.745 700.285 281.915 ;
        RECT 700.475 281.745 700.645 281.915 ;
        RECT 700.835 281.745 701.005 281.915 ;
        RECT 701.195 281.745 701.365 281.915 ;
        RECT 714.595 282.225 714.765 282.395 ;
        RECT 715.075 282.225 715.245 282.395 ;
        RECT 715.555 282.225 715.725 282.395 ;
        RECT 716.035 282.225 716.205 282.395 ;
        RECT 716.515 282.225 716.685 282.395 ;
        RECT 716.995 282.225 717.165 282.395 ;
        RECT 717.475 282.225 717.645 282.395 ;
        RECT 717.955 282.225 718.125 282.395 ;
        RECT 718.435 282.225 718.605 282.395 ;
        RECT 718.915 282.225 719.085 282.395 ;
        RECT 719.395 282.225 719.565 282.395 ;
        RECT 715.000 281.745 715.170 281.915 ;
        RECT 715.360 281.745 715.530 281.915 ;
        RECT 715.720 281.745 715.890 281.915 ;
        RECT 716.080 281.745 716.250 281.915 ;
        RECT 716.440 281.745 716.610 281.915 ;
        RECT 716.800 281.745 716.970 281.915 ;
        RECT 717.525 281.745 717.695 281.915 ;
        RECT 717.885 281.745 718.055 281.915 ;
        RECT 718.245 281.745 718.415 281.915 ;
        RECT 718.605 281.745 718.775 281.915 ;
        RECT 718.965 281.745 719.135 281.915 ;
        RECT 731.835 282.225 732.005 282.395 ;
        RECT 732.315 282.225 732.485 282.395 ;
        RECT 732.795 282.225 732.965 282.395 ;
        RECT 733.275 282.225 733.445 282.395 ;
        RECT 733.755 282.225 733.925 282.395 ;
        RECT 734.235 282.225 734.405 282.395 ;
        RECT 734.715 282.225 734.885 282.395 ;
        RECT 735.195 282.225 735.365 282.395 ;
        RECT 735.675 282.225 735.845 282.395 ;
        RECT 736.155 282.225 736.325 282.395 ;
        RECT 736.635 282.225 736.805 282.395 ;
        RECT 732.240 281.745 732.410 281.915 ;
        RECT 732.600 281.745 732.770 281.915 ;
        RECT 732.960 281.745 733.130 281.915 ;
        RECT 733.320 281.745 733.490 281.915 ;
        RECT 733.680 281.745 733.850 281.915 ;
        RECT 734.040 281.745 734.210 281.915 ;
        RECT 734.765 281.745 734.935 281.915 ;
        RECT 735.125 281.745 735.295 281.915 ;
        RECT 735.485 281.745 735.655 281.915 ;
        RECT 735.845 281.745 736.015 281.915 ;
        RECT 736.205 281.745 736.375 281.915 ;
        RECT 749.315 282.235 749.485 282.405 ;
        RECT 749.795 282.235 749.965 282.405 ;
        RECT 750.275 282.235 750.445 282.405 ;
        RECT 750.755 282.235 750.925 282.405 ;
        RECT 751.235 282.235 751.405 282.405 ;
        RECT 751.715 282.235 751.885 282.405 ;
        RECT 752.195 282.235 752.365 282.405 ;
        RECT 752.675 282.235 752.845 282.405 ;
        RECT 753.155 282.235 753.325 282.405 ;
        RECT 753.635 282.235 753.805 282.405 ;
        RECT 754.115 282.235 754.285 282.405 ;
        RECT 749.720 281.755 749.890 281.925 ;
        RECT 750.080 281.755 750.250 281.925 ;
        RECT 750.440 281.755 750.610 281.925 ;
        RECT 750.800 281.755 750.970 281.925 ;
        RECT 751.160 281.755 751.330 281.925 ;
        RECT 751.520 281.755 751.690 281.925 ;
        RECT 752.245 281.755 752.415 281.925 ;
        RECT 752.605 281.755 752.775 281.925 ;
        RECT 752.965 281.755 753.135 281.925 ;
        RECT 753.325 281.755 753.495 281.925 ;
        RECT 753.685 281.755 753.855 281.925 ;
        RECT 819.910 282.615 820.080 282.785 ;
        RECT 820.270 282.615 820.440 282.785 ;
        RECT 820.630 282.615 820.800 282.785 ;
        RECT 820.990 282.615 821.160 282.785 ;
        RECT 821.350 282.615 821.520 282.785 ;
        RECT 821.710 282.615 821.880 282.785 ;
        RECT 822.435 282.615 822.605 282.785 ;
        RECT 822.795 282.615 822.965 282.785 ;
        RECT 823.155 282.615 823.325 282.785 ;
        RECT 823.515 282.615 823.685 282.785 ;
        RECT 823.875 282.615 824.045 282.785 ;
        RECT 828.070 282.525 828.240 282.695 ;
        RECT 828.430 282.525 828.600 282.695 ;
        RECT 828.790 282.525 828.960 282.695 ;
        RECT 829.510 282.525 829.680 282.695 ;
        RECT 829.870 282.525 830.040 282.695 ;
        RECT 830.230 282.525 830.400 282.695 ;
        RECT 830.590 282.525 830.760 282.695 ;
        RECT 833.405 283.005 833.575 283.175 ;
        RECT 833.885 283.005 834.055 283.175 ;
        RECT 834.365 283.005 834.535 283.175 ;
        RECT 834.845 283.005 835.015 283.175 ;
        RECT 835.325 283.005 835.495 283.175 ;
        RECT 835.805 283.005 835.975 283.175 ;
        RECT 836.285 283.005 836.455 283.175 ;
        RECT 836.765 283.005 836.935 283.175 ;
        RECT 837.245 283.005 837.415 283.175 ;
        RECT 837.725 283.005 837.895 283.175 ;
        RECT 838.205 283.005 838.375 283.175 ;
        RECT 833.810 282.525 833.980 282.695 ;
        RECT 834.170 282.525 834.340 282.695 ;
        RECT 834.530 282.525 834.700 282.695 ;
        RECT 834.890 282.525 835.060 282.695 ;
        RECT 835.250 282.525 835.420 282.695 ;
        RECT 835.610 282.525 835.780 282.695 ;
        RECT 836.335 282.525 836.505 282.695 ;
        RECT 836.695 282.525 836.865 282.695 ;
        RECT 837.055 282.525 837.225 282.695 ;
        RECT 837.415 282.525 837.585 282.695 ;
        RECT 837.775 282.525 837.945 282.695 ;
        RECT 840.615 283.005 840.785 283.175 ;
        RECT 841.095 283.005 841.265 283.175 ;
        RECT 841.575 283.005 841.745 283.175 ;
        RECT 842.055 283.005 842.225 283.175 ;
        RECT 842.535 283.005 842.705 283.175 ;
        RECT 843.015 283.005 843.185 283.175 ;
        RECT 843.495 283.005 843.665 283.175 ;
        RECT 843.975 283.005 844.145 283.175 ;
        RECT 846.455 283.005 846.625 283.175 ;
        RECT 846.935 283.005 847.105 283.175 ;
        RECT 847.415 283.005 847.585 283.175 ;
        RECT 847.895 283.005 848.065 283.175 ;
        RECT 848.375 283.005 848.545 283.175 ;
        RECT 848.855 283.005 849.025 283.175 ;
        RECT 849.335 283.005 849.505 283.175 ;
        RECT 849.815 283.005 849.985 283.175 ;
        RECT 850.295 283.005 850.465 283.175 ;
        RECT 850.775 283.005 850.945 283.175 ;
        RECT 851.255 283.005 851.425 283.175 ;
        RECT 841.050 282.525 841.220 282.695 ;
        RECT 841.410 282.525 841.580 282.695 ;
        RECT 841.770 282.525 841.940 282.695 ;
        RECT 842.690 282.525 842.860 282.695 ;
        RECT 843.050 282.525 843.220 282.695 ;
        RECT 843.410 282.525 843.580 282.695 ;
        RECT 846.860 282.525 847.030 282.695 ;
        RECT 847.220 282.525 847.390 282.695 ;
        RECT 847.580 282.525 847.750 282.695 ;
        RECT 847.940 282.525 848.110 282.695 ;
        RECT 848.300 282.525 848.470 282.695 ;
        RECT 848.660 282.525 848.830 282.695 ;
        RECT 849.385 282.525 849.555 282.695 ;
        RECT 849.745 282.525 849.915 282.695 ;
        RECT 850.105 282.525 850.275 282.695 ;
        RECT 850.465 282.525 850.635 282.695 ;
        RECT 850.825 282.525 850.995 282.695 ;
        RECT 856.085 281.885 856.255 282.055 ;
        RECT 856.565 281.885 856.735 282.055 ;
        RECT 857.045 281.885 857.215 282.055 ;
        RECT 857.525 281.885 857.695 282.055 ;
        RECT 858.005 281.885 858.175 282.055 ;
        RECT 858.485 281.885 858.655 282.055 ;
        RECT 858.965 281.885 859.135 282.055 ;
        RECT 856.040 281.405 856.210 281.575 ;
        RECT 856.400 281.405 856.570 281.575 ;
        RECT 856.760 281.405 856.930 281.575 ;
        RECT 682.330 280.125 682.500 280.295 ;
        RECT 699.630 280.175 699.800 280.345 ;
        RECT 717.420 280.215 717.590 280.385 ;
        RECT 734.680 280.245 734.850 280.415 ;
        RECT 752.150 280.235 752.320 280.405 ;
        RECT 857.480 281.405 857.650 281.575 ;
        RECT 857.840 281.405 858.010 281.575 ;
        RECT 858.200 281.405 858.370 281.575 ;
        RECT 858.560 281.405 858.730 281.575 ;
        RECT 408.260 279.425 408.430 279.595 ;
        RECT 408.260 279.065 408.430 279.235 ;
        RECT 398.390 275.595 398.560 275.765 ;
        RECT 401.680 275.595 401.850 275.765 ;
        RECT 404.970 275.595 405.140 275.765 ;
        RECT 408.260 275.955 408.430 276.125 ;
        RECT 408.260 275.595 408.430 275.765 ;
        RECT 601.170 276.345 601.340 276.515 ;
        RECT 602.350 276.355 602.520 276.525 ;
        RECT 603.930 276.355 604.100 276.525 ;
        RECT 605.510 276.355 605.680 276.525 ;
        RECT 606.870 276.365 607.040 276.535 ;
        RECT 608.450 276.365 608.620 276.535 ;
        RECT 610.030 276.365 610.200 276.535 ;
        RECT 611.390 276.365 611.560 276.535 ;
        RECT 612.970 276.365 613.140 276.535 ;
        RECT 614.550 276.365 614.720 276.535 ;
        RECT 615.820 276.345 615.990 276.515 ;
        RECT 617.400 276.345 617.570 276.515 ;
        RECT 618.980 276.345 619.150 276.515 ;
        RECT 620.200 276.355 620.370 276.525 ;
        RECT 621.780 276.355 621.950 276.525 ;
        RECT 623.360 276.355 623.530 276.525 ;
        RECT 624.520 276.345 624.690 276.515 ;
        RECT 626.100 276.345 626.270 276.515 ;
        RECT 627.680 276.345 627.850 276.515 ;
        RECT 628.900 276.575 629.070 276.745 ;
        RECT 679.955 276.555 680.125 276.725 ;
        RECT 680.435 276.555 680.605 276.725 ;
        RECT 680.915 276.555 681.085 276.725 ;
        RECT 681.395 276.555 681.565 276.725 ;
        RECT 681.875 276.555 682.045 276.725 ;
        RECT 682.355 276.555 682.525 276.725 ;
        RECT 682.835 276.555 683.005 276.725 ;
        RECT 683.315 276.555 683.485 276.725 ;
        RECT 683.795 276.555 683.965 276.725 ;
        RECT 684.275 276.555 684.445 276.725 ;
        RECT 684.755 276.555 684.925 276.725 ;
        RECT 601.170 275.985 601.340 276.155 ;
        RECT 601.170 275.625 601.340 275.795 ;
        RECT 601.170 275.265 601.340 275.435 ;
        RECT 628.900 276.215 629.070 276.385 ;
        RECT 628.900 275.855 629.070 276.025 ;
        RECT 628.900 275.495 629.070 275.665 ;
        RECT 680.360 276.075 680.530 276.245 ;
        RECT 680.720 276.075 680.890 276.245 ;
        RECT 681.080 276.075 681.250 276.245 ;
        RECT 681.440 276.075 681.610 276.245 ;
        RECT 681.800 276.075 681.970 276.245 ;
        RECT 682.160 276.075 682.330 276.245 ;
        RECT 635.135 275.325 635.305 275.495 ;
        RECT 635.615 275.325 635.785 275.495 ;
        RECT 636.095 275.325 636.265 275.495 ;
        RECT 639.325 275.415 639.495 275.585 ;
        RECT 639.805 275.415 639.975 275.585 ;
        RECT 640.285 275.415 640.455 275.585 ;
        RECT 643.425 275.395 643.595 275.565 ;
        RECT 643.905 275.395 644.075 275.565 ;
        RECT 644.385 275.395 644.555 275.565 ;
        RECT 682.885 276.075 683.055 276.245 ;
        RECT 683.245 276.075 683.415 276.245 ;
        RECT 683.605 276.075 683.775 276.245 ;
        RECT 683.965 276.075 684.135 276.245 ;
        RECT 684.325 276.075 684.495 276.245 ;
        RECT 687.195 276.515 687.365 276.685 ;
        RECT 687.675 276.515 687.845 276.685 ;
        RECT 688.155 276.515 688.325 276.685 ;
        RECT 688.635 276.515 688.805 276.685 ;
        RECT 689.115 276.515 689.285 276.685 ;
        RECT 689.595 276.515 689.765 276.685 ;
        RECT 690.075 276.515 690.245 276.685 ;
        RECT 690.555 276.515 690.725 276.685 ;
        RECT 691.035 276.515 691.205 276.685 ;
        RECT 691.515 276.515 691.685 276.685 ;
        RECT 691.995 276.515 692.165 276.685 ;
        RECT 697.185 276.575 697.355 276.745 ;
        RECT 697.665 276.575 697.835 276.745 ;
        RECT 698.145 276.575 698.315 276.745 ;
        RECT 698.625 276.575 698.795 276.745 ;
        RECT 699.105 276.575 699.275 276.745 ;
        RECT 699.585 276.575 699.755 276.745 ;
        RECT 700.065 276.575 700.235 276.745 ;
        RECT 700.545 276.575 700.715 276.745 ;
        RECT 701.025 276.575 701.195 276.745 ;
        RECT 701.505 276.575 701.675 276.745 ;
        RECT 701.985 276.575 702.155 276.745 ;
        RECT 687.600 276.035 687.770 276.205 ;
        RECT 687.960 276.035 688.130 276.205 ;
        RECT 688.320 276.035 688.490 276.205 ;
        RECT 688.680 276.035 688.850 276.205 ;
        RECT 689.040 276.035 689.210 276.205 ;
        RECT 689.400 276.035 689.570 276.205 ;
        RECT 690.125 276.035 690.295 276.205 ;
        RECT 690.485 276.035 690.655 276.205 ;
        RECT 690.845 276.035 691.015 276.205 ;
        RECT 691.205 276.035 691.375 276.205 ;
        RECT 691.565 276.035 691.735 276.205 ;
        RECT 697.590 276.095 697.760 276.265 ;
        RECT 697.950 276.095 698.120 276.265 ;
        RECT 698.310 276.095 698.480 276.265 ;
        RECT 698.670 276.095 698.840 276.265 ;
        RECT 699.030 276.095 699.200 276.265 ;
        RECT 699.390 276.095 699.560 276.265 ;
        RECT 700.115 276.095 700.285 276.265 ;
        RECT 700.475 276.095 700.645 276.265 ;
        RECT 700.835 276.095 701.005 276.265 ;
        RECT 701.195 276.095 701.365 276.265 ;
        RECT 701.555 276.095 701.725 276.265 ;
        RECT 704.425 276.535 704.595 276.705 ;
        RECT 704.905 276.535 705.075 276.705 ;
        RECT 705.385 276.535 705.555 276.705 ;
        RECT 705.865 276.535 706.035 276.705 ;
        RECT 706.345 276.535 706.515 276.705 ;
        RECT 706.825 276.535 706.995 276.705 ;
        RECT 707.305 276.535 707.475 276.705 ;
        RECT 707.785 276.535 707.955 276.705 ;
        RECT 708.265 276.535 708.435 276.705 ;
        RECT 708.745 276.535 708.915 276.705 ;
        RECT 709.225 276.535 709.395 276.705 ;
        RECT 714.755 276.675 714.925 276.845 ;
        RECT 715.235 276.675 715.405 276.845 ;
        RECT 715.715 276.675 715.885 276.845 ;
        RECT 716.195 276.675 716.365 276.845 ;
        RECT 716.675 276.675 716.845 276.845 ;
        RECT 717.155 276.675 717.325 276.845 ;
        RECT 717.635 276.675 717.805 276.845 ;
        RECT 718.115 276.675 718.285 276.845 ;
        RECT 718.595 276.675 718.765 276.845 ;
        RECT 719.075 276.675 719.245 276.845 ;
        RECT 719.555 276.675 719.725 276.845 ;
        RECT 704.830 276.055 705.000 276.225 ;
        RECT 705.190 276.055 705.360 276.225 ;
        RECT 705.550 276.055 705.720 276.225 ;
        RECT 705.910 276.055 706.080 276.225 ;
        RECT 706.270 276.055 706.440 276.225 ;
        RECT 706.630 276.055 706.800 276.225 ;
        RECT 707.355 276.055 707.525 276.225 ;
        RECT 707.715 276.055 707.885 276.225 ;
        RECT 708.075 276.055 708.245 276.225 ;
        RECT 708.435 276.055 708.605 276.225 ;
        RECT 708.795 276.055 708.965 276.225 ;
        RECT 715.160 276.195 715.330 276.365 ;
        RECT 715.520 276.195 715.690 276.365 ;
        RECT 715.880 276.195 716.050 276.365 ;
        RECT 716.240 276.195 716.410 276.365 ;
        RECT 716.600 276.195 716.770 276.365 ;
        RECT 716.960 276.195 717.130 276.365 ;
        RECT 717.685 276.195 717.855 276.365 ;
        RECT 718.045 276.195 718.215 276.365 ;
        RECT 718.405 276.195 718.575 276.365 ;
        RECT 718.765 276.195 718.935 276.365 ;
        RECT 719.125 276.195 719.295 276.365 ;
        RECT 721.995 276.635 722.165 276.805 ;
        RECT 722.475 276.635 722.645 276.805 ;
        RECT 722.955 276.635 723.125 276.805 ;
        RECT 723.435 276.635 723.605 276.805 ;
        RECT 723.915 276.635 724.085 276.805 ;
        RECT 724.395 276.635 724.565 276.805 ;
        RECT 724.875 276.635 725.045 276.805 ;
        RECT 725.355 276.635 725.525 276.805 ;
        RECT 725.835 276.635 726.005 276.805 ;
        RECT 726.315 276.635 726.485 276.805 ;
        RECT 726.795 276.635 726.965 276.805 ;
        RECT 731.925 276.705 732.095 276.875 ;
        RECT 732.405 276.705 732.575 276.875 ;
        RECT 732.885 276.705 733.055 276.875 ;
        RECT 733.365 276.705 733.535 276.875 ;
        RECT 733.845 276.705 734.015 276.875 ;
        RECT 734.325 276.705 734.495 276.875 ;
        RECT 734.805 276.705 734.975 276.875 ;
        RECT 735.285 276.705 735.455 276.875 ;
        RECT 735.765 276.705 735.935 276.875 ;
        RECT 736.245 276.705 736.415 276.875 ;
        RECT 736.725 276.705 736.895 276.875 ;
        RECT 722.400 276.155 722.570 276.325 ;
        RECT 722.760 276.155 722.930 276.325 ;
        RECT 723.120 276.155 723.290 276.325 ;
        RECT 723.480 276.155 723.650 276.325 ;
        RECT 723.840 276.155 724.010 276.325 ;
        RECT 724.200 276.155 724.370 276.325 ;
        RECT 724.925 276.155 725.095 276.325 ;
        RECT 725.285 276.155 725.455 276.325 ;
        RECT 725.645 276.155 725.815 276.325 ;
        RECT 726.005 276.155 726.175 276.325 ;
        RECT 726.365 276.155 726.535 276.325 ;
        RECT 732.330 276.225 732.500 276.395 ;
        RECT 732.690 276.225 732.860 276.395 ;
        RECT 733.050 276.225 733.220 276.395 ;
        RECT 733.410 276.225 733.580 276.395 ;
        RECT 733.770 276.225 733.940 276.395 ;
        RECT 734.130 276.225 734.300 276.395 ;
        RECT 734.855 276.225 735.025 276.395 ;
        RECT 735.215 276.225 735.385 276.395 ;
        RECT 735.575 276.225 735.745 276.395 ;
        RECT 735.935 276.225 736.105 276.395 ;
        RECT 736.295 276.225 736.465 276.395 ;
        RECT 739.165 276.665 739.335 276.835 ;
        RECT 739.645 276.665 739.815 276.835 ;
        RECT 740.125 276.665 740.295 276.835 ;
        RECT 740.605 276.665 740.775 276.835 ;
        RECT 741.085 276.665 741.255 276.835 ;
        RECT 741.565 276.665 741.735 276.835 ;
        RECT 742.045 276.665 742.215 276.835 ;
        RECT 742.525 276.665 742.695 276.835 ;
        RECT 743.005 276.665 743.175 276.835 ;
        RECT 743.485 276.665 743.655 276.835 ;
        RECT 743.965 276.665 744.135 276.835 ;
        RECT 749.735 276.765 749.905 276.935 ;
        RECT 750.215 276.765 750.385 276.935 ;
        RECT 750.695 276.765 750.865 276.935 ;
        RECT 751.175 276.765 751.345 276.935 ;
        RECT 751.655 276.765 751.825 276.935 ;
        RECT 752.135 276.765 752.305 276.935 ;
        RECT 752.615 276.765 752.785 276.935 ;
        RECT 753.095 276.765 753.265 276.935 ;
        RECT 753.575 276.765 753.745 276.935 ;
        RECT 754.055 276.765 754.225 276.935 ;
        RECT 754.535 276.765 754.705 276.935 ;
        RECT 739.570 276.185 739.740 276.355 ;
        RECT 739.930 276.185 740.100 276.355 ;
        RECT 740.290 276.185 740.460 276.355 ;
        RECT 740.650 276.185 740.820 276.355 ;
        RECT 741.010 276.185 741.180 276.355 ;
        RECT 741.370 276.185 741.540 276.355 ;
        RECT 742.095 276.185 742.265 276.355 ;
        RECT 742.455 276.185 742.625 276.355 ;
        RECT 742.815 276.185 742.985 276.355 ;
        RECT 743.175 276.185 743.345 276.355 ;
        RECT 743.535 276.185 743.705 276.355 ;
        RECT 750.140 276.285 750.310 276.455 ;
        RECT 750.500 276.285 750.670 276.455 ;
        RECT 750.860 276.285 751.030 276.455 ;
        RECT 751.220 276.285 751.390 276.455 ;
        RECT 751.580 276.285 751.750 276.455 ;
        RECT 751.940 276.285 752.110 276.455 ;
        RECT 752.665 276.285 752.835 276.455 ;
        RECT 753.025 276.285 753.195 276.455 ;
        RECT 753.385 276.285 753.555 276.455 ;
        RECT 753.745 276.285 753.915 276.455 ;
        RECT 754.105 276.285 754.275 276.455 ;
        RECT 756.975 276.725 757.145 276.895 ;
        RECT 757.455 276.725 757.625 276.895 ;
        RECT 757.935 276.725 758.105 276.895 ;
        RECT 758.415 276.725 758.585 276.895 ;
        RECT 758.895 276.725 759.065 276.895 ;
        RECT 759.375 276.725 759.545 276.895 ;
        RECT 759.855 276.725 760.025 276.895 ;
        RECT 760.335 276.725 760.505 276.895 ;
        RECT 760.815 276.725 760.985 276.895 ;
        RECT 761.295 276.725 761.465 276.895 ;
        RECT 761.775 276.725 761.945 276.895 ;
        RECT 757.380 276.245 757.550 276.415 ;
        RECT 757.740 276.245 757.910 276.415 ;
        RECT 758.100 276.245 758.270 276.415 ;
        RECT 758.460 276.245 758.630 276.415 ;
        RECT 758.820 276.245 758.990 276.415 ;
        RECT 759.180 276.245 759.350 276.415 ;
        RECT 759.905 276.245 760.075 276.415 ;
        RECT 760.265 276.245 760.435 276.415 ;
        RECT 760.625 276.245 760.795 276.415 ;
        RECT 760.985 276.245 761.155 276.415 ;
        RECT 761.345 276.245 761.515 276.415 ;
        RECT 781.115 275.395 781.285 275.565 ;
        RECT 781.595 275.395 781.765 275.565 ;
        RECT 782.075 275.395 782.245 275.565 ;
        RECT 782.555 275.395 782.725 275.565 ;
        RECT 783.035 275.395 783.205 275.565 ;
        RECT 783.515 275.395 783.685 275.565 ;
        RECT 783.995 275.395 784.165 275.565 ;
        RECT 784.475 275.395 784.645 275.565 ;
        RECT 784.955 275.395 785.125 275.565 ;
        RECT 785.435 275.395 785.605 275.565 ;
        RECT 785.915 275.395 786.085 275.565 ;
        RECT 786.395 275.395 786.565 275.565 ;
        RECT 786.875 275.395 787.045 275.565 ;
        RECT 787.355 275.395 787.525 275.565 ;
        RECT 787.835 275.395 788.005 275.565 ;
        RECT 788.315 275.395 788.485 275.565 ;
        RECT 788.795 275.395 788.965 275.565 ;
        RECT 789.275 275.395 789.445 275.565 ;
        RECT 789.755 275.395 789.925 275.565 ;
        RECT 790.235 275.395 790.405 275.565 ;
        RECT 790.715 275.395 790.885 275.565 ;
        RECT 791.195 275.395 791.365 275.565 ;
        RECT 791.675 275.395 791.845 275.565 ;
        RECT 792.155 275.395 792.325 275.565 ;
        RECT 792.635 275.395 792.805 275.565 ;
        RECT 793.115 275.395 793.285 275.565 ;
        RECT 793.595 275.395 793.765 275.565 ;
        RECT 794.075 275.395 794.245 275.565 ;
        RECT 794.555 275.395 794.725 275.565 ;
        RECT 795.035 275.395 795.205 275.565 ;
        RECT 795.515 275.395 795.685 275.565 ;
        RECT 795.995 275.395 796.165 275.565 ;
        RECT 595.245 274.875 595.415 275.045 ;
        RECT 595.725 274.875 595.895 275.045 ;
        RECT 596.205 274.875 596.375 275.045 ;
        RECT 601.170 274.905 601.340 275.075 ;
        RECT 355.455 270.405 355.625 270.575 ;
        RECT 355.455 270.045 355.625 270.215 ;
        RECT 355.455 269.685 355.625 269.855 ;
        RECT 355.455 269.325 355.625 269.495 ;
        RECT 355.455 268.965 355.625 269.135 ;
        RECT 355.455 268.605 355.625 268.775 ;
        RECT 355.455 268.245 355.625 268.415 ;
        RECT 355.455 267.885 355.625 268.055 ;
        RECT 355.455 267.525 355.625 267.695 ;
        RECT 355.455 267.165 355.625 267.335 ;
        RECT 355.455 266.805 355.625 266.975 ;
        RECT 271.985 266.500 272.155 266.670 ;
        RECT 272.345 266.500 272.515 266.670 ;
        RECT 275.455 266.500 275.625 266.670 ;
        RECT 275.815 266.500 275.985 266.670 ;
        RECT 278.925 266.500 279.095 266.670 ;
        RECT 279.285 266.500 279.455 266.670 ;
        RECT 282.395 266.500 282.565 266.670 ;
        RECT 282.755 266.500 282.925 266.670 ;
        RECT 285.865 266.500 286.035 266.670 ;
        RECT 286.225 266.500 286.395 266.670 ;
        RECT 355.455 266.445 355.625 266.615 ;
        RECT 211.835 263.220 212.005 263.390 ;
        RECT 212.195 263.220 212.365 263.390 ;
        RECT 215.305 263.220 215.475 263.390 ;
        RECT 215.665 263.220 215.835 263.390 ;
        RECT 218.775 263.220 218.945 263.390 ;
        RECT 219.135 263.220 219.305 263.390 ;
        RECT 222.245 263.220 222.415 263.390 ;
        RECT 222.605 263.220 222.775 263.390 ;
        RECT 225.715 263.220 225.885 263.390 ;
        RECT 226.075 263.220 226.245 263.390 ;
        RECT 231.875 263.210 232.045 263.380 ;
        RECT 232.235 263.210 232.405 263.380 ;
        RECT 235.345 263.210 235.515 263.380 ;
        RECT 235.705 263.210 235.875 263.380 ;
        RECT 238.815 263.210 238.985 263.380 ;
        RECT 239.175 263.210 239.345 263.380 ;
        RECT 242.285 263.210 242.455 263.380 ;
        RECT 242.645 263.210 242.815 263.380 ;
        RECT 245.755 263.210 245.925 263.380 ;
        RECT 246.115 263.210 246.285 263.380 ;
        RECT 251.935 263.210 252.105 263.380 ;
        RECT 252.295 263.210 252.465 263.380 ;
        RECT 255.405 263.210 255.575 263.380 ;
        RECT 255.765 263.210 255.935 263.380 ;
        RECT 258.875 263.210 259.045 263.380 ;
        RECT 259.235 263.210 259.405 263.380 ;
        RECT 262.345 263.210 262.515 263.380 ;
        RECT 262.705 263.210 262.875 263.380 ;
        RECT 265.815 263.210 265.985 263.380 ;
        RECT 266.175 263.210 266.345 263.380 ;
        RECT 271.985 263.210 272.155 263.380 ;
        RECT 272.345 263.210 272.515 263.380 ;
        RECT 275.455 263.210 275.625 263.380 ;
        RECT 275.815 263.210 275.985 263.380 ;
        RECT 278.925 263.210 279.095 263.380 ;
        RECT 279.285 263.210 279.455 263.380 ;
        RECT 282.395 263.210 282.565 263.380 ;
        RECT 282.755 263.210 282.925 263.380 ;
        RECT 285.865 263.210 286.035 263.380 ;
        RECT 286.225 263.210 286.395 263.380 ;
        RECT 214.970 260.160 225.580 261.050 ;
        RECT 234.940 260.160 245.550 261.050 ;
        RECT 255.050 260.160 265.660 261.050 ;
        RECT 275.160 260.160 285.770 261.050 ;
        RECT 355.455 266.085 355.625 266.255 ;
        RECT 355.455 265.725 355.625 265.895 ;
        RECT 355.455 265.365 355.625 265.535 ;
        RECT 355.455 265.005 355.625 265.175 ;
        RECT 355.455 264.645 355.625 264.815 ;
        RECT 355.455 264.285 355.625 264.455 ;
        RECT 355.455 263.925 355.625 264.095 ;
        RECT 355.455 263.565 355.625 263.735 ;
        RECT 355.455 263.205 355.625 263.375 ;
        RECT 355.455 262.845 355.625 263.015 ;
        RECT 355.455 262.485 355.625 262.655 ;
        RECT 288.225 260.260 288.755 261.510 ;
        RECT 355.455 262.125 355.625 262.295 ;
        RECT 355.455 261.765 355.625 261.935 ;
        RECT 355.455 261.405 355.625 261.575 ;
        RECT 355.455 261.045 355.625 261.215 ;
        RECT 355.455 260.685 355.625 260.855 ;
        RECT 355.455 260.325 355.625 260.495 ;
        RECT 355.455 259.965 355.625 260.135 ;
        RECT 355.455 259.605 355.625 259.775 ;
        RECT 211.795 258.680 211.965 258.850 ;
        RECT 212.155 258.680 212.325 258.850 ;
        RECT 215.265 258.680 215.435 258.850 ;
        RECT 215.625 258.680 215.795 258.850 ;
        RECT 218.735 258.680 218.905 258.850 ;
        RECT 219.095 258.680 219.265 258.850 ;
        RECT 222.205 258.680 222.375 258.850 ;
        RECT 222.565 258.680 222.735 258.850 ;
        RECT 225.675 258.680 225.845 258.850 ;
        RECT 226.035 258.680 226.205 258.850 ;
        RECT 231.765 258.680 231.935 258.850 ;
        RECT 232.125 258.680 232.295 258.850 ;
        RECT 235.235 258.680 235.405 258.850 ;
        RECT 235.595 258.680 235.765 258.850 ;
        RECT 238.705 258.680 238.875 258.850 ;
        RECT 239.065 258.680 239.235 258.850 ;
        RECT 242.175 258.680 242.345 258.850 ;
        RECT 242.535 258.680 242.705 258.850 ;
        RECT 245.645 258.680 245.815 258.850 ;
        RECT 246.005 258.680 246.175 258.850 ;
        RECT 251.875 258.680 252.045 258.850 ;
        RECT 252.235 258.680 252.405 258.850 ;
        RECT 255.345 258.680 255.515 258.850 ;
        RECT 255.705 258.680 255.875 258.850 ;
        RECT 258.815 258.680 258.985 258.850 ;
        RECT 259.175 258.680 259.345 258.850 ;
        RECT 262.285 258.680 262.455 258.850 ;
        RECT 262.645 258.680 262.815 258.850 ;
        RECT 265.755 258.680 265.925 258.850 ;
        RECT 266.115 258.680 266.285 258.850 ;
        RECT 271.985 258.680 272.155 258.850 ;
        RECT 272.345 258.680 272.515 258.850 ;
        RECT 275.455 258.680 275.625 258.850 ;
        RECT 275.815 258.680 275.985 258.850 ;
        RECT 278.925 258.680 279.095 258.850 ;
        RECT 279.285 258.680 279.455 258.850 ;
        RECT 282.395 258.680 282.565 258.850 ;
        RECT 282.755 258.680 282.925 258.850 ;
        RECT 285.865 258.680 286.035 258.850 ;
        RECT 286.225 258.680 286.395 258.850 ;
        RECT 355.455 259.245 355.625 259.415 ;
        RECT 355.455 258.885 355.625 259.055 ;
        RECT 211.795 255.390 211.965 255.560 ;
        RECT 212.155 255.390 212.325 255.560 ;
        RECT 215.265 255.390 215.435 255.560 ;
        RECT 215.625 255.390 215.795 255.560 ;
        RECT 218.735 255.390 218.905 255.560 ;
        RECT 219.095 255.390 219.265 255.560 ;
        RECT 222.205 255.390 222.375 255.560 ;
        RECT 222.565 255.390 222.735 255.560 ;
        RECT 225.675 255.390 225.845 255.560 ;
        RECT 226.035 255.390 226.205 255.560 ;
        RECT 97.885 251.600 98.055 251.770 ;
        RECT 98.245 251.600 98.415 251.770 ;
        RECT 101.355 251.600 101.525 251.770 ;
        RECT 101.715 251.600 101.885 251.770 ;
        RECT 97.885 248.310 98.055 248.480 ;
        RECT 98.245 248.310 98.415 248.480 ;
        RECT 101.355 248.310 101.525 248.480 ;
        RECT 101.715 248.310 101.885 248.480 ;
        RECT 84.465 244.800 84.635 244.970 ;
        RECT 84.825 244.800 84.995 244.970 ;
        RECT 87.935 244.800 88.105 244.970 ;
        RECT 88.295 244.800 88.465 244.970 ;
        RECT 91.405 244.800 91.575 244.970 ;
        RECT 91.765 244.800 91.935 244.970 ;
        RECT 84.465 241.510 84.635 241.680 ;
        RECT 84.825 241.510 84.995 241.680 ;
        RECT 87.935 241.510 88.105 241.680 ;
        RECT 88.295 241.510 88.465 241.680 ;
        RECT 91.405 241.510 91.575 241.680 ;
        RECT 91.765 241.510 91.935 241.680 ;
        RECT 94.300 240.970 95.190 242.580 ;
        RECT 231.765 255.390 231.935 255.560 ;
        RECT 232.125 255.390 232.295 255.560 ;
        RECT 235.235 255.390 235.405 255.560 ;
        RECT 235.595 255.390 235.765 255.560 ;
        RECT 238.705 255.390 238.875 255.560 ;
        RECT 239.065 255.390 239.235 255.560 ;
        RECT 242.175 255.390 242.345 255.560 ;
        RECT 242.535 255.390 242.705 255.560 ;
        RECT 245.645 255.390 245.815 255.560 ;
        RECT 246.005 255.390 246.175 255.560 ;
        RECT 211.795 252.100 211.965 252.270 ;
        RECT 212.155 252.100 212.325 252.270 ;
        RECT 215.265 252.100 215.435 252.270 ;
        RECT 215.625 252.100 215.795 252.270 ;
        RECT 218.735 252.100 218.905 252.270 ;
        RECT 219.095 252.100 219.265 252.270 ;
        RECT 222.205 252.100 222.375 252.270 ;
        RECT 222.565 252.100 222.735 252.270 ;
        RECT 225.675 252.100 225.845 252.270 ;
        RECT 226.035 252.100 226.205 252.270 ;
        RECT 211.795 248.810 211.965 248.980 ;
        RECT 212.155 248.810 212.325 248.980 ;
        RECT 215.265 248.810 215.435 248.980 ;
        RECT 215.625 248.810 215.795 248.980 ;
        RECT 218.735 248.810 218.905 248.980 ;
        RECT 219.095 248.810 219.265 248.980 ;
        RECT 222.205 248.810 222.375 248.980 ;
        RECT 222.565 248.810 222.735 248.980 ;
        RECT 225.675 248.810 225.845 248.980 ;
        RECT 226.035 248.810 226.205 248.980 ;
        RECT 97.885 245.020 98.055 245.190 ;
        RECT 98.245 245.020 98.415 245.190 ;
        RECT 101.355 245.020 101.525 245.190 ;
        RECT 101.715 245.020 101.885 245.190 ;
        RECT 103.495 243.470 103.665 243.640 ;
        RECT 251.875 255.390 252.045 255.560 ;
        RECT 252.235 255.390 252.405 255.560 ;
        RECT 255.345 255.390 255.515 255.560 ;
        RECT 255.705 255.390 255.875 255.560 ;
        RECT 258.815 255.390 258.985 255.560 ;
        RECT 259.175 255.390 259.345 255.560 ;
        RECT 262.285 255.390 262.455 255.560 ;
        RECT 262.645 255.390 262.815 255.560 ;
        RECT 265.755 255.390 265.925 255.560 ;
        RECT 266.115 255.390 266.285 255.560 ;
        RECT 231.765 252.100 231.935 252.270 ;
        RECT 232.125 252.100 232.295 252.270 ;
        RECT 235.235 252.100 235.405 252.270 ;
        RECT 235.595 252.100 235.765 252.270 ;
        RECT 238.705 252.100 238.875 252.270 ;
        RECT 239.065 252.100 239.235 252.270 ;
        RECT 242.175 252.100 242.345 252.270 ;
        RECT 242.535 252.100 242.705 252.270 ;
        RECT 245.645 252.100 245.815 252.270 ;
        RECT 246.005 252.100 246.175 252.270 ;
        RECT 231.765 248.810 231.935 248.980 ;
        RECT 232.125 248.810 232.295 248.980 ;
        RECT 235.235 248.810 235.405 248.980 ;
        RECT 235.595 248.810 235.765 248.980 ;
        RECT 238.705 248.810 238.875 248.980 ;
        RECT 239.065 248.810 239.235 248.980 ;
        RECT 242.175 248.810 242.345 248.980 ;
        RECT 242.535 248.810 242.705 248.980 ;
        RECT 245.645 248.810 245.815 248.980 ;
        RECT 246.005 248.810 246.175 248.980 ;
        RECT 211.795 245.520 211.965 245.690 ;
        RECT 212.155 245.520 212.325 245.690 ;
        RECT 215.265 245.520 215.435 245.690 ;
        RECT 215.625 245.520 215.795 245.690 ;
        RECT 218.735 245.520 218.905 245.690 ;
        RECT 219.095 245.520 219.265 245.690 ;
        RECT 222.205 245.520 222.375 245.690 ;
        RECT 222.565 245.520 222.735 245.690 ;
        RECT 225.675 245.520 225.845 245.690 ;
        RECT 226.035 245.520 226.205 245.690 ;
        RECT 271.985 255.390 272.155 255.560 ;
        RECT 272.345 255.390 272.515 255.560 ;
        RECT 275.455 255.390 275.625 255.560 ;
        RECT 275.815 255.390 275.985 255.560 ;
        RECT 278.925 255.390 279.095 255.560 ;
        RECT 279.285 255.390 279.455 255.560 ;
        RECT 282.395 255.390 282.565 255.560 ;
        RECT 282.755 255.390 282.925 255.560 ;
        RECT 285.865 255.390 286.035 255.560 ;
        RECT 286.225 255.390 286.395 255.560 ;
        RECT 251.875 252.100 252.045 252.270 ;
        RECT 252.235 252.100 252.405 252.270 ;
        RECT 255.345 252.100 255.515 252.270 ;
        RECT 255.705 252.100 255.875 252.270 ;
        RECT 258.815 252.100 258.985 252.270 ;
        RECT 259.175 252.100 259.345 252.270 ;
        RECT 262.285 252.100 262.455 252.270 ;
        RECT 262.645 252.100 262.815 252.270 ;
        RECT 265.755 252.100 265.925 252.270 ;
        RECT 266.115 252.100 266.285 252.270 ;
        RECT 251.875 248.810 252.045 248.980 ;
        RECT 252.235 248.810 252.405 248.980 ;
        RECT 255.345 248.810 255.515 248.980 ;
        RECT 255.705 248.810 255.875 248.980 ;
        RECT 258.815 248.810 258.985 248.980 ;
        RECT 259.175 248.810 259.345 248.980 ;
        RECT 262.285 248.810 262.455 248.980 ;
        RECT 262.645 248.810 262.815 248.980 ;
        RECT 265.755 248.810 265.925 248.980 ;
        RECT 266.115 248.810 266.285 248.980 ;
        RECT 231.765 245.520 231.935 245.690 ;
        RECT 232.125 245.520 232.295 245.690 ;
        RECT 235.235 245.520 235.405 245.690 ;
        RECT 235.595 245.520 235.765 245.690 ;
        RECT 238.705 245.520 238.875 245.690 ;
        RECT 239.065 245.520 239.235 245.690 ;
        RECT 242.175 245.520 242.345 245.690 ;
        RECT 242.535 245.520 242.705 245.690 ;
        RECT 245.645 245.520 245.815 245.690 ;
        RECT 246.005 245.520 246.175 245.690 ;
        RECT 355.455 258.525 355.625 258.695 ;
        RECT 355.455 258.165 355.625 258.335 ;
        RECT 355.455 257.805 355.625 257.975 ;
        RECT 356.550 271.005 356.720 271.175 ;
        RECT 356.550 270.645 356.720 270.815 ;
        RECT 356.550 267.535 356.720 267.705 ;
        RECT 356.550 267.175 356.720 267.345 ;
        RECT 356.550 264.065 356.720 264.235 ;
        RECT 356.550 263.705 356.720 263.875 ;
        RECT 356.550 260.595 356.720 260.765 ;
        RECT 356.550 260.235 356.720 260.405 ;
        RECT 356.550 257.125 356.720 257.295 ;
        RECT 359.840 271.005 360.010 271.175 ;
        RECT 359.840 270.645 360.010 270.815 ;
        RECT 359.840 267.535 360.010 267.705 ;
        RECT 359.840 267.175 360.010 267.345 ;
        RECT 359.840 264.065 360.010 264.235 ;
        RECT 359.840 263.705 360.010 263.875 ;
        RECT 359.840 260.595 360.010 260.765 ;
        RECT 359.840 260.235 360.010 260.405 ;
        RECT 359.840 257.125 360.010 257.295 ;
        RECT 356.550 256.765 356.720 256.935 ;
        RECT 363.130 271.005 363.300 271.175 ;
        RECT 363.130 270.645 363.300 270.815 ;
        RECT 363.130 267.535 363.300 267.705 ;
        RECT 363.130 267.175 363.300 267.345 ;
        RECT 363.130 264.065 363.300 264.235 ;
        RECT 363.130 263.705 363.300 263.875 ;
        RECT 363.130 260.595 363.300 260.765 ;
        RECT 363.130 260.235 363.300 260.405 ;
        RECT 363.130 257.125 363.300 257.295 ;
        RECT 366.420 271.005 366.590 271.175 ;
        RECT 369.710 271.005 369.880 271.175 ;
        RECT 366.420 270.645 366.590 270.815 ;
        RECT 366.420 267.535 366.590 267.705 ;
        RECT 366.420 267.175 366.590 267.345 ;
        RECT 366.420 264.065 366.590 264.235 ;
        RECT 366.420 263.705 366.590 263.875 ;
        RECT 366.420 260.595 366.590 260.765 ;
        RECT 366.420 260.235 366.590 260.405 ;
        RECT 366.420 257.125 366.590 257.295 ;
        RECT 369.710 270.645 369.880 270.815 ;
        RECT 369.710 267.535 369.880 267.705 ;
        RECT 369.710 267.175 369.880 267.345 ;
        RECT 369.710 264.065 369.880 264.235 ;
        RECT 369.710 263.705 369.880 263.875 ;
        RECT 369.710 260.595 369.880 260.765 ;
        RECT 369.710 260.235 369.880 260.405 ;
        RECT 359.840 256.765 360.010 256.935 ;
        RECT 363.130 256.765 363.300 256.935 ;
        RECT 366.420 256.765 366.590 256.935 ;
        RECT 369.710 257.125 369.880 257.295 ;
        RECT 374.775 270.305 374.945 270.475 ;
        RECT 374.775 269.945 374.945 270.115 ;
        RECT 374.775 269.585 374.945 269.755 ;
        RECT 374.775 269.225 374.945 269.395 ;
        RECT 374.775 268.865 374.945 269.035 ;
        RECT 374.775 268.505 374.945 268.675 ;
        RECT 374.775 268.145 374.945 268.315 ;
        RECT 374.775 267.785 374.945 267.955 ;
        RECT 374.775 267.425 374.945 267.595 ;
        RECT 374.775 267.065 374.945 267.235 ;
        RECT 374.775 266.705 374.945 266.875 ;
        RECT 374.775 266.345 374.945 266.515 ;
        RECT 374.775 265.985 374.945 266.155 ;
        RECT 374.775 265.625 374.945 265.795 ;
        RECT 374.775 265.265 374.945 265.435 ;
        RECT 374.775 264.905 374.945 265.075 ;
        RECT 374.775 264.545 374.945 264.715 ;
        RECT 374.775 264.185 374.945 264.355 ;
        RECT 374.775 263.825 374.945 263.995 ;
        RECT 374.775 263.465 374.945 263.635 ;
        RECT 374.775 263.105 374.945 263.275 ;
        RECT 374.775 262.745 374.945 262.915 ;
        RECT 374.775 262.385 374.945 262.555 ;
        RECT 374.775 262.025 374.945 262.195 ;
        RECT 374.775 261.665 374.945 261.835 ;
        RECT 374.775 261.305 374.945 261.475 ;
        RECT 374.775 260.945 374.945 261.115 ;
        RECT 374.775 260.585 374.945 260.755 ;
        RECT 374.775 260.225 374.945 260.395 ;
        RECT 374.775 259.865 374.945 260.035 ;
        RECT 374.775 259.505 374.945 259.675 ;
        RECT 374.775 259.145 374.945 259.315 ;
        RECT 374.775 258.785 374.945 258.955 ;
        RECT 374.775 258.425 374.945 258.595 ;
        RECT 374.775 258.065 374.945 258.235 ;
        RECT 374.775 257.705 374.945 257.875 ;
        RECT 375.870 270.905 376.040 271.075 ;
        RECT 375.870 270.545 376.040 270.715 ;
        RECT 375.870 267.435 376.040 267.605 ;
        RECT 375.870 267.075 376.040 267.245 ;
        RECT 375.870 263.965 376.040 264.135 ;
        RECT 375.870 263.605 376.040 263.775 ;
        RECT 375.870 260.495 376.040 260.665 ;
        RECT 375.870 260.135 376.040 260.305 ;
        RECT 375.870 257.025 376.040 257.195 ;
        RECT 382.450 270.905 382.620 271.075 ;
        RECT 389.030 270.905 389.200 271.075 ;
        RECT 382.450 270.545 382.620 270.715 ;
        RECT 382.450 267.435 382.620 267.605 ;
        RECT 382.450 267.075 382.620 267.245 ;
        RECT 382.450 263.965 382.620 264.135 ;
        RECT 382.450 263.605 382.620 263.775 ;
        RECT 382.450 260.495 382.620 260.665 ;
        RECT 382.450 260.135 382.620 260.305 ;
        RECT 382.450 257.025 382.620 257.195 ;
        RECT 369.710 256.765 369.880 256.935 ;
        RECT 389.030 270.545 389.200 270.715 ;
        RECT 389.030 267.435 389.200 267.605 ;
        RECT 389.030 267.075 389.200 267.245 ;
        RECT 389.030 263.965 389.200 264.135 ;
        RECT 389.030 263.605 389.200 263.775 ;
        RECT 389.030 260.495 389.200 260.665 ;
        RECT 389.030 260.135 389.200 260.305 ;
        RECT 389.030 257.025 389.200 257.195 ;
        RECT 375.870 256.665 376.040 256.835 ;
        RECT 382.450 256.665 382.620 256.835 ;
        RECT 394.025 270.375 394.195 270.545 ;
        RECT 394.025 270.015 394.195 270.185 ;
        RECT 394.025 269.655 394.195 269.825 ;
        RECT 394.025 269.295 394.195 269.465 ;
        RECT 394.025 268.935 394.195 269.105 ;
        RECT 394.025 268.575 394.195 268.745 ;
        RECT 394.025 268.215 394.195 268.385 ;
        RECT 394.025 267.855 394.195 268.025 ;
        RECT 394.025 267.495 394.195 267.665 ;
        RECT 394.025 267.135 394.195 267.305 ;
        RECT 394.025 266.775 394.195 266.945 ;
        RECT 394.025 266.415 394.195 266.585 ;
        RECT 394.025 266.055 394.195 266.225 ;
        RECT 394.025 265.695 394.195 265.865 ;
        RECT 394.025 265.335 394.195 265.505 ;
        RECT 394.025 264.975 394.195 265.145 ;
        RECT 394.025 264.615 394.195 264.785 ;
        RECT 394.025 264.255 394.195 264.425 ;
        RECT 394.025 263.895 394.195 264.065 ;
        RECT 394.025 263.535 394.195 263.705 ;
        RECT 394.025 263.175 394.195 263.345 ;
        RECT 394.025 262.815 394.195 262.985 ;
        RECT 394.025 262.455 394.195 262.625 ;
        RECT 394.025 262.095 394.195 262.265 ;
        RECT 394.025 261.735 394.195 261.905 ;
        RECT 394.025 261.375 394.195 261.545 ;
        RECT 394.025 261.015 394.195 261.185 ;
        RECT 394.025 260.655 394.195 260.825 ;
        RECT 394.025 260.295 394.195 260.465 ;
        RECT 394.025 259.935 394.195 260.105 ;
        RECT 394.025 259.575 394.195 259.745 ;
        RECT 394.025 259.215 394.195 259.385 ;
        RECT 394.025 258.855 394.195 259.025 ;
        RECT 394.025 258.495 394.195 258.665 ;
        RECT 394.025 258.135 394.195 258.305 ;
        RECT 394.025 257.775 394.195 257.945 ;
        RECT 395.120 270.975 395.290 271.145 ;
        RECT 395.120 270.615 395.290 270.785 ;
        RECT 395.120 267.505 395.290 267.675 ;
        RECT 395.120 267.145 395.290 267.315 ;
        RECT 395.120 264.035 395.290 264.205 ;
        RECT 395.120 263.675 395.290 263.845 ;
        RECT 395.120 260.565 395.290 260.735 ;
        RECT 395.120 260.205 395.290 260.375 ;
        RECT 395.120 257.095 395.290 257.265 ;
        RECT 398.410 270.975 398.580 271.145 ;
        RECT 398.410 270.615 398.580 270.785 ;
        RECT 398.410 267.505 398.580 267.675 ;
        RECT 398.410 267.145 398.580 267.315 ;
        RECT 398.410 264.035 398.580 264.205 ;
        RECT 398.410 263.675 398.580 263.845 ;
        RECT 398.410 260.565 398.580 260.735 ;
        RECT 398.410 260.205 398.580 260.375 ;
        RECT 398.410 257.095 398.580 257.265 ;
        RECT 389.030 256.665 389.200 256.835 ;
        RECT 395.120 256.735 395.290 256.905 ;
        RECT 401.700 270.975 401.870 271.145 ;
        RECT 401.700 270.615 401.870 270.785 ;
        RECT 401.700 267.505 401.870 267.675 ;
        RECT 401.700 267.145 401.870 267.315 ;
        RECT 401.700 264.035 401.870 264.205 ;
        RECT 401.700 263.675 401.870 263.845 ;
        RECT 401.700 260.565 401.870 260.735 ;
        RECT 401.700 260.205 401.870 260.375 ;
        RECT 401.700 257.095 401.870 257.265 ;
        RECT 404.990 270.975 405.160 271.145 ;
        RECT 408.280 270.975 408.450 271.145 ;
        RECT 409.665 271.245 410.195 274.295 ;
        RECT 595.880 274.395 596.050 274.565 ;
        RECT 596.240 274.395 596.410 274.565 ;
        RECT 602.350 274.885 602.520 275.055 ;
        RECT 603.930 274.885 604.100 275.055 ;
        RECT 605.510 274.885 605.680 275.055 ;
        RECT 606.870 274.895 607.040 275.065 ;
        RECT 608.450 274.895 608.620 275.065 ;
        RECT 610.030 274.895 610.200 275.065 ;
        RECT 611.390 274.895 611.560 275.065 ;
        RECT 612.970 274.895 613.140 275.065 ;
        RECT 614.550 274.895 614.720 275.065 ;
        RECT 615.820 274.875 615.990 275.045 ;
        RECT 617.400 274.875 617.570 275.045 ;
        RECT 618.980 274.875 619.150 275.045 ;
        RECT 620.200 274.885 620.370 275.055 ;
        RECT 621.780 274.885 621.950 275.055 ;
        RECT 623.360 274.885 623.530 275.055 ;
        RECT 624.520 274.875 624.690 275.045 ;
        RECT 626.100 274.875 626.270 275.045 ;
        RECT 627.680 274.875 627.850 275.045 ;
        RECT 628.900 275.135 629.070 275.305 ;
        RECT 628.900 274.775 629.070 274.945 ;
        RECT 635.100 274.845 635.270 275.015 ;
        RECT 635.460 274.845 635.630 275.015 ;
        RECT 639.290 274.935 639.460 275.105 ;
        RECT 639.650 274.935 639.820 275.105 ;
        RECT 643.390 274.915 643.560 275.085 ;
        RECT 643.750 274.915 643.920 275.085 ;
        RECT 781.620 274.915 781.790 275.085 ;
        RECT 781.980 274.915 782.150 275.085 ;
        RECT 760.315 274.330 760.485 274.500 ;
        RECT 784.010 274.915 784.180 275.085 ;
        RECT 786.440 274.915 786.610 275.085 ;
        RECT 786.800 274.915 786.970 275.085 ;
        RECT 787.160 274.915 787.330 275.085 ;
        RECT 788.780 274.915 788.950 275.085 ;
        RECT 789.140 274.915 789.310 275.085 ;
        RECT 789.500 274.915 789.670 275.085 ;
        RECT 791.475 274.915 791.645 275.085 ;
        RECT 791.835 274.915 792.005 275.085 ;
        RECT 792.195 274.915 792.365 275.085 ;
        RECT 793.230 274.915 793.400 275.085 ;
        RECT 793.590 274.915 793.760 275.085 ;
        RECT 793.950 274.915 794.120 275.085 ;
        RECT 794.760 274.915 794.930 275.085 ;
        RECT 795.120 274.915 795.290 275.085 ;
        RECT 795.480 274.915 795.650 275.085 ;
        RECT 800.005 275.385 800.175 275.555 ;
        RECT 800.485 275.385 800.655 275.555 ;
        RECT 800.965 275.385 801.135 275.555 ;
        RECT 801.445 275.385 801.615 275.555 ;
        RECT 801.925 275.385 802.095 275.555 ;
        RECT 802.405 275.385 802.575 275.555 ;
        RECT 802.885 275.385 803.055 275.555 ;
        RECT 803.365 275.385 803.535 275.555 ;
        RECT 803.845 275.385 804.015 275.555 ;
        RECT 804.325 275.385 804.495 275.555 ;
        RECT 804.805 275.385 804.975 275.555 ;
        RECT 805.285 275.385 805.455 275.555 ;
        RECT 805.765 275.385 805.935 275.555 ;
        RECT 806.245 275.385 806.415 275.555 ;
        RECT 806.725 275.385 806.895 275.555 ;
        RECT 807.205 275.385 807.375 275.555 ;
        RECT 807.685 275.385 807.855 275.555 ;
        RECT 808.165 275.385 808.335 275.555 ;
        RECT 808.645 275.385 808.815 275.555 ;
        RECT 809.125 275.385 809.295 275.555 ;
        RECT 809.605 275.385 809.775 275.555 ;
        RECT 810.085 275.385 810.255 275.555 ;
        RECT 810.565 275.385 810.735 275.555 ;
        RECT 811.045 275.385 811.215 275.555 ;
        RECT 811.525 275.385 811.695 275.555 ;
        RECT 812.005 275.385 812.175 275.555 ;
        RECT 812.485 275.385 812.655 275.555 ;
        RECT 812.965 275.385 813.135 275.555 ;
        RECT 813.445 275.385 813.615 275.555 ;
        RECT 813.925 275.385 814.095 275.555 ;
        RECT 814.405 275.385 814.575 275.555 ;
        RECT 814.885 275.385 815.055 275.555 ;
        RECT 800.510 274.905 800.680 275.075 ;
        RECT 800.870 274.905 801.040 275.075 ;
        RECT 802.900 274.905 803.070 275.075 ;
        RECT 805.330 274.905 805.500 275.075 ;
        RECT 805.690 274.905 805.860 275.075 ;
        RECT 806.050 274.905 806.220 275.075 ;
        RECT 807.670 274.905 807.840 275.075 ;
        RECT 808.030 274.905 808.200 275.075 ;
        RECT 808.390 274.905 808.560 275.075 ;
        RECT 810.365 274.905 810.535 275.075 ;
        RECT 810.725 274.905 810.895 275.075 ;
        RECT 811.085 274.905 811.255 275.075 ;
        RECT 812.120 274.905 812.290 275.075 ;
        RECT 812.480 274.905 812.650 275.075 ;
        RECT 812.840 274.905 813.010 275.075 ;
        RECT 813.650 274.905 813.820 275.075 ;
        RECT 814.010 274.905 814.180 275.075 ;
        RECT 814.370 274.905 814.540 275.075 ;
        RECT 818.855 275.355 819.025 275.525 ;
        RECT 819.335 275.355 819.505 275.525 ;
        RECT 819.815 275.355 819.985 275.525 ;
        RECT 820.295 275.355 820.465 275.525 ;
        RECT 820.775 275.355 820.945 275.525 ;
        RECT 821.255 275.355 821.425 275.525 ;
        RECT 821.735 275.355 821.905 275.525 ;
        RECT 822.215 275.355 822.385 275.525 ;
        RECT 822.695 275.355 822.865 275.525 ;
        RECT 823.175 275.355 823.345 275.525 ;
        RECT 823.655 275.355 823.825 275.525 ;
        RECT 824.135 275.355 824.305 275.525 ;
        RECT 824.615 275.355 824.785 275.525 ;
        RECT 825.095 275.355 825.265 275.525 ;
        RECT 825.575 275.355 825.745 275.525 ;
        RECT 826.055 275.355 826.225 275.525 ;
        RECT 826.535 275.355 826.705 275.525 ;
        RECT 827.015 275.355 827.185 275.525 ;
        RECT 827.495 275.355 827.665 275.525 ;
        RECT 827.975 275.355 828.145 275.525 ;
        RECT 828.455 275.355 828.625 275.525 ;
        RECT 828.935 275.355 829.105 275.525 ;
        RECT 829.415 275.355 829.585 275.525 ;
        RECT 829.895 275.355 830.065 275.525 ;
        RECT 830.375 275.355 830.545 275.525 ;
        RECT 830.855 275.355 831.025 275.525 ;
        RECT 831.335 275.355 831.505 275.525 ;
        RECT 831.815 275.355 831.985 275.525 ;
        RECT 832.295 275.355 832.465 275.525 ;
        RECT 832.775 275.355 832.945 275.525 ;
        RECT 833.255 275.355 833.425 275.525 ;
        RECT 833.735 275.355 833.905 275.525 ;
        RECT 819.360 274.875 819.530 275.045 ;
        RECT 819.720 274.875 819.890 275.045 ;
        RECT 821.750 274.875 821.920 275.045 ;
        RECT 824.180 274.875 824.350 275.045 ;
        RECT 824.540 274.875 824.710 275.045 ;
        RECT 824.900 274.875 825.070 275.045 ;
        RECT 826.520 274.875 826.690 275.045 ;
        RECT 826.880 274.875 827.050 275.045 ;
        RECT 827.240 274.875 827.410 275.045 ;
        RECT 829.215 274.875 829.385 275.045 ;
        RECT 829.575 274.875 829.745 275.045 ;
        RECT 829.935 274.875 830.105 275.045 ;
        RECT 830.970 274.875 831.140 275.045 ;
        RECT 831.330 274.875 831.500 275.045 ;
        RECT 831.690 274.875 831.860 275.045 ;
        RECT 832.500 274.875 832.670 275.045 ;
        RECT 832.860 274.875 833.030 275.045 ;
        RECT 833.220 274.875 833.390 275.045 ;
        RECT 838.575 275.395 838.745 275.565 ;
        RECT 839.055 275.395 839.225 275.565 ;
        RECT 839.535 275.395 839.705 275.565 ;
        RECT 840.015 275.395 840.185 275.565 ;
        RECT 840.495 275.395 840.665 275.565 ;
        RECT 840.975 275.395 841.145 275.565 ;
        RECT 841.455 275.395 841.625 275.565 ;
        RECT 841.935 275.395 842.105 275.565 ;
        RECT 856.085 275.345 856.255 275.515 ;
        RECT 856.565 275.345 856.735 275.515 ;
        RECT 857.045 275.345 857.215 275.515 ;
        RECT 857.525 275.345 857.695 275.515 ;
        RECT 858.005 275.345 858.175 275.515 ;
        RECT 858.485 275.345 858.655 275.515 ;
        RECT 858.965 275.345 859.135 275.515 ;
        RECT 839.010 274.915 839.180 275.085 ;
        RECT 839.370 274.915 839.540 275.085 ;
        RECT 839.730 274.915 839.900 275.085 ;
        RECT 840.650 274.915 840.820 275.085 ;
        RECT 841.010 274.915 841.180 275.085 ;
        RECT 841.370 274.915 841.540 275.085 ;
        RECT 856.040 274.865 856.210 275.035 ;
        RECT 856.400 274.865 856.570 275.035 ;
        RECT 856.760 274.865 856.930 275.035 ;
        RECT 857.480 274.865 857.650 275.035 ;
        RECT 857.840 274.865 858.010 275.035 ;
        RECT 858.200 274.865 858.370 275.035 ;
        RECT 858.560 274.865 858.730 275.035 ;
        RECT 844.825 273.135 844.995 273.305 ;
        RECT 845.305 273.135 845.475 273.305 ;
        RECT 845.785 273.135 845.955 273.305 ;
        RECT 846.265 273.135 846.435 273.305 ;
        RECT 846.745 273.135 846.915 273.305 ;
        RECT 847.225 273.135 847.395 273.305 ;
        RECT 847.705 273.135 847.875 273.305 ;
        RECT 850.235 273.145 850.405 273.315 ;
        RECT 850.715 273.145 850.885 273.315 ;
        RECT 851.195 273.145 851.365 273.315 ;
        RECT 844.780 272.655 844.950 272.825 ;
        RECT 845.140 272.655 845.310 272.825 ;
        RECT 845.500 272.655 845.670 272.825 ;
        RECT 846.220 272.655 846.390 272.825 ;
        RECT 846.580 272.655 846.750 272.825 ;
        RECT 846.940 272.655 847.110 272.825 ;
        RECT 847.300 272.655 847.470 272.825 ;
        RECT 850.200 272.665 850.370 272.835 ;
        RECT 850.560 272.665 850.730 272.835 ;
        RECT 861.405 271.955 861.575 272.125 ;
        RECT 861.885 271.955 862.055 272.125 ;
        RECT 862.365 271.955 862.535 272.125 ;
        RECT 862.845 271.955 863.015 272.125 ;
        RECT 863.325 271.955 863.495 272.125 ;
        RECT 863.805 271.955 863.975 272.125 ;
        RECT 864.285 271.955 864.455 272.125 ;
        RECT 862.080 271.475 862.250 271.645 ;
        RECT 862.440 271.475 862.610 271.645 ;
        RECT 862.800 271.475 862.970 271.645 ;
        RECT 863.160 271.475 863.330 271.645 ;
        RECT 863.520 271.475 863.690 271.645 ;
        RECT 863.880 271.475 864.050 271.645 ;
        RECT 404.990 270.615 405.160 270.785 ;
        RECT 404.990 267.505 405.160 267.675 ;
        RECT 404.990 267.145 405.160 267.315 ;
        RECT 404.990 264.035 405.160 264.205 ;
        RECT 404.990 263.675 405.160 263.845 ;
        RECT 404.990 260.565 405.160 260.735 ;
        RECT 404.990 260.205 405.160 260.375 ;
        RECT 404.990 257.095 405.160 257.265 ;
        RECT 408.280 270.615 408.450 270.785 ;
        RECT 680.075 270.875 680.245 271.045 ;
        RECT 680.555 270.875 680.725 271.045 ;
        RECT 681.035 270.875 681.205 271.045 ;
        RECT 681.515 270.875 681.685 271.045 ;
        RECT 681.995 270.875 682.165 271.045 ;
        RECT 682.475 270.875 682.645 271.045 ;
        RECT 682.955 270.875 683.125 271.045 ;
        RECT 685.735 270.885 685.905 271.055 ;
        RECT 686.215 270.885 686.385 271.055 ;
        RECT 686.695 270.885 686.865 271.055 ;
        RECT 687.175 270.885 687.345 271.055 ;
        RECT 687.655 270.885 687.825 271.055 ;
        RECT 688.135 270.885 688.305 271.055 ;
        RECT 688.615 270.885 688.785 271.055 ;
        RECT 680.030 270.395 680.200 270.565 ;
        RECT 680.390 270.395 680.560 270.565 ;
        RECT 680.750 270.395 680.920 270.565 ;
        RECT 681.470 270.395 681.640 270.565 ;
        RECT 681.830 270.395 682.000 270.565 ;
        RECT 682.190 270.395 682.360 270.565 ;
        RECT 682.550 270.395 682.720 270.565 ;
        RECT 685.690 270.405 685.860 270.575 ;
        RECT 686.050 270.405 686.220 270.575 ;
        RECT 686.410 270.405 686.580 270.575 ;
        RECT 687.130 270.405 687.300 270.575 ;
        RECT 687.490 270.405 687.660 270.575 ;
        RECT 687.850 270.405 688.020 270.575 ;
        RECT 688.210 270.405 688.380 270.575 ;
        RECT 691.085 270.905 691.255 271.075 ;
        RECT 691.565 270.905 691.735 271.075 ;
        RECT 692.045 270.905 692.215 271.075 ;
        RECT 692.525 270.905 692.695 271.075 ;
        RECT 693.005 270.905 693.175 271.075 ;
        RECT 693.485 270.905 693.655 271.075 ;
        RECT 693.965 270.905 694.135 271.075 ;
        RECT 697.305 270.895 697.475 271.065 ;
        RECT 697.785 270.895 697.955 271.065 ;
        RECT 698.265 270.895 698.435 271.065 ;
        RECT 698.745 270.895 698.915 271.065 ;
        RECT 699.225 270.895 699.395 271.065 ;
        RECT 699.705 270.895 699.875 271.065 ;
        RECT 700.185 270.895 700.355 271.065 ;
        RECT 691.760 270.425 691.930 270.595 ;
        RECT 692.120 270.425 692.290 270.595 ;
        RECT 692.480 270.425 692.650 270.595 ;
        RECT 692.840 270.425 693.010 270.595 ;
        RECT 693.200 270.425 693.370 270.595 ;
        RECT 693.560 270.425 693.730 270.595 ;
        RECT 697.260 270.415 697.430 270.585 ;
        RECT 697.620 270.415 697.790 270.585 ;
        RECT 697.980 270.415 698.150 270.585 ;
        RECT 698.700 270.415 698.870 270.585 ;
        RECT 699.060 270.415 699.230 270.585 ;
        RECT 699.420 270.415 699.590 270.585 ;
        RECT 699.780 270.415 699.950 270.585 ;
        RECT 702.965 270.905 703.135 271.075 ;
        RECT 703.445 270.905 703.615 271.075 ;
        RECT 703.925 270.905 704.095 271.075 ;
        RECT 704.405 270.905 704.575 271.075 ;
        RECT 704.885 270.905 705.055 271.075 ;
        RECT 705.365 270.905 705.535 271.075 ;
        RECT 705.845 270.905 706.015 271.075 ;
        RECT 708.315 270.925 708.485 271.095 ;
        RECT 708.795 270.925 708.965 271.095 ;
        RECT 709.275 270.925 709.445 271.095 ;
        RECT 709.755 270.925 709.925 271.095 ;
        RECT 710.235 270.925 710.405 271.095 ;
        RECT 710.715 270.925 710.885 271.095 ;
        RECT 711.195 270.925 711.365 271.095 ;
        RECT 714.875 270.995 715.045 271.165 ;
        RECT 715.355 270.995 715.525 271.165 ;
        RECT 715.835 270.995 716.005 271.165 ;
        RECT 716.315 270.995 716.485 271.165 ;
        RECT 716.795 270.995 716.965 271.165 ;
        RECT 717.275 270.995 717.445 271.165 ;
        RECT 717.755 270.995 717.925 271.165 ;
        RECT 702.920 270.425 703.090 270.595 ;
        RECT 703.280 270.425 703.450 270.595 ;
        RECT 703.640 270.425 703.810 270.595 ;
        RECT 704.360 270.425 704.530 270.595 ;
        RECT 704.720 270.425 704.890 270.595 ;
        RECT 705.080 270.425 705.250 270.595 ;
        RECT 705.440 270.425 705.610 270.595 ;
        RECT 708.990 270.445 709.160 270.615 ;
        RECT 709.350 270.445 709.520 270.615 ;
        RECT 709.710 270.445 709.880 270.615 ;
        RECT 710.070 270.445 710.240 270.615 ;
        RECT 710.430 270.445 710.600 270.615 ;
        RECT 710.790 270.445 710.960 270.615 ;
        RECT 714.830 270.515 715.000 270.685 ;
        RECT 715.190 270.515 715.360 270.685 ;
        RECT 715.550 270.515 715.720 270.685 ;
        RECT 716.270 270.515 716.440 270.685 ;
        RECT 716.630 270.515 716.800 270.685 ;
        RECT 716.990 270.515 717.160 270.685 ;
        RECT 717.350 270.515 717.520 270.685 ;
        RECT 720.535 271.005 720.705 271.175 ;
        RECT 721.015 271.005 721.185 271.175 ;
        RECT 721.495 271.005 721.665 271.175 ;
        RECT 721.975 271.005 722.145 271.175 ;
        RECT 722.455 271.005 722.625 271.175 ;
        RECT 722.935 271.005 723.105 271.175 ;
        RECT 723.415 271.005 723.585 271.175 ;
        RECT 725.885 271.025 726.055 271.195 ;
        RECT 726.365 271.025 726.535 271.195 ;
        RECT 726.845 271.025 727.015 271.195 ;
        RECT 727.325 271.025 727.495 271.195 ;
        RECT 727.805 271.025 727.975 271.195 ;
        RECT 728.285 271.025 728.455 271.195 ;
        RECT 728.765 271.025 728.935 271.195 ;
        RECT 732.045 271.025 732.215 271.195 ;
        RECT 732.525 271.025 732.695 271.195 ;
        RECT 733.005 271.025 733.175 271.195 ;
        RECT 733.485 271.025 733.655 271.195 ;
        RECT 733.965 271.025 734.135 271.195 ;
        RECT 734.445 271.025 734.615 271.195 ;
        RECT 734.925 271.025 735.095 271.195 ;
        RECT 720.490 270.525 720.660 270.695 ;
        RECT 720.850 270.525 721.020 270.695 ;
        RECT 721.210 270.525 721.380 270.695 ;
        RECT 721.930 270.525 722.100 270.695 ;
        RECT 722.290 270.525 722.460 270.695 ;
        RECT 722.650 270.525 722.820 270.695 ;
        RECT 723.010 270.525 723.180 270.695 ;
        RECT 726.560 270.545 726.730 270.715 ;
        RECT 726.920 270.545 727.090 270.715 ;
        RECT 727.280 270.545 727.450 270.715 ;
        RECT 727.640 270.545 727.810 270.715 ;
        RECT 728.000 270.545 728.170 270.715 ;
        RECT 728.360 270.545 728.530 270.715 ;
        RECT 732.000 270.545 732.170 270.715 ;
        RECT 732.360 270.545 732.530 270.715 ;
        RECT 732.720 270.545 732.890 270.715 ;
        RECT 733.440 270.545 733.610 270.715 ;
        RECT 733.800 270.545 733.970 270.715 ;
        RECT 734.160 270.545 734.330 270.715 ;
        RECT 734.520 270.545 734.690 270.715 ;
        RECT 737.705 271.035 737.875 271.205 ;
        RECT 738.185 271.035 738.355 271.205 ;
        RECT 738.665 271.035 738.835 271.205 ;
        RECT 739.145 271.035 739.315 271.205 ;
        RECT 739.625 271.035 739.795 271.205 ;
        RECT 740.105 271.035 740.275 271.205 ;
        RECT 740.585 271.035 740.755 271.205 ;
        RECT 743.055 271.055 743.225 271.225 ;
        RECT 743.535 271.055 743.705 271.225 ;
        RECT 744.015 271.055 744.185 271.225 ;
        RECT 744.495 271.055 744.665 271.225 ;
        RECT 744.975 271.055 745.145 271.225 ;
        RECT 745.455 271.055 745.625 271.225 ;
        RECT 745.935 271.055 746.105 271.225 ;
        RECT 749.855 271.085 750.025 271.255 ;
        RECT 750.335 271.085 750.505 271.255 ;
        RECT 750.815 271.085 750.985 271.255 ;
        RECT 751.295 271.085 751.465 271.255 ;
        RECT 751.775 271.085 751.945 271.255 ;
        RECT 752.255 271.085 752.425 271.255 ;
        RECT 752.735 271.085 752.905 271.255 ;
        RECT 737.660 270.555 737.830 270.725 ;
        RECT 738.020 270.555 738.190 270.725 ;
        RECT 738.380 270.555 738.550 270.725 ;
        RECT 739.100 270.555 739.270 270.725 ;
        RECT 739.460 270.555 739.630 270.725 ;
        RECT 739.820 270.555 739.990 270.725 ;
        RECT 740.180 270.555 740.350 270.725 ;
        RECT 743.730 270.575 743.900 270.745 ;
        RECT 744.090 270.575 744.260 270.745 ;
        RECT 744.450 270.575 744.620 270.745 ;
        RECT 744.810 270.575 744.980 270.745 ;
        RECT 745.170 270.575 745.340 270.745 ;
        RECT 745.530 270.575 745.700 270.745 ;
        RECT 749.810 270.605 749.980 270.775 ;
        RECT 750.170 270.605 750.340 270.775 ;
        RECT 750.530 270.605 750.700 270.775 ;
        RECT 751.250 270.605 751.420 270.775 ;
        RECT 751.610 270.605 751.780 270.775 ;
        RECT 751.970 270.605 752.140 270.775 ;
        RECT 752.330 270.605 752.500 270.775 ;
        RECT 755.515 271.095 755.685 271.265 ;
        RECT 755.995 271.095 756.165 271.265 ;
        RECT 756.475 271.095 756.645 271.265 ;
        RECT 756.955 271.095 757.125 271.265 ;
        RECT 757.435 271.095 757.605 271.265 ;
        RECT 757.915 271.095 758.085 271.265 ;
        RECT 758.395 271.095 758.565 271.265 ;
        RECT 760.865 271.115 761.035 271.285 ;
        RECT 761.345 271.115 761.515 271.285 ;
        RECT 761.825 271.115 761.995 271.285 ;
        RECT 762.305 271.115 762.475 271.285 ;
        RECT 762.785 271.115 762.955 271.285 ;
        RECT 763.265 271.115 763.435 271.285 ;
        RECT 763.745 271.115 763.915 271.285 ;
        RECT 755.470 270.615 755.640 270.785 ;
        RECT 755.830 270.615 756.000 270.785 ;
        RECT 756.190 270.615 756.360 270.785 ;
        RECT 756.910 270.615 757.080 270.785 ;
        RECT 757.270 270.615 757.440 270.785 ;
        RECT 757.630 270.615 757.800 270.785 ;
        RECT 757.990 270.615 758.160 270.785 ;
        RECT 761.540 270.635 761.710 270.805 ;
        RECT 761.900 270.635 762.070 270.805 ;
        RECT 762.260 270.635 762.430 270.805 ;
        RECT 762.620 270.635 762.790 270.805 ;
        RECT 762.980 270.635 763.150 270.805 ;
        RECT 763.340 270.635 763.510 270.805 ;
        RECT 838.585 269.835 838.755 270.005 ;
        RECT 839.065 269.835 839.235 270.005 ;
        RECT 839.545 269.835 839.715 270.005 ;
        RECT 840.025 269.835 840.195 270.005 ;
        RECT 840.505 269.835 840.675 270.005 ;
        RECT 840.985 269.835 841.155 270.005 ;
        RECT 841.465 269.835 841.635 270.005 ;
        RECT 838.540 269.355 838.710 269.525 ;
        RECT 838.900 269.355 839.070 269.525 ;
        RECT 839.260 269.355 839.430 269.525 ;
        RECT 756.555 268.445 756.725 268.615 ;
        RECT 756.555 268.085 756.725 268.255 ;
        RECT 839.980 269.355 840.150 269.525 ;
        RECT 840.340 269.355 840.510 269.525 ;
        RECT 840.700 269.355 840.870 269.525 ;
        RECT 841.060 269.355 841.230 269.525 ;
        RECT 856.165 268.675 856.335 268.845 ;
        RECT 856.645 268.675 856.815 268.845 ;
        RECT 857.125 268.675 857.295 268.845 ;
        RECT 857.605 268.675 857.775 268.845 ;
        RECT 858.085 268.675 858.255 268.845 ;
        RECT 858.565 268.675 858.735 268.845 ;
        RECT 859.045 268.675 859.215 268.845 ;
        RECT 856.120 268.195 856.290 268.365 ;
        RECT 856.480 268.195 856.650 268.365 ;
        RECT 856.840 268.195 857.010 268.365 ;
        RECT 781.125 267.835 781.295 268.005 ;
        RECT 781.605 267.835 781.775 268.005 ;
        RECT 782.085 267.835 782.255 268.005 ;
        RECT 782.565 267.835 782.735 268.005 ;
        RECT 783.045 267.835 783.215 268.005 ;
        RECT 783.525 267.835 783.695 268.005 ;
        RECT 784.005 267.835 784.175 268.005 ;
        RECT 784.485 267.835 784.655 268.005 ;
        RECT 784.965 267.835 785.135 268.005 ;
        RECT 785.445 267.835 785.615 268.005 ;
        RECT 785.925 267.835 786.095 268.005 ;
        RECT 786.405 267.835 786.575 268.005 ;
        RECT 786.885 267.835 787.055 268.005 ;
        RECT 787.365 267.835 787.535 268.005 ;
        RECT 787.845 267.835 788.015 268.005 ;
        RECT 788.325 267.835 788.495 268.005 ;
        RECT 788.805 267.835 788.975 268.005 ;
        RECT 789.285 267.835 789.455 268.005 ;
        RECT 789.765 267.835 789.935 268.005 ;
        RECT 790.245 267.835 790.415 268.005 ;
        RECT 790.725 267.835 790.895 268.005 ;
        RECT 791.205 267.835 791.375 268.005 ;
        RECT 791.685 267.835 791.855 268.005 ;
        RECT 792.165 267.835 792.335 268.005 ;
        RECT 792.645 267.835 792.815 268.005 ;
        RECT 793.125 267.835 793.295 268.005 ;
        RECT 793.605 267.835 793.775 268.005 ;
        RECT 794.085 267.835 794.255 268.005 ;
        RECT 794.565 267.835 794.735 268.005 ;
        RECT 795.045 267.835 795.215 268.005 ;
        RECT 795.525 267.835 795.695 268.005 ;
        RECT 796.005 267.835 796.175 268.005 ;
        RECT 408.280 267.505 408.450 267.675 ;
        RECT 408.280 267.145 408.450 267.315 ;
        RECT 781.630 267.355 781.800 267.525 ;
        RECT 781.990 267.355 782.160 267.525 ;
        RECT 784.020 267.355 784.190 267.525 ;
        RECT 786.450 267.355 786.620 267.525 ;
        RECT 786.810 267.355 786.980 267.525 ;
        RECT 787.170 267.355 787.340 267.525 ;
        RECT 788.790 267.355 788.960 267.525 ;
        RECT 789.150 267.355 789.320 267.525 ;
        RECT 789.510 267.355 789.680 267.525 ;
        RECT 791.485 267.355 791.655 267.525 ;
        RECT 791.845 267.355 792.015 267.525 ;
        RECT 792.205 267.355 792.375 267.525 ;
        RECT 793.240 267.355 793.410 267.525 ;
        RECT 793.600 267.355 793.770 267.525 ;
        RECT 793.960 267.355 794.130 267.525 ;
        RECT 794.770 267.355 794.940 267.525 ;
        RECT 795.130 267.355 795.300 267.525 ;
        RECT 795.490 267.355 795.660 267.525 ;
        RECT 799.655 267.895 799.825 268.065 ;
        RECT 800.135 267.895 800.305 268.065 ;
        RECT 800.615 267.895 800.785 268.065 ;
        RECT 801.095 267.895 801.265 268.065 ;
        RECT 801.575 267.895 801.745 268.065 ;
        RECT 802.055 267.895 802.225 268.065 ;
        RECT 802.535 267.895 802.705 268.065 ;
        RECT 803.015 267.895 803.185 268.065 ;
        RECT 803.495 267.895 803.665 268.065 ;
        RECT 803.975 267.895 804.145 268.065 ;
        RECT 804.455 267.895 804.625 268.065 ;
        RECT 804.935 267.895 805.105 268.065 ;
        RECT 805.415 267.895 805.585 268.065 ;
        RECT 805.895 267.895 806.065 268.065 ;
        RECT 806.375 267.895 806.545 268.065 ;
        RECT 806.855 267.895 807.025 268.065 ;
        RECT 807.335 267.895 807.505 268.065 ;
        RECT 807.815 267.895 807.985 268.065 ;
        RECT 808.295 267.895 808.465 268.065 ;
        RECT 808.775 267.895 808.945 268.065 ;
        RECT 809.255 267.895 809.425 268.065 ;
        RECT 809.735 267.895 809.905 268.065 ;
        RECT 810.215 267.895 810.385 268.065 ;
        RECT 810.695 267.895 810.865 268.065 ;
        RECT 811.175 267.895 811.345 268.065 ;
        RECT 811.655 267.895 811.825 268.065 ;
        RECT 812.135 267.895 812.305 268.065 ;
        RECT 812.615 267.895 812.785 268.065 ;
        RECT 813.095 267.895 813.265 268.065 ;
        RECT 813.575 267.895 813.745 268.065 ;
        RECT 814.055 267.895 814.225 268.065 ;
        RECT 814.535 267.895 814.705 268.065 ;
        RECT 800.160 267.415 800.330 267.585 ;
        RECT 800.520 267.415 800.690 267.585 ;
        RECT 802.550 267.415 802.720 267.585 ;
        RECT 804.980 267.415 805.150 267.585 ;
        RECT 805.340 267.415 805.510 267.585 ;
        RECT 805.700 267.415 805.870 267.585 ;
        RECT 807.320 267.415 807.490 267.585 ;
        RECT 807.680 267.415 807.850 267.585 ;
        RECT 808.040 267.415 808.210 267.585 ;
        RECT 810.015 267.415 810.185 267.585 ;
        RECT 810.375 267.415 810.545 267.585 ;
        RECT 810.735 267.415 810.905 267.585 ;
        RECT 811.770 267.415 811.940 267.585 ;
        RECT 812.130 267.415 812.300 267.585 ;
        RECT 812.490 267.415 812.660 267.585 ;
        RECT 813.300 267.415 813.470 267.585 ;
        RECT 813.660 267.415 813.830 267.585 ;
        RECT 814.020 267.415 814.190 267.585 ;
        RECT 857.560 268.195 857.730 268.365 ;
        RECT 857.920 268.195 858.090 268.365 ;
        RECT 858.280 268.195 858.450 268.365 ;
        RECT 858.640 268.195 858.810 268.365 ;
        RECT 408.280 264.035 408.450 264.205 ;
        RECT 408.280 263.675 408.450 263.845 ;
        RECT 408.280 260.565 408.450 260.735 ;
        RECT 679.525 260.685 679.695 260.855 ;
        RECT 680.005 260.685 680.175 260.855 ;
        RECT 680.485 260.685 680.655 260.855 ;
        RECT 680.965 260.685 681.135 260.855 ;
        RECT 681.445 260.685 681.615 260.855 ;
        RECT 681.925 260.685 682.095 260.855 ;
        RECT 682.405 260.685 682.575 260.855 ;
        RECT 682.885 260.685 683.055 260.855 ;
        RECT 683.365 260.685 683.535 260.855 ;
        RECT 683.845 260.685 684.015 260.855 ;
        RECT 684.325 260.685 684.495 260.855 ;
        RECT 408.280 260.205 408.450 260.375 ;
        RECT 679.930 260.205 680.100 260.375 ;
        RECT 680.290 260.205 680.460 260.375 ;
        RECT 680.650 260.205 680.820 260.375 ;
        RECT 681.010 260.205 681.180 260.375 ;
        RECT 681.370 260.205 681.540 260.375 ;
        RECT 681.730 260.205 681.900 260.375 ;
        RECT 682.455 260.205 682.625 260.375 ;
        RECT 682.815 260.205 682.985 260.375 ;
        RECT 683.175 260.205 683.345 260.375 ;
        RECT 683.535 260.205 683.705 260.375 ;
        RECT 683.895 260.205 684.065 260.375 ;
        RECT 696.805 260.695 696.975 260.865 ;
        RECT 697.285 260.695 697.455 260.865 ;
        RECT 697.765 260.695 697.935 260.865 ;
        RECT 698.245 260.695 698.415 260.865 ;
        RECT 698.725 260.695 698.895 260.865 ;
        RECT 699.205 260.695 699.375 260.865 ;
        RECT 699.685 260.695 699.855 260.865 ;
        RECT 700.165 260.695 700.335 260.865 ;
        RECT 700.645 260.695 700.815 260.865 ;
        RECT 701.125 260.695 701.295 260.865 ;
        RECT 701.605 260.695 701.775 260.865 ;
        RECT 697.210 260.215 697.380 260.385 ;
        RECT 697.570 260.215 697.740 260.385 ;
        RECT 697.930 260.215 698.100 260.385 ;
        RECT 698.290 260.215 698.460 260.385 ;
        RECT 698.650 260.215 698.820 260.385 ;
        RECT 699.010 260.215 699.180 260.385 ;
        RECT 699.735 260.215 699.905 260.385 ;
        RECT 700.095 260.215 700.265 260.385 ;
        RECT 700.455 260.215 700.625 260.385 ;
        RECT 700.815 260.215 700.985 260.385 ;
        RECT 701.175 260.215 701.345 260.385 ;
        RECT 714.575 260.695 714.745 260.865 ;
        RECT 715.055 260.695 715.225 260.865 ;
        RECT 715.535 260.695 715.705 260.865 ;
        RECT 716.015 260.695 716.185 260.865 ;
        RECT 716.495 260.695 716.665 260.865 ;
        RECT 716.975 260.695 717.145 260.865 ;
        RECT 717.455 260.695 717.625 260.865 ;
        RECT 717.935 260.695 718.105 260.865 ;
        RECT 718.415 260.695 718.585 260.865 ;
        RECT 718.895 260.695 719.065 260.865 ;
        RECT 719.375 260.695 719.545 260.865 ;
        RECT 714.980 260.215 715.150 260.385 ;
        RECT 715.340 260.215 715.510 260.385 ;
        RECT 715.700 260.215 715.870 260.385 ;
        RECT 716.060 260.215 716.230 260.385 ;
        RECT 716.420 260.215 716.590 260.385 ;
        RECT 716.780 260.215 716.950 260.385 ;
        RECT 717.505 260.215 717.675 260.385 ;
        RECT 717.865 260.215 718.035 260.385 ;
        RECT 718.225 260.215 718.395 260.385 ;
        RECT 718.585 260.215 718.755 260.385 ;
        RECT 718.945 260.215 719.115 260.385 ;
        RECT 731.815 260.695 731.985 260.865 ;
        RECT 732.295 260.695 732.465 260.865 ;
        RECT 732.775 260.695 732.945 260.865 ;
        RECT 733.255 260.695 733.425 260.865 ;
        RECT 733.735 260.695 733.905 260.865 ;
        RECT 734.215 260.695 734.385 260.865 ;
        RECT 734.695 260.695 734.865 260.865 ;
        RECT 735.175 260.695 735.345 260.865 ;
        RECT 735.655 260.695 735.825 260.865 ;
        RECT 736.135 260.695 736.305 260.865 ;
        RECT 736.615 260.695 736.785 260.865 ;
        RECT 732.220 260.215 732.390 260.385 ;
        RECT 732.580 260.215 732.750 260.385 ;
        RECT 732.940 260.215 733.110 260.385 ;
        RECT 733.300 260.215 733.470 260.385 ;
        RECT 733.660 260.215 733.830 260.385 ;
        RECT 734.020 260.215 734.190 260.385 ;
        RECT 749.295 260.705 749.465 260.875 ;
        RECT 749.775 260.705 749.945 260.875 ;
        RECT 750.255 260.705 750.425 260.875 ;
        RECT 750.735 260.705 750.905 260.875 ;
        RECT 751.215 260.705 751.385 260.875 ;
        RECT 751.695 260.705 751.865 260.875 ;
        RECT 752.175 260.705 752.345 260.875 ;
        RECT 752.655 260.705 752.825 260.875 ;
        RECT 753.135 260.705 753.305 260.875 ;
        RECT 753.615 260.705 753.785 260.875 ;
        RECT 754.095 260.705 754.265 260.875 ;
        RECT 734.745 260.215 734.915 260.385 ;
        RECT 735.105 260.215 735.275 260.385 ;
        RECT 735.465 260.215 735.635 260.385 ;
        RECT 735.825 260.215 735.995 260.385 ;
        RECT 736.185 260.215 736.355 260.385 ;
        RECT 749.700 260.225 749.870 260.395 ;
        RECT 750.060 260.225 750.230 260.395 ;
        RECT 750.420 260.225 750.590 260.395 ;
        RECT 750.780 260.225 750.950 260.395 ;
        RECT 751.140 260.225 751.310 260.395 ;
        RECT 751.500 260.225 751.670 260.395 ;
        RECT 752.225 260.225 752.395 260.395 ;
        RECT 752.585 260.225 752.755 260.395 ;
        RECT 752.945 260.225 753.115 260.395 ;
        RECT 753.305 260.225 753.475 260.395 ;
        RECT 753.665 260.225 753.835 260.395 ;
        RECT 856.035 259.365 856.205 259.535 ;
        RECT 856.515 259.365 856.685 259.535 ;
        RECT 856.995 259.365 857.165 259.535 ;
        RECT 857.475 259.365 857.645 259.535 ;
        RECT 857.955 259.365 858.125 259.535 ;
        RECT 858.435 259.365 858.605 259.535 ;
        RECT 858.915 259.365 859.085 259.535 ;
        RECT 601.020 258.615 601.190 258.785 ;
        RECT 602.200 258.625 602.370 258.795 ;
        RECT 603.780 258.625 603.950 258.795 ;
        RECT 605.360 258.625 605.530 258.795 ;
        RECT 606.720 258.635 606.890 258.805 ;
        RECT 608.300 258.635 608.470 258.805 ;
        RECT 609.880 258.635 610.050 258.805 ;
        RECT 611.240 258.635 611.410 258.805 ;
        RECT 612.820 258.635 612.990 258.805 ;
        RECT 614.400 258.635 614.570 258.805 ;
        RECT 615.670 258.615 615.840 258.785 ;
        RECT 617.250 258.615 617.420 258.785 ;
        RECT 618.830 258.615 619.000 258.785 ;
        RECT 620.050 258.625 620.220 258.795 ;
        RECT 621.630 258.625 621.800 258.795 ;
        RECT 623.210 258.625 623.380 258.795 ;
        RECT 624.370 258.615 624.540 258.785 ;
        RECT 625.950 258.615 626.120 258.785 ;
        RECT 627.530 258.615 627.700 258.785 ;
        RECT 628.750 258.845 628.920 259.015 ;
        RECT 601.020 258.255 601.190 258.425 ;
        RECT 601.020 257.895 601.190 258.065 ;
        RECT 601.020 257.535 601.190 257.705 ;
        RECT 628.750 258.485 628.920 258.655 ;
        RECT 628.750 258.125 628.920 258.295 ;
        RECT 628.750 257.765 628.920 257.935 ;
        RECT 855.990 258.885 856.160 259.055 ;
        RECT 856.350 258.885 856.520 259.055 ;
        RECT 856.710 258.885 856.880 259.055 ;
        RECT 634.985 257.595 635.155 257.765 ;
        RECT 635.465 257.595 635.635 257.765 ;
        RECT 635.945 257.595 636.115 257.765 ;
        RECT 639.175 257.685 639.345 257.855 ;
        RECT 639.655 257.685 639.825 257.855 ;
        RECT 640.135 257.685 640.305 257.855 ;
        RECT 643.275 257.665 643.445 257.835 ;
        RECT 643.755 257.665 643.925 257.835 ;
        RECT 644.235 257.665 644.405 257.835 ;
        RECT 857.430 258.885 857.600 259.055 ;
        RECT 857.790 258.885 857.960 259.055 ;
        RECT 858.150 258.885 858.320 259.055 ;
        RECT 858.510 258.885 858.680 259.055 ;
        RECT 398.410 256.735 398.580 256.905 ;
        RECT 401.700 256.735 401.870 256.905 ;
        RECT 404.990 256.735 405.160 256.905 ;
        RECT 408.280 257.095 408.450 257.265 ;
        RECT 595.095 257.145 595.265 257.315 ;
        RECT 595.575 257.145 595.745 257.315 ;
        RECT 596.055 257.145 596.225 257.315 ;
        RECT 601.020 257.175 601.190 257.345 ;
        RECT 408.280 256.735 408.450 256.905 ;
        RECT 595.730 256.665 595.900 256.835 ;
        RECT 596.090 256.665 596.260 256.835 ;
        RECT 602.200 257.155 602.370 257.325 ;
        RECT 603.780 257.155 603.950 257.325 ;
        RECT 605.360 257.155 605.530 257.325 ;
        RECT 606.720 257.165 606.890 257.335 ;
        RECT 608.300 257.165 608.470 257.335 ;
        RECT 609.880 257.165 610.050 257.335 ;
        RECT 611.240 257.165 611.410 257.335 ;
        RECT 612.820 257.165 612.990 257.335 ;
        RECT 614.400 257.165 614.570 257.335 ;
        RECT 615.670 257.145 615.840 257.315 ;
        RECT 617.250 257.145 617.420 257.315 ;
        RECT 618.830 257.145 619.000 257.315 ;
        RECT 620.050 257.155 620.220 257.325 ;
        RECT 621.630 257.155 621.800 257.325 ;
        RECT 623.210 257.155 623.380 257.325 ;
        RECT 624.370 257.145 624.540 257.315 ;
        RECT 625.950 257.145 626.120 257.315 ;
        RECT 627.530 257.145 627.700 257.315 ;
        RECT 628.750 257.405 628.920 257.575 ;
        RECT 628.750 257.045 628.920 257.215 ;
        RECT 634.950 257.115 635.120 257.285 ;
        RECT 635.310 257.115 635.480 257.285 ;
        RECT 639.140 257.205 639.310 257.375 ;
        RECT 639.500 257.205 639.670 257.375 ;
        RECT 643.240 257.185 643.410 257.355 ;
        RECT 643.600 257.185 643.770 257.355 ;
        RECT 861.345 256.875 861.515 257.045 ;
        RECT 861.825 256.875 861.995 257.045 ;
        RECT 862.305 256.875 862.475 257.045 ;
        RECT 862.785 256.875 862.955 257.045 ;
        RECT 863.265 256.875 863.435 257.045 ;
        RECT 863.745 256.875 863.915 257.045 ;
        RECT 864.225 256.875 864.395 257.045 ;
        RECT 862.020 256.395 862.190 256.565 ;
        RECT 862.380 256.395 862.550 256.565 ;
        RECT 862.740 256.395 862.910 256.565 ;
        RECT 863.100 256.395 863.270 256.565 ;
        RECT 863.460 256.395 863.630 256.565 ;
        RECT 863.820 256.395 863.990 256.565 ;
        RECT 679.935 255.025 680.105 255.195 ;
        RECT 680.415 255.025 680.585 255.195 ;
        RECT 680.895 255.025 681.065 255.195 ;
        RECT 681.375 255.025 681.545 255.195 ;
        RECT 681.855 255.025 682.025 255.195 ;
        RECT 682.335 255.025 682.505 255.195 ;
        RECT 682.815 255.025 682.985 255.195 ;
        RECT 683.295 255.025 683.465 255.195 ;
        RECT 683.775 255.025 683.945 255.195 ;
        RECT 684.255 255.025 684.425 255.195 ;
        RECT 684.735 255.025 684.905 255.195 ;
        RECT 680.340 254.545 680.510 254.715 ;
        RECT 680.700 254.545 680.870 254.715 ;
        RECT 681.060 254.545 681.230 254.715 ;
        RECT 681.420 254.545 681.590 254.715 ;
        RECT 681.780 254.545 681.950 254.715 ;
        RECT 682.140 254.545 682.310 254.715 ;
        RECT 682.865 254.545 683.035 254.715 ;
        RECT 683.225 254.545 683.395 254.715 ;
        RECT 683.585 254.545 683.755 254.715 ;
        RECT 683.945 254.545 684.115 254.715 ;
        RECT 684.305 254.545 684.475 254.715 ;
        RECT 687.175 254.985 687.345 255.155 ;
        RECT 687.655 254.985 687.825 255.155 ;
        RECT 688.135 254.985 688.305 255.155 ;
        RECT 688.615 254.985 688.785 255.155 ;
        RECT 689.095 254.985 689.265 255.155 ;
        RECT 689.575 254.985 689.745 255.155 ;
        RECT 690.055 254.985 690.225 255.155 ;
        RECT 690.535 254.985 690.705 255.155 ;
        RECT 691.015 254.985 691.185 255.155 ;
        RECT 691.495 254.985 691.665 255.155 ;
        RECT 691.975 254.985 692.145 255.155 ;
        RECT 697.165 255.045 697.335 255.215 ;
        RECT 697.645 255.045 697.815 255.215 ;
        RECT 698.125 255.045 698.295 255.215 ;
        RECT 698.605 255.045 698.775 255.215 ;
        RECT 699.085 255.045 699.255 255.215 ;
        RECT 699.565 255.045 699.735 255.215 ;
        RECT 700.045 255.045 700.215 255.215 ;
        RECT 700.525 255.045 700.695 255.215 ;
        RECT 701.005 255.045 701.175 255.215 ;
        RECT 701.485 255.045 701.655 255.215 ;
        RECT 701.965 255.045 702.135 255.215 ;
        RECT 687.580 254.505 687.750 254.675 ;
        RECT 687.940 254.505 688.110 254.675 ;
        RECT 688.300 254.505 688.470 254.675 ;
        RECT 688.660 254.505 688.830 254.675 ;
        RECT 689.020 254.505 689.190 254.675 ;
        RECT 689.380 254.505 689.550 254.675 ;
        RECT 690.105 254.505 690.275 254.675 ;
        RECT 690.465 254.505 690.635 254.675 ;
        RECT 690.825 254.505 690.995 254.675 ;
        RECT 691.185 254.505 691.355 254.675 ;
        RECT 691.545 254.505 691.715 254.675 ;
        RECT 697.570 254.565 697.740 254.735 ;
        RECT 697.930 254.565 698.100 254.735 ;
        RECT 698.290 254.565 698.460 254.735 ;
        RECT 698.650 254.565 698.820 254.735 ;
        RECT 699.010 254.565 699.180 254.735 ;
        RECT 699.370 254.565 699.540 254.735 ;
        RECT 700.095 254.565 700.265 254.735 ;
        RECT 700.455 254.565 700.625 254.735 ;
        RECT 700.815 254.565 700.985 254.735 ;
        RECT 701.175 254.565 701.345 254.735 ;
        RECT 701.535 254.565 701.705 254.735 ;
        RECT 704.405 255.005 704.575 255.175 ;
        RECT 704.885 255.005 705.055 255.175 ;
        RECT 705.365 255.005 705.535 255.175 ;
        RECT 705.845 255.005 706.015 255.175 ;
        RECT 706.325 255.005 706.495 255.175 ;
        RECT 706.805 255.005 706.975 255.175 ;
        RECT 707.285 255.005 707.455 255.175 ;
        RECT 707.765 255.005 707.935 255.175 ;
        RECT 708.245 255.005 708.415 255.175 ;
        RECT 708.725 255.005 708.895 255.175 ;
        RECT 709.205 255.005 709.375 255.175 ;
        RECT 714.735 255.145 714.905 255.315 ;
        RECT 715.215 255.145 715.385 255.315 ;
        RECT 715.695 255.145 715.865 255.315 ;
        RECT 716.175 255.145 716.345 255.315 ;
        RECT 716.655 255.145 716.825 255.315 ;
        RECT 717.135 255.145 717.305 255.315 ;
        RECT 717.615 255.145 717.785 255.315 ;
        RECT 718.095 255.145 718.265 255.315 ;
        RECT 718.575 255.145 718.745 255.315 ;
        RECT 719.055 255.145 719.225 255.315 ;
        RECT 719.535 255.145 719.705 255.315 ;
        RECT 704.810 254.525 704.980 254.695 ;
        RECT 705.170 254.525 705.340 254.695 ;
        RECT 705.530 254.525 705.700 254.695 ;
        RECT 705.890 254.525 706.060 254.695 ;
        RECT 706.250 254.525 706.420 254.695 ;
        RECT 706.610 254.525 706.780 254.695 ;
        RECT 707.335 254.525 707.505 254.695 ;
        RECT 707.695 254.525 707.865 254.695 ;
        RECT 708.055 254.525 708.225 254.695 ;
        RECT 708.415 254.525 708.585 254.695 ;
        RECT 708.775 254.525 708.945 254.695 ;
        RECT 715.140 254.665 715.310 254.835 ;
        RECT 715.500 254.665 715.670 254.835 ;
        RECT 715.860 254.665 716.030 254.835 ;
        RECT 716.220 254.665 716.390 254.835 ;
        RECT 716.580 254.665 716.750 254.835 ;
        RECT 716.940 254.665 717.110 254.835 ;
        RECT 717.665 254.665 717.835 254.835 ;
        RECT 718.025 254.665 718.195 254.835 ;
        RECT 718.385 254.665 718.555 254.835 ;
        RECT 718.745 254.665 718.915 254.835 ;
        RECT 719.105 254.665 719.275 254.835 ;
        RECT 721.975 255.105 722.145 255.275 ;
        RECT 722.455 255.105 722.625 255.275 ;
        RECT 722.935 255.105 723.105 255.275 ;
        RECT 723.415 255.105 723.585 255.275 ;
        RECT 723.895 255.105 724.065 255.275 ;
        RECT 724.375 255.105 724.545 255.275 ;
        RECT 724.855 255.105 725.025 255.275 ;
        RECT 725.335 255.105 725.505 255.275 ;
        RECT 725.815 255.105 725.985 255.275 ;
        RECT 726.295 255.105 726.465 255.275 ;
        RECT 726.775 255.105 726.945 255.275 ;
        RECT 731.905 255.175 732.075 255.345 ;
        RECT 732.385 255.175 732.555 255.345 ;
        RECT 732.865 255.175 733.035 255.345 ;
        RECT 733.345 255.175 733.515 255.345 ;
        RECT 733.825 255.175 733.995 255.345 ;
        RECT 734.305 255.175 734.475 255.345 ;
        RECT 734.785 255.175 734.955 255.345 ;
        RECT 735.265 255.175 735.435 255.345 ;
        RECT 735.745 255.175 735.915 255.345 ;
        RECT 736.225 255.175 736.395 255.345 ;
        RECT 736.705 255.175 736.875 255.345 ;
        RECT 722.380 254.625 722.550 254.795 ;
        RECT 722.740 254.625 722.910 254.795 ;
        RECT 723.100 254.625 723.270 254.795 ;
        RECT 723.460 254.625 723.630 254.795 ;
        RECT 723.820 254.625 723.990 254.795 ;
        RECT 724.180 254.625 724.350 254.795 ;
        RECT 724.905 254.625 725.075 254.795 ;
        RECT 725.265 254.625 725.435 254.795 ;
        RECT 725.625 254.625 725.795 254.795 ;
        RECT 725.985 254.625 726.155 254.795 ;
        RECT 726.345 254.625 726.515 254.795 ;
        RECT 732.310 254.695 732.480 254.865 ;
        RECT 732.670 254.695 732.840 254.865 ;
        RECT 733.030 254.695 733.200 254.865 ;
        RECT 733.390 254.695 733.560 254.865 ;
        RECT 733.750 254.695 733.920 254.865 ;
        RECT 734.110 254.695 734.280 254.865 ;
        RECT 734.835 254.695 735.005 254.865 ;
        RECT 735.195 254.695 735.365 254.865 ;
        RECT 735.555 254.695 735.725 254.865 ;
        RECT 735.915 254.695 736.085 254.865 ;
        RECT 736.275 254.695 736.445 254.865 ;
        RECT 739.145 255.135 739.315 255.305 ;
        RECT 739.625 255.135 739.795 255.305 ;
        RECT 740.105 255.135 740.275 255.305 ;
        RECT 740.585 255.135 740.755 255.305 ;
        RECT 741.065 255.135 741.235 255.305 ;
        RECT 741.545 255.135 741.715 255.305 ;
        RECT 742.025 255.135 742.195 255.305 ;
        RECT 742.505 255.135 742.675 255.305 ;
        RECT 742.985 255.135 743.155 255.305 ;
        RECT 743.465 255.135 743.635 255.305 ;
        RECT 743.945 255.135 744.115 255.305 ;
        RECT 749.715 255.235 749.885 255.405 ;
        RECT 750.195 255.235 750.365 255.405 ;
        RECT 750.675 255.235 750.845 255.405 ;
        RECT 751.155 255.235 751.325 255.405 ;
        RECT 751.635 255.235 751.805 255.405 ;
        RECT 752.115 255.235 752.285 255.405 ;
        RECT 752.595 255.235 752.765 255.405 ;
        RECT 753.075 255.235 753.245 255.405 ;
        RECT 753.555 255.235 753.725 255.405 ;
        RECT 754.035 255.235 754.205 255.405 ;
        RECT 754.515 255.235 754.685 255.405 ;
        RECT 739.550 254.655 739.720 254.825 ;
        RECT 739.910 254.655 740.080 254.825 ;
        RECT 740.270 254.655 740.440 254.825 ;
        RECT 740.630 254.655 740.800 254.825 ;
        RECT 740.990 254.655 741.160 254.825 ;
        RECT 741.350 254.655 741.520 254.825 ;
        RECT 742.075 254.655 742.245 254.825 ;
        RECT 742.435 254.655 742.605 254.825 ;
        RECT 742.795 254.655 742.965 254.825 ;
        RECT 743.155 254.655 743.325 254.825 ;
        RECT 743.515 254.655 743.685 254.825 ;
        RECT 750.120 254.755 750.290 254.925 ;
        RECT 750.480 254.755 750.650 254.925 ;
        RECT 750.840 254.755 751.010 254.925 ;
        RECT 751.200 254.755 751.370 254.925 ;
        RECT 751.560 254.755 751.730 254.925 ;
        RECT 751.920 254.755 752.090 254.925 ;
        RECT 752.645 254.755 752.815 254.925 ;
        RECT 753.005 254.755 753.175 254.925 ;
        RECT 753.365 254.755 753.535 254.925 ;
        RECT 753.725 254.755 753.895 254.925 ;
        RECT 754.085 254.755 754.255 254.925 ;
        RECT 756.955 255.195 757.125 255.365 ;
        RECT 757.435 255.195 757.605 255.365 ;
        RECT 757.915 255.195 758.085 255.365 ;
        RECT 758.395 255.195 758.565 255.365 ;
        RECT 758.875 255.195 759.045 255.365 ;
        RECT 759.355 255.195 759.525 255.365 ;
        RECT 759.835 255.195 760.005 255.365 ;
        RECT 760.315 255.195 760.485 255.365 ;
        RECT 760.795 255.195 760.965 255.365 ;
        RECT 761.275 255.195 761.445 255.365 ;
        RECT 761.755 255.195 761.925 255.365 ;
        RECT 757.360 254.715 757.530 254.885 ;
        RECT 757.720 254.715 757.890 254.885 ;
        RECT 758.080 254.715 758.250 254.885 ;
        RECT 758.440 254.715 758.610 254.885 ;
        RECT 758.800 254.715 758.970 254.885 ;
        RECT 759.160 254.715 759.330 254.885 ;
        RECT 759.885 254.715 760.055 254.885 ;
        RECT 760.245 254.715 760.415 254.885 ;
        RECT 760.605 254.715 760.775 254.885 ;
        RECT 760.965 254.715 761.135 254.885 ;
        RECT 761.325 254.715 761.495 254.885 ;
        RECT 856.095 253.595 856.265 253.765 ;
        RECT 856.575 253.595 856.745 253.765 ;
        RECT 857.055 253.595 857.225 253.765 ;
        RECT 857.535 253.595 857.705 253.765 ;
        RECT 858.015 253.595 858.185 253.765 ;
        RECT 858.495 253.595 858.665 253.765 ;
        RECT 858.975 253.595 859.145 253.765 ;
        RECT 699.095 253.000 699.265 253.170 ;
        RECT 856.050 253.115 856.220 253.285 ;
        RECT 856.410 253.115 856.580 253.285 ;
        RECT 856.770 253.115 856.940 253.285 ;
        RECT 271.985 252.100 272.155 252.270 ;
        RECT 272.345 252.100 272.515 252.270 ;
        RECT 275.455 252.100 275.625 252.270 ;
        RECT 275.815 252.100 275.985 252.270 ;
        RECT 278.925 252.100 279.095 252.270 ;
        RECT 279.285 252.100 279.455 252.270 ;
        RECT 282.395 252.100 282.565 252.270 ;
        RECT 282.755 252.100 282.925 252.270 ;
        RECT 285.865 252.100 286.035 252.270 ;
        RECT 286.225 252.100 286.395 252.270 ;
        RECT 271.985 248.810 272.155 248.980 ;
        RECT 272.345 248.810 272.515 248.980 ;
        RECT 275.455 248.810 275.625 248.980 ;
        RECT 275.815 248.810 275.985 248.980 ;
        RECT 278.925 248.810 279.095 248.980 ;
        RECT 279.285 248.810 279.455 248.980 ;
        RECT 282.395 248.810 282.565 248.980 ;
        RECT 282.755 248.810 282.925 248.980 ;
        RECT 285.865 248.810 286.035 248.980 ;
        RECT 286.225 248.810 286.395 248.980 ;
        RECT 251.875 245.520 252.045 245.690 ;
        RECT 252.235 245.520 252.405 245.690 ;
        RECT 255.345 245.520 255.515 245.690 ;
        RECT 255.705 245.520 255.875 245.690 ;
        RECT 258.815 245.520 258.985 245.690 ;
        RECT 259.175 245.520 259.345 245.690 ;
        RECT 262.285 245.520 262.455 245.690 ;
        RECT 262.645 245.520 262.815 245.690 ;
        RECT 265.755 245.520 265.925 245.690 ;
        RECT 266.115 245.520 266.285 245.690 ;
        RECT 857.490 253.115 857.660 253.285 ;
        RECT 857.850 253.115 858.020 253.285 ;
        RECT 858.210 253.115 858.380 253.285 ;
        RECT 858.570 253.115 858.740 253.285 ;
        RECT 680.055 249.345 680.225 249.515 ;
        RECT 680.535 249.345 680.705 249.515 ;
        RECT 681.015 249.345 681.185 249.515 ;
        RECT 681.495 249.345 681.665 249.515 ;
        RECT 681.975 249.345 682.145 249.515 ;
        RECT 682.455 249.345 682.625 249.515 ;
        RECT 682.935 249.345 683.105 249.515 ;
        RECT 680.010 248.865 680.180 249.035 ;
        RECT 680.370 248.865 680.540 249.035 ;
        RECT 680.730 248.865 680.900 249.035 ;
        RECT 681.450 248.865 681.620 249.035 ;
        RECT 681.810 248.865 681.980 249.035 ;
        RECT 682.170 248.865 682.340 249.035 ;
        RECT 682.530 248.865 682.700 249.035 ;
        RECT 685.715 249.355 685.885 249.525 ;
        RECT 686.195 249.355 686.365 249.525 ;
        RECT 686.675 249.355 686.845 249.525 ;
        RECT 687.155 249.355 687.325 249.525 ;
        RECT 687.635 249.355 687.805 249.525 ;
        RECT 688.115 249.355 688.285 249.525 ;
        RECT 688.595 249.355 688.765 249.525 ;
        RECT 691.065 249.375 691.235 249.545 ;
        RECT 691.545 249.375 691.715 249.545 ;
        RECT 692.025 249.375 692.195 249.545 ;
        RECT 692.505 249.375 692.675 249.545 ;
        RECT 692.985 249.375 693.155 249.545 ;
        RECT 693.465 249.375 693.635 249.545 ;
        RECT 693.945 249.375 694.115 249.545 ;
        RECT 697.285 249.365 697.455 249.535 ;
        RECT 697.765 249.365 697.935 249.535 ;
        RECT 698.245 249.365 698.415 249.535 ;
        RECT 698.725 249.365 698.895 249.535 ;
        RECT 699.205 249.365 699.375 249.535 ;
        RECT 699.685 249.365 699.855 249.535 ;
        RECT 700.165 249.365 700.335 249.535 ;
        RECT 685.670 248.875 685.840 249.045 ;
        RECT 686.030 248.875 686.200 249.045 ;
        RECT 686.390 248.875 686.560 249.045 ;
        RECT 687.110 248.875 687.280 249.045 ;
        RECT 687.470 248.875 687.640 249.045 ;
        RECT 687.830 248.875 688.000 249.045 ;
        RECT 688.190 248.875 688.360 249.045 ;
        RECT 691.740 248.895 691.910 249.065 ;
        RECT 692.100 248.895 692.270 249.065 ;
        RECT 692.460 248.895 692.630 249.065 ;
        RECT 692.820 248.895 692.990 249.065 ;
        RECT 693.180 248.895 693.350 249.065 ;
        RECT 693.540 248.895 693.710 249.065 ;
        RECT 697.240 248.885 697.410 249.055 ;
        RECT 697.600 248.885 697.770 249.055 ;
        RECT 697.960 248.885 698.130 249.055 ;
        RECT 698.680 248.885 698.850 249.055 ;
        RECT 699.040 248.885 699.210 249.055 ;
        RECT 699.400 248.885 699.570 249.055 ;
        RECT 699.760 248.885 699.930 249.055 ;
        RECT 702.945 249.375 703.115 249.545 ;
        RECT 703.425 249.375 703.595 249.545 ;
        RECT 703.905 249.375 704.075 249.545 ;
        RECT 704.385 249.375 704.555 249.545 ;
        RECT 704.865 249.375 705.035 249.545 ;
        RECT 705.345 249.375 705.515 249.545 ;
        RECT 705.825 249.375 705.995 249.545 ;
        RECT 708.295 249.395 708.465 249.565 ;
        RECT 708.775 249.395 708.945 249.565 ;
        RECT 709.255 249.395 709.425 249.565 ;
        RECT 709.735 249.395 709.905 249.565 ;
        RECT 710.215 249.395 710.385 249.565 ;
        RECT 710.695 249.395 710.865 249.565 ;
        RECT 711.175 249.395 711.345 249.565 ;
        RECT 714.855 249.465 715.025 249.635 ;
        RECT 715.335 249.465 715.505 249.635 ;
        RECT 715.815 249.465 715.985 249.635 ;
        RECT 716.295 249.465 716.465 249.635 ;
        RECT 716.775 249.465 716.945 249.635 ;
        RECT 717.255 249.465 717.425 249.635 ;
        RECT 717.735 249.465 717.905 249.635 ;
        RECT 702.900 248.895 703.070 249.065 ;
        RECT 703.260 248.895 703.430 249.065 ;
        RECT 703.620 248.895 703.790 249.065 ;
        RECT 704.340 248.895 704.510 249.065 ;
        RECT 704.700 248.895 704.870 249.065 ;
        RECT 705.060 248.895 705.230 249.065 ;
        RECT 705.420 248.895 705.590 249.065 ;
        RECT 708.970 248.915 709.140 249.085 ;
        RECT 709.330 248.915 709.500 249.085 ;
        RECT 709.690 248.915 709.860 249.085 ;
        RECT 710.050 248.915 710.220 249.085 ;
        RECT 710.410 248.915 710.580 249.085 ;
        RECT 710.770 248.915 710.940 249.085 ;
        RECT 714.810 248.985 714.980 249.155 ;
        RECT 715.170 248.985 715.340 249.155 ;
        RECT 715.530 248.985 715.700 249.155 ;
        RECT 716.250 248.985 716.420 249.155 ;
        RECT 716.610 248.985 716.780 249.155 ;
        RECT 716.970 248.985 717.140 249.155 ;
        RECT 717.330 248.985 717.500 249.155 ;
        RECT 720.515 249.475 720.685 249.645 ;
        RECT 720.995 249.475 721.165 249.645 ;
        RECT 721.475 249.475 721.645 249.645 ;
        RECT 721.955 249.475 722.125 249.645 ;
        RECT 722.435 249.475 722.605 249.645 ;
        RECT 722.915 249.475 723.085 249.645 ;
        RECT 723.395 249.475 723.565 249.645 ;
        RECT 725.865 249.495 726.035 249.665 ;
        RECT 726.345 249.495 726.515 249.665 ;
        RECT 726.825 249.495 726.995 249.665 ;
        RECT 727.305 249.495 727.475 249.665 ;
        RECT 727.785 249.495 727.955 249.665 ;
        RECT 728.265 249.495 728.435 249.665 ;
        RECT 728.745 249.495 728.915 249.665 ;
        RECT 732.025 249.495 732.195 249.665 ;
        RECT 732.505 249.495 732.675 249.665 ;
        RECT 732.985 249.495 733.155 249.665 ;
        RECT 733.465 249.495 733.635 249.665 ;
        RECT 733.945 249.495 734.115 249.665 ;
        RECT 734.425 249.495 734.595 249.665 ;
        RECT 734.905 249.495 735.075 249.665 ;
        RECT 720.470 248.995 720.640 249.165 ;
        RECT 720.830 248.995 721.000 249.165 ;
        RECT 721.190 248.995 721.360 249.165 ;
        RECT 721.910 248.995 722.080 249.165 ;
        RECT 722.270 248.995 722.440 249.165 ;
        RECT 722.630 248.995 722.800 249.165 ;
        RECT 722.990 248.995 723.160 249.165 ;
        RECT 726.540 249.015 726.710 249.185 ;
        RECT 726.900 249.015 727.070 249.185 ;
        RECT 727.260 249.015 727.430 249.185 ;
        RECT 727.620 249.015 727.790 249.185 ;
        RECT 727.980 249.015 728.150 249.185 ;
        RECT 728.340 249.015 728.510 249.185 ;
        RECT 731.980 249.015 732.150 249.185 ;
        RECT 732.340 249.015 732.510 249.185 ;
        RECT 732.700 249.015 732.870 249.185 ;
        RECT 733.420 249.015 733.590 249.185 ;
        RECT 733.780 249.015 733.950 249.185 ;
        RECT 734.140 249.015 734.310 249.185 ;
        RECT 734.500 249.015 734.670 249.185 ;
        RECT 737.685 249.505 737.855 249.675 ;
        RECT 738.165 249.505 738.335 249.675 ;
        RECT 738.645 249.505 738.815 249.675 ;
        RECT 739.125 249.505 739.295 249.675 ;
        RECT 739.605 249.505 739.775 249.675 ;
        RECT 740.085 249.505 740.255 249.675 ;
        RECT 740.565 249.505 740.735 249.675 ;
        RECT 743.035 249.525 743.205 249.695 ;
        RECT 743.515 249.525 743.685 249.695 ;
        RECT 743.995 249.525 744.165 249.695 ;
        RECT 744.475 249.525 744.645 249.695 ;
        RECT 744.955 249.525 745.125 249.695 ;
        RECT 745.435 249.525 745.605 249.695 ;
        RECT 745.915 249.525 746.085 249.695 ;
        RECT 749.835 249.555 750.005 249.725 ;
        RECT 750.315 249.555 750.485 249.725 ;
        RECT 750.795 249.555 750.965 249.725 ;
        RECT 751.275 249.555 751.445 249.725 ;
        RECT 751.755 249.555 751.925 249.725 ;
        RECT 752.235 249.555 752.405 249.725 ;
        RECT 752.715 249.555 752.885 249.725 ;
        RECT 737.640 249.025 737.810 249.195 ;
        RECT 738.000 249.025 738.170 249.195 ;
        RECT 738.360 249.025 738.530 249.195 ;
        RECT 739.080 249.025 739.250 249.195 ;
        RECT 739.440 249.025 739.610 249.195 ;
        RECT 739.800 249.025 739.970 249.195 ;
        RECT 740.160 249.025 740.330 249.195 ;
        RECT 743.710 249.045 743.880 249.215 ;
        RECT 744.070 249.045 744.240 249.215 ;
        RECT 744.430 249.045 744.600 249.215 ;
        RECT 744.790 249.045 744.960 249.215 ;
        RECT 745.150 249.045 745.320 249.215 ;
        RECT 745.510 249.045 745.680 249.215 ;
        RECT 749.790 249.075 749.960 249.245 ;
        RECT 750.150 249.075 750.320 249.245 ;
        RECT 750.510 249.075 750.680 249.245 ;
        RECT 751.230 249.075 751.400 249.245 ;
        RECT 751.590 249.075 751.760 249.245 ;
        RECT 751.950 249.075 752.120 249.245 ;
        RECT 752.310 249.075 752.480 249.245 ;
        RECT 755.495 249.565 755.665 249.735 ;
        RECT 755.975 249.565 756.145 249.735 ;
        RECT 756.455 249.565 756.625 249.735 ;
        RECT 756.935 249.565 757.105 249.735 ;
        RECT 757.415 249.565 757.585 249.735 ;
        RECT 757.895 249.565 758.065 249.735 ;
        RECT 758.375 249.565 758.545 249.735 ;
        RECT 760.845 249.585 761.015 249.755 ;
        RECT 761.325 249.585 761.495 249.755 ;
        RECT 761.805 249.585 761.975 249.755 ;
        RECT 762.285 249.585 762.455 249.755 ;
        RECT 762.765 249.585 762.935 249.755 ;
        RECT 763.245 249.585 763.415 249.755 ;
        RECT 763.725 249.585 763.895 249.755 ;
        RECT 755.450 249.085 755.620 249.255 ;
        RECT 755.810 249.085 755.980 249.255 ;
        RECT 756.170 249.085 756.340 249.255 ;
        RECT 756.890 249.085 757.060 249.255 ;
        RECT 757.250 249.085 757.420 249.255 ;
        RECT 757.610 249.085 757.780 249.255 ;
        RECT 757.970 249.085 758.140 249.255 ;
        RECT 761.520 249.105 761.690 249.275 ;
        RECT 761.880 249.105 762.050 249.275 ;
        RECT 762.240 249.105 762.410 249.275 ;
        RECT 762.600 249.105 762.770 249.275 ;
        RECT 762.960 249.105 763.130 249.275 ;
        RECT 763.320 249.105 763.490 249.275 ;
        RECT 697.355 246.830 697.525 247.000 ;
        RECT 271.985 245.520 272.155 245.690 ;
        RECT 272.345 245.520 272.515 245.690 ;
        RECT 275.455 245.520 275.625 245.690 ;
        RECT 275.815 245.520 275.985 245.690 ;
        RECT 278.925 245.520 279.095 245.690 ;
        RECT 279.285 245.520 279.455 245.690 ;
        RECT 282.395 245.520 282.565 245.690 ;
        RECT 282.755 245.520 282.925 245.690 ;
        RECT 285.865 245.520 286.035 245.690 ;
        RECT 286.225 245.520 286.395 245.690 ;
        RECT 211.795 242.230 211.965 242.400 ;
        RECT 212.155 242.230 212.325 242.400 ;
        RECT 215.265 242.230 215.435 242.400 ;
        RECT 215.625 242.230 215.795 242.400 ;
        RECT 218.735 242.230 218.905 242.400 ;
        RECT 219.095 242.230 219.265 242.400 ;
        RECT 222.205 242.230 222.375 242.400 ;
        RECT 222.565 242.230 222.735 242.400 ;
        RECT 225.675 242.230 225.845 242.400 ;
        RECT 226.035 242.230 226.205 242.400 ;
        RECT 231.765 242.230 231.935 242.400 ;
        RECT 232.125 242.230 232.295 242.400 ;
        RECT 235.235 242.230 235.405 242.400 ;
        RECT 235.595 242.230 235.765 242.400 ;
        RECT 238.705 242.230 238.875 242.400 ;
        RECT 239.065 242.230 239.235 242.400 ;
        RECT 242.175 242.230 242.345 242.400 ;
        RECT 242.535 242.230 242.705 242.400 ;
        RECT 245.645 242.230 245.815 242.400 ;
        RECT 246.005 242.230 246.175 242.400 ;
        RECT 251.875 242.230 252.045 242.400 ;
        RECT 252.235 242.230 252.405 242.400 ;
        RECT 255.345 242.230 255.515 242.400 ;
        RECT 255.705 242.230 255.875 242.400 ;
        RECT 258.815 242.230 258.985 242.400 ;
        RECT 259.175 242.230 259.345 242.400 ;
        RECT 262.285 242.230 262.455 242.400 ;
        RECT 262.645 242.230 262.815 242.400 ;
        RECT 265.755 242.230 265.925 242.400 ;
        RECT 266.115 242.230 266.285 242.400 ;
        RECT 271.985 242.230 272.155 242.400 ;
        RECT 272.345 242.230 272.515 242.400 ;
        RECT 275.455 242.230 275.625 242.400 ;
        RECT 275.815 242.230 275.985 242.400 ;
        RECT 278.925 242.230 279.095 242.400 ;
        RECT 279.285 242.230 279.455 242.400 ;
        RECT 282.395 242.230 282.565 242.400 ;
        RECT 282.755 242.230 282.925 242.400 ;
        RECT 285.865 242.230 286.035 242.400 ;
        RECT 286.225 242.230 286.395 242.400 ;
        RECT 97.885 241.730 98.055 241.900 ;
        RECT 98.245 241.730 98.415 241.900 ;
        RECT 101.355 241.730 101.525 241.900 ;
        RECT 101.715 241.730 101.885 241.900 ;
        RECT 214.380 240.000 223.910 240.530 ;
        RECT 234.415 239.970 246.105 240.500 ;
        RECT 254.345 239.835 266.035 240.365 ;
        RECT 272.865 239.790 285.275 240.680 ;
        RECT 97.885 238.440 98.055 238.610 ;
        RECT 98.245 238.440 98.415 238.610 ;
        RECT 101.355 238.440 101.525 238.610 ;
        RECT 101.715 238.440 101.885 238.610 ;
        RECT 4.855 238.190 5.025 238.360 ;
        RECT 5.215 238.190 5.385 238.360 ;
        RECT 8.325 238.190 8.495 238.360 ;
        RECT 8.685 238.190 8.855 238.360 ;
        RECT 11.795 238.190 11.965 238.360 ;
        RECT 12.155 238.190 12.325 238.360 ;
        RECT 18.195 238.170 18.365 238.340 ;
        RECT 18.555 238.170 18.725 238.340 ;
        RECT 21.665 238.170 21.835 238.340 ;
        RECT 22.025 238.170 22.195 238.340 ;
        RECT 25.135 238.170 25.305 238.340 ;
        RECT 25.495 238.170 25.665 238.340 ;
        RECT 31.565 238.200 31.735 238.370 ;
        RECT 31.925 238.200 32.095 238.370 ;
        RECT 35.035 238.200 35.205 238.370 ;
        RECT 35.395 238.200 35.565 238.370 ;
        RECT 38.505 238.200 38.675 238.370 ;
        RECT 38.865 238.200 39.035 238.370 ;
        RECT 44.795 238.200 44.965 238.370 ;
        RECT 45.155 238.200 45.325 238.370 ;
        RECT 48.265 238.200 48.435 238.370 ;
        RECT 48.625 238.200 48.795 238.370 ;
        RECT 51.735 238.200 51.905 238.370 ;
        RECT 52.095 238.200 52.265 238.370 ;
        RECT 58.065 238.170 58.235 238.340 ;
        RECT 58.425 238.170 58.595 238.340 ;
        RECT 61.535 238.170 61.705 238.340 ;
        RECT 61.895 238.170 62.065 238.340 ;
        RECT 65.005 238.170 65.175 238.340 ;
        RECT 65.365 238.170 65.535 238.340 ;
        RECT 71.335 238.200 71.505 238.370 ;
        RECT 71.695 238.200 71.865 238.370 ;
        RECT 74.805 238.200 74.975 238.370 ;
        RECT 75.165 238.200 75.335 238.370 ;
        RECT 78.275 238.200 78.445 238.370 ;
        RECT 78.635 238.200 78.805 238.370 ;
        RECT 84.465 238.220 84.635 238.390 ;
        RECT 84.825 238.220 84.995 238.390 ;
        RECT 87.935 238.220 88.105 238.390 ;
        RECT 88.295 238.220 88.465 238.390 ;
        RECT 91.405 238.220 91.575 238.390 ;
        RECT 91.765 238.220 91.935 238.390 ;
        RECT 13.705 236.395 13.875 236.565 ;
        RECT 14.065 236.395 14.235 236.565 ;
        RECT 14.425 236.395 14.595 236.565 ;
        RECT 14.785 236.395 14.955 236.565 ;
        RECT 15.145 236.395 15.315 236.565 ;
        RECT 15.505 236.395 15.675 236.565 ;
        RECT 15.865 236.395 16.035 236.565 ;
        RECT 16.225 236.395 16.395 236.565 ;
        RECT 16.585 236.395 16.755 236.565 ;
        RECT 16.945 236.395 17.115 236.565 ;
        RECT 17.305 236.395 17.475 236.565 ;
        RECT 17.665 236.395 17.835 236.565 ;
        RECT 18.025 236.395 18.195 236.565 ;
        RECT 18.385 236.395 18.555 236.565 ;
        RECT 18.745 236.395 18.915 236.565 ;
        RECT 19.105 236.395 19.275 236.565 ;
        RECT 19.465 236.395 19.635 236.565 ;
        RECT 19.825 236.395 19.995 236.565 ;
        RECT 20.185 236.395 20.355 236.565 ;
        RECT 20.545 236.395 20.715 236.565 ;
        RECT 20.905 236.395 21.075 236.565 ;
        RECT 21.265 236.395 21.435 236.565 ;
        RECT -51.765 236.080 -51.595 236.250 ;
        RECT -50.475 236.080 -50.305 236.250 ;
        RECT -49.185 236.080 -49.015 236.250 ;
        RECT -47.895 236.080 -47.725 236.250 ;
        RECT -46.605 236.080 -46.435 236.250 ;
        RECT -45.315 236.080 -45.145 236.250 ;
        RECT -44.025 236.080 -43.855 236.250 ;
        RECT -42.735 236.080 -42.565 236.250 ;
        RECT -41.445 236.080 -41.275 236.250 ;
        RECT -40.155 236.080 -39.985 236.250 ;
        RECT -38.865 236.080 -38.695 236.250 ;
        RECT -37.575 236.080 -37.405 236.250 ;
        RECT -36.285 236.080 -36.115 236.250 ;
        RECT -34.995 236.080 -34.825 236.250 ;
        RECT -33.705 236.080 -33.535 236.250 ;
        RECT -32.415 236.080 -32.245 236.250 ;
        RECT -31.125 236.080 -30.955 236.250 ;
        RECT -29.835 236.080 -29.665 236.250 ;
        RECT -28.545 236.080 -28.375 236.250 ;
        RECT -27.255 236.080 -27.085 236.250 ;
        RECT 46.185 236.385 52.475 236.915 ;
        RECT 72.055 236.245 77.265 236.775 ;
        RECT 85.650 236.630 85.820 236.800 ;
        RECT 86.010 236.630 86.180 236.800 ;
        RECT 86.370 236.630 86.540 236.800 ;
        RECT 86.730 236.630 86.900 236.800 ;
        RECT 87.090 236.630 87.260 236.800 ;
        RECT 87.450 236.630 87.620 236.800 ;
        RECT 87.810 236.630 87.980 236.800 ;
        RECT 88.170 236.630 88.340 236.800 ;
        RECT 88.530 236.630 88.700 236.800 ;
        RECT 88.890 236.630 89.060 236.800 ;
        RECT 89.250 236.630 89.420 236.800 ;
        RECT 89.610 236.630 89.780 236.800 ;
        RECT 89.970 236.630 90.140 236.800 ;
        RECT 90.330 236.630 90.500 236.800 ;
        RECT 90.690 236.630 90.860 236.800 ;
        RECT 91.050 236.630 91.220 236.800 ;
        RECT 91.410 236.630 91.580 236.800 ;
        RECT 97.955 236.285 102.085 236.815 ;
        RECT -52.410 233.800 -52.240 233.970 ;
        RECT -52.410 233.440 -52.240 233.610 ;
        RECT -52.410 233.080 -52.240 233.250 ;
        RECT -52.410 232.720 -52.240 232.890 ;
        RECT -49.830 233.800 -49.660 233.970 ;
        RECT -49.830 233.440 -49.660 233.610 ;
        RECT -49.830 233.080 -49.660 233.250 ;
        RECT -49.830 232.720 -49.660 232.890 ;
        RECT -47.250 233.800 -47.080 233.970 ;
        RECT -47.250 233.440 -47.080 233.610 ;
        RECT -47.250 233.080 -47.080 233.250 ;
        RECT -47.250 232.720 -47.080 232.890 ;
        RECT -44.670 233.800 -44.500 233.970 ;
        RECT -44.670 233.440 -44.500 233.610 ;
        RECT -44.670 233.080 -44.500 233.250 ;
        RECT -44.670 232.720 -44.500 232.890 ;
        RECT -42.090 233.800 -41.920 233.970 ;
        RECT -42.090 233.440 -41.920 233.610 ;
        RECT -42.090 233.080 -41.920 233.250 ;
        RECT -42.090 232.720 -41.920 232.890 ;
        RECT -39.510 233.800 -39.340 233.970 ;
        RECT -39.510 233.440 -39.340 233.610 ;
        RECT -39.510 233.080 -39.340 233.250 ;
        RECT -39.510 232.720 -39.340 232.890 ;
        RECT -36.930 233.800 -36.760 233.970 ;
        RECT -36.930 233.440 -36.760 233.610 ;
        RECT -36.930 233.080 -36.760 233.250 ;
        RECT -36.930 232.720 -36.760 232.890 ;
        RECT -34.350 233.800 -34.180 233.970 ;
        RECT -34.350 233.440 -34.180 233.610 ;
        RECT -34.350 233.080 -34.180 233.250 ;
        RECT -34.350 232.720 -34.180 232.890 ;
        RECT -31.770 233.800 -31.600 233.970 ;
        RECT -31.770 233.440 -31.600 233.610 ;
        RECT -31.770 233.080 -31.600 233.250 ;
        RECT -31.770 232.720 -31.600 232.890 ;
        RECT -29.190 233.800 -29.020 233.970 ;
        RECT -29.190 233.440 -29.020 233.610 ;
        RECT -29.190 233.080 -29.020 233.250 ;
        RECT -29.190 232.720 -29.020 232.890 ;
        RECT -26.610 233.800 -26.440 233.970 ;
        RECT -26.610 233.440 -26.440 233.610 ;
        RECT -26.610 233.080 -26.440 233.250 ;
        RECT -26.610 232.720 -26.440 232.890 ;
        RECT -46.010 224.695 -32.520 227.025 ;
        RECT -51.655 223.930 -51.485 224.100 ;
        RECT -50.365 223.930 -50.195 224.100 ;
        RECT -49.075 223.930 -48.905 224.100 ;
        RECT -47.785 223.930 -47.615 224.100 ;
        RECT -46.495 223.930 -46.325 224.100 ;
        RECT -45.205 223.930 -45.035 224.100 ;
        RECT -43.915 223.930 -43.745 224.100 ;
        RECT -42.625 223.930 -42.455 224.100 ;
        RECT -41.335 223.930 -41.165 224.100 ;
        RECT -40.045 223.930 -39.875 224.100 ;
        RECT -38.755 223.930 -38.585 224.100 ;
        RECT -37.465 223.930 -37.295 224.100 ;
        RECT -36.175 223.930 -36.005 224.100 ;
        RECT -34.885 223.930 -34.715 224.100 ;
        RECT -33.595 223.930 -33.425 224.100 ;
        RECT -32.305 223.930 -32.135 224.100 ;
        RECT -31.015 223.930 -30.845 224.100 ;
        RECT -29.725 223.930 -29.555 224.100 ;
        RECT -28.435 223.930 -28.265 224.100 ;
        RECT -27.145 223.930 -26.975 224.100 ;
        RECT -52.300 221.650 -52.130 221.820 ;
        RECT -52.300 221.290 -52.130 221.460 ;
        RECT -52.300 220.930 -52.130 221.100 ;
        RECT -52.300 220.570 -52.130 220.740 ;
        RECT -49.720 221.650 -49.550 221.820 ;
        RECT -49.720 221.290 -49.550 221.460 ;
        RECT -49.720 220.930 -49.550 221.100 ;
        RECT -49.720 220.570 -49.550 220.740 ;
        RECT -47.140 221.650 -46.970 221.820 ;
        RECT -47.140 221.290 -46.970 221.460 ;
        RECT -47.140 220.930 -46.970 221.100 ;
        RECT -47.140 220.570 -46.970 220.740 ;
        RECT -44.560 221.650 -44.390 221.820 ;
        RECT -44.560 221.290 -44.390 221.460 ;
        RECT -44.560 220.930 -44.390 221.100 ;
        RECT -44.560 220.570 -44.390 220.740 ;
        RECT -41.980 221.650 -41.810 221.820 ;
        RECT -41.980 221.290 -41.810 221.460 ;
        RECT -41.980 220.930 -41.810 221.100 ;
        RECT -41.980 220.570 -41.810 220.740 ;
        RECT -39.400 221.650 -39.230 221.820 ;
        RECT -39.400 221.290 -39.230 221.460 ;
        RECT -39.400 220.930 -39.230 221.100 ;
        RECT -39.400 220.570 -39.230 220.740 ;
        RECT -36.820 221.650 -36.650 221.820 ;
        RECT -36.820 221.290 -36.650 221.460 ;
        RECT -36.820 220.930 -36.650 221.100 ;
        RECT -36.820 220.570 -36.650 220.740 ;
        RECT -34.240 221.650 -34.070 221.820 ;
        RECT -34.240 221.290 -34.070 221.460 ;
        RECT -34.240 220.930 -34.070 221.100 ;
        RECT -34.240 220.570 -34.070 220.740 ;
        RECT -31.660 221.650 -31.490 221.820 ;
        RECT -31.660 221.290 -31.490 221.460 ;
        RECT -31.660 220.930 -31.490 221.100 ;
        RECT -31.660 220.570 -31.490 220.740 ;
        RECT -29.080 221.650 -28.910 221.820 ;
        RECT -29.080 221.290 -28.910 221.460 ;
        RECT -29.080 220.930 -28.910 221.100 ;
        RECT -29.080 220.570 -28.910 220.740 ;
        RECT -26.500 221.650 -26.330 221.820 ;
        RECT -26.500 221.290 -26.330 221.460 ;
        RECT -26.500 220.930 -26.330 221.100 ;
        RECT -26.500 220.570 -26.330 220.740 ;
        RECT -46.010 137.085 -32.520 139.415 ;
        RECT -51.695 136.280 -51.525 136.450 ;
        RECT -50.405 136.280 -50.235 136.450 ;
        RECT -49.115 136.280 -48.945 136.450 ;
        RECT -47.825 136.280 -47.655 136.450 ;
        RECT -46.535 136.280 -46.365 136.450 ;
        RECT -45.245 136.280 -45.075 136.450 ;
        RECT -43.955 136.280 -43.785 136.450 ;
        RECT -42.665 136.280 -42.495 136.450 ;
        RECT -41.375 136.280 -41.205 136.450 ;
        RECT -40.085 136.280 -39.915 136.450 ;
        RECT -38.795 136.280 -38.625 136.450 ;
        RECT -37.505 136.280 -37.335 136.450 ;
        RECT -36.215 136.280 -36.045 136.450 ;
        RECT -34.925 136.280 -34.755 136.450 ;
        RECT -33.635 136.280 -33.465 136.450 ;
        RECT -32.345 136.280 -32.175 136.450 ;
        RECT -31.055 136.280 -30.885 136.450 ;
        RECT -29.765 136.280 -29.595 136.450 ;
        RECT -28.475 136.280 -28.305 136.450 ;
        RECT -27.185 136.280 -27.015 136.450 ;
        RECT -52.340 134.000 -52.170 134.170 ;
        RECT -52.340 133.640 -52.170 133.810 ;
        RECT -52.340 133.280 -52.170 133.450 ;
        RECT -52.340 132.920 -52.170 133.090 ;
        RECT -49.760 134.000 -49.590 134.170 ;
        RECT -49.760 133.640 -49.590 133.810 ;
        RECT -49.760 133.280 -49.590 133.450 ;
        RECT -49.760 132.920 -49.590 133.090 ;
        RECT -47.180 134.000 -47.010 134.170 ;
        RECT -47.180 133.640 -47.010 133.810 ;
        RECT -47.180 133.280 -47.010 133.450 ;
        RECT -47.180 132.920 -47.010 133.090 ;
        RECT -44.600 134.000 -44.430 134.170 ;
        RECT -44.600 133.640 -44.430 133.810 ;
        RECT -44.600 133.280 -44.430 133.450 ;
        RECT -44.600 132.920 -44.430 133.090 ;
        RECT -42.020 134.000 -41.850 134.170 ;
        RECT -42.020 133.640 -41.850 133.810 ;
        RECT -42.020 133.280 -41.850 133.450 ;
        RECT -42.020 132.920 -41.850 133.090 ;
        RECT -39.440 134.000 -39.270 134.170 ;
        RECT -39.440 133.640 -39.270 133.810 ;
        RECT -39.440 133.280 -39.270 133.450 ;
        RECT -39.440 132.920 -39.270 133.090 ;
        RECT -36.860 134.000 -36.690 134.170 ;
        RECT -36.860 133.640 -36.690 133.810 ;
        RECT -36.860 133.280 -36.690 133.450 ;
        RECT -36.860 132.920 -36.690 133.090 ;
        RECT -34.280 134.000 -34.110 134.170 ;
        RECT -34.280 133.640 -34.110 133.810 ;
        RECT -34.280 133.280 -34.110 133.450 ;
        RECT -34.280 132.920 -34.110 133.090 ;
        RECT -31.700 134.000 -31.530 134.170 ;
        RECT -31.700 133.640 -31.530 133.810 ;
        RECT -31.700 133.280 -31.530 133.450 ;
        RECT -31.700 132.920 -31.530 133.090 ;
        RECT -29.120 134.000 -28.950 134.170 ;
        RECT -29.120 133.640 -28.950 133.810 ;
        RECT -29.120 133.280 -28.950 133.450 ;
        RECT -29.120 132.920 -28.950 133.090 ;
        RECT -26.540 134.000 -26.370 134.170 ;
        RECT -26.540 133.640 -26.370 133.810 ;
        RECT -26.540 133.280 -26.370 133.450 ;
        RECT -26.540 132.920 -26.370 133.090 ;
        RECT -45.890 17.645 -32.400 19.975 ;
        RECT -51.575 16.840 -51.405 17.010 ;
        RECT -50.285 16.840 -50.115 17.010 ;
        RECT -48.995 16.840 -48.825 17.010 ;
        RECT -47.705 16.840 -47.535 17.010 ;
        RECT -46.415 16.840 -46.245 17.010 ;
        RECT -45.125 16.840 -44.955 17.010 ;
        RECT -43.835 16.840 -43.665 17.010 ;
        RECT -42.545 16.840 -42.375 17.010 ;
        RECT -41.255 16.840 -41.085 17.010 ;
        RECT -39.965 16.840 -39.795 17.010 ;
        RECT -38.675 16.840 -38.505 17.010 ;
        RECT -37.385 16.840 -37.215 17.010 ;
        RECT -36.095 16.840 -35.925 17.010 ;
        RECT -34.805 16.840 -34.635 17.010 ;
        RECT -33.515 16.840 -33.345 17.010 ;
        RECT -32.225 16.840 -32.055 17.010 ;
        RECT -30.935 16.840 -30.765 17.010 ;
        RECT -29.645 16.840 -29.475 17.010 ;
        RECT -28.355 16.840 -28.185 17.010 ;
        RECT -27.065 16.840 -26.895 17.010 ;
        RECT -52.220 14.560 -52.050 14.730 ;
        RECT -52.220 14.200 -52.050 14.370 ;
        RECT -52.220 13.840 -52.050 14.010 ;
        RECT -52.220 13.480 -52.050 13.650 ;
        RECT -49.640 14.560 -49.470 14.730 ;
        RECT -49.640 14.200 -49.470 14.370 ;
        RECT -49.640 13.840 -49.470 14.010 ;
        RECT -49.640 13.480 -49.470 13.650 ;
        RECT -47.060 14.560 -46.890 14.730 ;
        RECT -47.060 14.200 -46.890 14.370 ;
        RECT -47.060 13.840 -46.890 14.010 ;
        RECT -47.060 13.480 -46.890 13.650 ;
        RECT -44.480 14.560 -44.310 14.730 ;
        RECT -44.480 14.200 -44.310 14.370 ;
        RECT -44.480 13.840 -44.310 14.010 ;
        RECT -44.480 13.480 -44.310 13.650 ;
        RECT -41.900 14.560 -41.730 14.730 ;
        RECT -41.900 14.200 -41.730 14.370 ;
        RECT -41.900 13.840 -41.730 14.010 ;
        RECT -41.900 13.480 -41.730 13.650 ;
        RECT -39.320 14.560 -39.150 14.730 ;
        RECT -39.320 14.200 -39.150 14.370 ;
        RECT -39.320 13.840 -39.150 14.010 ;
        RECT -39.320 13.480 -39.150 13.650 ;
        RECT -36.740 14.560 -36.570 14.730 ;
        RECT -36.740 14.200 -36.570 14.370 ;
        RECT -36.740 13.840 -36.570 14.010 ;
        RECT -36.740 13.480 -36.570 13.650 ;
        RECT -34.160 14.560 -33.990 14.730 ;
        RECT -34.160 14.200 -33.990 14.370 ;
        RECT -34.160 13.840 -33.990 14.010 ;
        RECT -34.160 13.480 -33.990 13.650 ;
        RECT -31.580 14.560 -31.410 14.730 ;
        RECT -31.580 14.200 -31.410 14.370 ;
        RECT -31.580 13.840 -31.410 14.010 ;
        RECT -31.580 13.480 -31.410 13.650 ;
        RECT -29.000 14.560 -28.830 14.730 ;
        RECT -29.000 14.200 -28.830 14.370 ;
        RECT -29.000 13.840 -28.830 14.010 ;
        RECT -29.000 13.480 -28.830 13.650 ;
        RECT -26.420 14.560 -26.250 14.730 ;
        RECT -26.420 14.200 -26.250 14.370 ;
        RECT -26.420 13.840 -26.250 14.010 ;
        RECT -26.420 13.480 -26.250 13.650 ;
      LAYER met1 ;
        RECT -34.750 409.540 29.620 410.950 ;
        RECT -34.750 409.430 944.550 409.540 ;
        RECT 1072.580 409.430 1130.800 409.810 ;
        RECT -34.750 380.150 1130.800 409.430 ;
        RECT -34.750 379.880 1085.940 380.150 ;
        RECT -34.750 379.370 32.450 379.880 ;
        RECT -34.750 378.470 29.620 379.370 ;
        RECT 18.880 378.150 22.880 378.470 ;
        RECT -44.650 357.960 -34.300 359.660 ;
        RECT -51.960 357.430 -51.420 357.660 ;
        RECT -50.670 357.430 -50.130 357.660 ;
        RECT -49.380 357.430 -48.840 357.660 ;
        RECT -48.090 357.430 -47.550 357.660 ;
        RECT -46.800 357.430 -46.260 357.660 ;
        RECT -45.510 357.430 -44.970 357.660 ;
        RECT -44.220 357.430 -43.680 357.660 ;
        RECT -42.930 357.430 -42.390 357.660 ;
        RECT -41.640 357.430 -41.100 357.660 ;
        RECT -40.350 357.430 -39.810 357.660 ;
        RECT -39.060 357.430 -38.520 357.660 ;
        RECT -37.770 357.430 -37.230 357.660 ;
        RECT -36.480 357.430 -35.940 357.660 ;
        RECT -35.190 357.430 -34.650 357.660 ;
        RECT -33.900 357.430 -33.360 357.660 ;
        RECT -32.610 357.430 -32.070 357.660 ;
        RECT -31.320 357.430 -30.780 357.660 ;
        RECT -30.030 357.430 -29.490 357.660 ;
        RECT -28.740 357.430 -28.200 357.660 ;
        RECT -27.450 357.430 -26.910 357.660 ;
        RECT -52.485 356.770 -52.215 356.790 ;
        RECT -44.045 356.770 -43.895 357.430 ;
        RECT -52.555 356.430 -26.305 356.770 ;
        RECT -52.485 355.310 -52.215 356.430 ;
        RECT -49.845 355.515 -49.575 356.430 ;
        RECT -52.450 353.935 -52.220 355.310 ;
        RECT -49.870 355.270 -49.575 355.515 ;
        RECT -49.870 353.935 -49.640 355.270 ;
        RECT -47.315 355.250 -47.045 356.430 ;
        RECT -47.290 353.935 -47.060 355.250 ;
        RECT -44.725 355.190 -44.455 356.430 ;
        RECT -42.145 355.190 -41.875 356.430 ;
        RECT -44.710 353.935 -44.480 355.190 ;
        RECT -42.130 353.935 -41.900 355.190 ;
        RECT -39.575 355.130 -39.305 356.430 ;
        RECT -39.550 353.935 -39.320 355.130 ;
        RECT -36.985 355.110 -36.715 356.430 ;
        RECT -34.405 355.250 -34.135 356.430 ;
        RECT -36.970 353.935 -36.740 355.110 ;
        RECT -34.390 353.935 -34.160 355.250 ;
        RECT -31.835 355.230 -31.565 356.430 ;
        RECT -29.235 355.230 -28.965 356.430 ;
        RECT -26.645 355.515 -26.375 356.430 ;
        RECT -31.810 353.935 -31.580 355.230 ;
        RECT -29.230 353.935 -29.000 355.230 ;
        RECT -26.650 355.190 -26.375 355.515 ;
        RECT -26.650 353.935 -26.420 355.190 ;
        RECT 18.890 346.010 22.880 378.150 ;
        RECT 205.900 369.210 207.630 369.470 ;
        RECT 205.900 368.840 215.940 369.210 ;
        RECT 205.900 368.440 227.000 368.840 ;
        RECT 281.100 368.830 283.020 379.880 ;
        RECT 293.960 379.560 1085.940 379.880 ;
        RECT 233.810 368.440 247.040 368.830 ;
        RECT 253.870 368.440 267.100 368.830 ;
        RECT 273.920 368.440 287.150 368.830 ;
        RECT 205.900 367.520 287.150 368.440 ;
        RECT 205.900 366.930 227.000 367.520 ;
        RECT 18.890 343.020 23.000 346.010 ;
        RECT 4.860 329.790 13.020 329.810 ;
        RECT 19.390 329.790 23.000 343.020 ;
        RECT 31.570 329.790 39.730 329.820 ;
        RECT 44.800 329.790 52.960 329.820 ;
        RECT 71.340 329.790 79.500 329.820 ;
        RECT 84.470 329.790 92.630 329.840 ;
        RECT 96.960 329.790 103.140 329.970 ;
        RECT 4.860 329.650 103.140 329.790 ;
        RECT 1.310 329.620 103.140 329.650 ;
        RECT 1.170 328.950 103.140 329.620 ;
        RECT 1.170 328.790 13.020 328.950 ;
        RECT 1.170 328.480 9.310 328.790 ;
        RECT 18.200 328.770 26.360 328.950 ;
        RECT 31.570 328.800 39.730 328.950 ;
        RECT 44.800 328.800 52.960 328.950 ;
        RECT 58.070 328.770 66.230 328.950 ;
        RECT 71.340 328.800 79.500 328.950 ;
        RECT 84.470 328.820 92.630 328.950 ;
        RECT 96.960 328.620 103.140 328.950 ;
        RECT 1.170 298.870 2.470 328.480 ;
        RECT 4.770 327.650 5.750 327.880 ;
        RECT 8.240 327.650 9.220 327.880 ;
        RECT 11.710 327.650 12.690 327.880 ;
        RECT 18.110 327.630 19.090 327.860 ;
        RECT 21.580 327.630 22.560 327.860 ;
        RECT 25.050 327.630 26.030 327.860 ;
        RECT 31.480 327.660 32.460 327.890 ;
        RECT 34.950 327.660 35.930 327.890 ;
        RECT 38.420 327.660 39.400 327.890 ;
        RECT 44.710 327.660 45.690 327.890 ;
        RECT 48.180 327.660 49.160 327.890 ;
        RECT 51.650 327.660 52.630 327.890 ;
        RECT 57.980 327.630 58.960 327.860 ;
        RECT 61.450 327.630 62.430 327.860 ;
        RECT 64.920 327.630 65.900 327.860 ;
        RECT 71.250 327.660 72.230 327.890 ;
        RECT 74.720 327.660 75.700 327.890 ;
        RECT 78.190 327.660 79.170 327.890 ;
        RECT 84.380 327.680 85.360 327.910 ;
        RECT 87.850 327.680 88.830 327.910 ;
        RECT 91.320 327.680 92.300 327.910 ;
        RECT 97.800 327.900 98.780 328.130 ;
        RECT 101.270 327.900 102.250 328.130 ;
        RECT 205.900 325.040 207.630 366.930 ;
        RECT 213.770 366.830 227.000 366.930 ;
        RECT 233.810 366.820 247.040 367.520 ;
        RECT 253.870 366.820 267.100 367.520 ;
        RECT 273.920 366.820 287.150 367.520 ;
        RECT 211.990 365.940 212.970 366.170 ;
        RECT 215.460 365.940 216.440 366.170 ;
        RECT 218.930 365.940 219.910 366.170 ;
        RECT 222.400 365.940 223.380 366.170 ;
        RECT 225.870 365.940 226.850 366.170 ;
        RECT 282.680 366.160 283.610 366.820 ;
        RECT 232.030 365.930 233.010 366.160 ;
        RECT 235.500 365.930 236.480 366.160 ;
        RECT 238.970 365.930 239.950 366.160 ;
        RECT 242.440 365.930 243.420 366.160 ;
        RECT 245.910 365.930 246.890 366.160 ;
        RECT 252.090 365.930 253.070 366.160 ;
        RECT 255.560 365.930 256.540 366.160 ;
        RECT 259.030 365.930 260.010 366.160 ;
        RECT 262.500 365.930 263.480 366.160 ;
        RECT 265.970 365.930 266.950 366.160 ;
        RECT 272.140 365.930 273.120 366.160 ;
        RECT 275.610 365.930 276.590 366.160 ;
        RECT 279.080 365.930 280.060 366.160 ;
        RECT 282.550 366.010 283.610 366.160 ;
        RECT 282.550 365.930 283.530 366.010 ;
        RECT 286.020 365.930 287.000 366.160 ;
        RECT 354.920 363.890 356.240 379.560 ;
        RECT 362.820 371.640 364.540 372.690 ;
        RECT 356.660 369.280 356.890 370.260 ;
        RECT 359.950 369.280 360.180 370.260 ;
        RECT 363.240 369.280 363.470 370.260 ;
        RECT 366.530 369.620 366.760 370.260 ;
        RECT 366.200 367.660 366.830 369.620 ;
        RECT 369.820 369.280 370.050 370.260 ;
        RECT 366.190 367.500 366.830 367.660 ;
        RECT 366.190 367.330 366.690 367.500 ;
        RECT 356.520 364.710 356.750 365.690 ;
        RECT 359.810 364.710 360.040 365.690 ;
        RECT 363.100 364.710 363.330 365.690 ;
        RECT 366.200 365.360 366.690 367.330 ;
        RECT 366.330 365.350 366.690 365.360 ;
        RECT 366.390 364.710 366.620 365.350 ;
        RECT 369.680 364.710 369.910 365.690 ;
        RECT 374.370 365.530 374.950 379.560 ;
        RECT 375.980 369.180 376.210 370.160 ;
        RECT 382.560 369.180 382.790 370.160 ;
        RECT 388.850 369.720 389.650 379.560 ;
        RECT 389.140 369.180 389.370 369.720 ;
        RECT 393.730 365.600 394.310 379.560 ;
        RECT 401.570 371.830 404.570 373.040 ;
        RECT 395.230 369.250 395.460 370.230 ;
        RECT 398.520 369.250 398.750 370.230 ;
        RECT 401.810 369.250 402.040 370.230 ;
        RECT 405.100 369.590 405.330 370.230 ;
        RECT 404.770 367.630 405.400 369.590 ;
        RECT 408.390 369.250 408.620 370.230 ;
        RECT 404.760 367.470 405.400 367.630 ;
        RECT 404.760 367.300 405.260 367.470 ;
        RECT 211.990 362.650 212.970 362.880 ;
        RECT 215.460 362.650 216.440 362.880 ;
        RECT 218.930 362.650 219.910 362.880 ;
        RECT 222.400 362.650 223.380 362.880 ;
        RECT 225.870 362.650 226.850 362.880 ;
        RECT 232.030 362.640 233.010 362.870 ;
        RECT 235.500 362.640 236.480 362.870 ;
        RECT 238.970 362.640 239.950 362.870 ;
        RECT 242.440 362.640 243.420 362.870 ;
        RECT 245.910 362.640 246.890 362.870 ;
        RECT 252.090 362.640 253.070 362.870 ;
        RECT 255.560 362.640 256.540 362.870 ;
        RECT 259.030 362.640 260.010 362.870 ;
        RECT 262.500 362.640 263.480 362.870 ;
        RECT 265.970 362.640 266.950 362.870 ;
        RECT 272.140 362.640 273.120 362.870 ;
        RECT 275.610 362.640 276.590 362.870 ;
        RECT 279.080 362.640 280.060 362.870 ;
        RECT 282.550 362.640 283.530 362.870 ;
        RECT 286.020 362.640 287.000 362.870 ;
        RECT 211.990 359.360 212.970 359.590 ;
        RECT 215.460 359.360 216.440 359.590 ;
        RECT 218.930 359.360 219.910 359.590 ;
        RECT 222.400 359.360 223.380 359.590 ;
        RECT 225.870 359.360 226.850 359.590 ;
        RECT 232.030 359.350 233.010 359.580 ;
        RECT 235.500 359.350 236.480 359.580 ;
        RECT 238.970 359.350 239.950 359.580 ;
        RECT 242.440 359.350 243.420 359.580 ;
        RECT 245.910 359.350 246.890 359.580 ;
        RECT 252.090 359.350 253.070 359.580 ;
        RECT 255.560 359.350 256.540 359.580 ;
        RECT 259.030 359.350 260.010 359.580 ;
        RECT 262.500 359.350 263.480 359.580 ;
        RECT 265.970 359.350 266.950 359.580 ;
        RECT 272.140 359.350 273.120 359.580 ;
        RECT 275.610 359.350 276.590 359.580 ;
        RECT 279.080 359.350 280.060 359.580 ;
        RECT 282.550 359.350 283.530 359.580 ;
        RECT 286.020 359.350 287.000 359.580 ;
        RECT 211.990 356.070 212.970 356.300 ;
        RECT 215.460 356.070 216.440 356.300 ;
        RECT 218.930 356.070 219.910 356.300 ;
        RECT 222.400 356.070 223.380 356.300 ;
        RECT 225.870 356.070 226.850 356.300 ;
        RECT 232.030 356.060 233.010 356.290 ;
        RECT 235.500 356.060 236.480 356.290 ;
        RECT 238.970 356.060 239.950 356.290 ;
        RECT 242.440 356.060 243.420 356.290 ;
        RECT 245.910 356.060 246.890 356.290 ;
        RECT 252.090 356.060 253.070 356.290 ;
        RECT 255.560 356.060 256.540 356.290 ;
        RECT 259.030 356.060 260.010 356.290 ;
        RECT 262.500 356.060 263.480 356.290 ;
        RECT 265.970 356.060 266.950 356.290 ;
        RECT 272.140 356.060 273.120 356.290 ;
        RECT 275.610 356.060 276.590 356.290 ;
        RECT 279.080 356.060 280.060 356.290 ;
        RECT 282.550 356.060 283.530 356.290 ;
        RECT 286.020 356.060 287.000 356.290 ;
        RECT 211.990 352.780 212.970 353.010 ;
        RECT 215.460 352.780 216.440 353.010 ;
        RECT 218.930 352.780 219.910 353.010 ;
        RECT 222.400 352.780 223.380 353.010 ;
        RECT 225.870 352.780 226.850 353.010 ;
        RECT 232.030 352.770 233.010 353.000 ;
        RECT 235.500 352.770 236.480 353.000 ;
        RECT 238.970 352.770 239.950 353.000 ;
        RECT 242.440 352.770 243.420 353.000 ;
        RECT 245.910 352.770 246.890 353.000 ;
        RECT 252.090 352.770 253.070 353.000 ;
        RECT 255.560 352.770 256.540 353.000 ;
        RECT 259.030 352.770 260.010 353.000 ;
        RECT 262.500 352.770 263.480 353.000 ;
        RECT 265.970 352.770 266.950 353.000 ;
        RECT 272.140 352.770 273.120 353.000 ;
        RECT 275.610 352.770 276.590 353.000 ;
        RECT 279.080 352.770 280.060 353.000 ;
        RECT 282.550 352.770 283.530 353.000 ;
        RECT 286.020 352.770 287.000 353.000 ;
        RECT 355.060 351.330 356.140 363.890 ;
        RECT 356.520 361.240 356.750 362.220 ;
        RECT 359.810 361.240 360.040 362.220 ;
        RECT 363.100 361.240 363.330 362.220 ;
        RECT 366.390 361.240 366.620 362.220 ;
        RECT 369.680 361.240 369.910 362.220 ;
        RECT 356.520 357.770 356.750 358.750 ;
        RECT 359.810 357.770 360.040 358.750 ;
        RECT 363.100 357.770 363.330 358.750 ;
        RECT 366.390 357.770 366.620 358.750 ;
        RECT 369.680 357.770 369.910 358.750 ;
        RECT 356.520 354.300 356.750 355.280 ;
        RECT 359.810 354.300 360.040 355.280 ;
        RECT 363.100 354.300 363.330 355.280 ;
        RECT 366.390 354.300 366.620 355.280 ;
        RECT 369.680 354.300 369.910 355.280 ;
        RECT 356.520 350.830 356.750 351.810 ;
        RECT 359.810 350.830 360.040 351.810 ;
        RECT 363.100 350.830 363.330 351.810 ;
        RECT 366.390 351.180 366.620 351.810 ;
        RECT 211.990 349.490 212.970 349.720 ;
        RECT 215.460 349.490 216.440 349.720 ;
        RECT 218.930 349.490 219.910 349.720 ;
        RECT 222.400 349.490 223.380 349.720 ;
        RECT 225.870 349.490 226.850 349.720 ;
        RECT 232.030 349.480 233.010 349.710 ;
        RECT 235.500 349.480 236.480 349.710 ;
        RECT 238.970 349.480 239.950 349.710 ;
        RECT 242.440 349.480 243.420 349.710 ;
        RECT 245.910 349.480 246.890 349.710 ;
        RECT 252.090 349.480 253.070 349.710 ;
        RECT 255.560 349.480 256.540 349.710 ;
        RECT 259.030 349.480 260.010 349.710 ;
        RECT 262.500 349.480 263.480 349.710 ;
        RECT 265.970 349.480 266.950 349.710 ;
        RECT 272.140 349.480 273.120 349.710 ;
        RECT 275.610 349.480 276.590 349.710 ;
        RECT 279.080 349.480 280.060 349.710 ;
        RECT 282.550 349.480 283.530 349.710 ;
        RECT 286.020 349.480 287.000 349.710 ;
        RECT 213.730 347.280 226.960 347.850 ;
        RECT 233.700 347.280 246.930 347.850 ;
        RECT 253.810 347.280 267.040 347.850 ;
        RECT 273.920 347.280 287.150 347.850 ;
        RECT 213.730 346.360 287.150 347.280 ;
        RECT 288.460 347.040 289.350 348.760 ;
        RECT 213.730 345.840 226.960 346.360 ;
        RECT 233.700 345.840 246.930 346.360 ;
        RECT 253.810 345.840 267.040 346.360 ;
        RECT 273.920 345.840 287.150 346.360 ;
        RECT 285.930 345.180 286.860 345.840 ;
        RECT 211.950 344.950 212.930 345.180 ;
        RECT 215.420 344.950 216.400 345.180 ;
        RECT 218.890 344.950 219.870 345.180 ;
        RECT 222.360 344.950 223.340 345.180 ;
        RECT 225.830 344.950 226.810 345.180 ;
        RECT 231.920 344.950 232.900 345.180 ;
        RECT 235.390 344.950 236.370 345.180 ;
        RECT 238.860 344.950 239.840 345.180 ;
        RECT 242.330 344.950 243.310 345.180 ;
        RECT 245.800 344.950 246.780 345.180 ;
        RECT 252.030 344.950 253.010 345.180 ;
        RECT 255.500 344.950 256.480 345.180 ;
        RECT 258.970 344.950 259.950 345.180 ;
        RECT 262.440 344.950 263.420 345.180 ;
        RECT 265.910 344.950 266.890 345.180 ;
        RECT 272.140 344.950 273.120 345.180 ;
        RECT 275.610 344.950 276.590 345.180 ;
        RECT 279.080 344.950 280.060 345.180 ;
        RECT 282.550 344.950 283.530 345.180 ;
        RECT 285.930 344.970 287.000 345.180 ;
        RECT 286.020 344.950 287.000 344.970 ;
        RECT 211.950 341.660 212.930 341.890 ;
        RECT 215.420 341.660 216.400 341.890 ;
        RECT 218.890 341.660 219.870 341.890 ;
        RECT 222.360 341.660 223.340 341.890 ;
        RECT 225.830 341.660 226.810 341.890 ;
        RECT 231.920 341.660 232.900 341.890 ;
        RECT 235.390 341.660 236.370 341.890 ;
        RECT 238.860 341.660 239.840 341.890 ;
        RECT 242.330 341.660 243.310 341.890 ;
        RECT 245.800 341.660 246.780 341.890 ;
        RECT 252.030 341.660 253.010 341.890 ;
        RECT 255.500 341.660 256.480 341.890 ;
        RECT 258.970 341.660 259.950 341.890 ;
        RECT 262.440 341.660 263.420 341.890 ;
        RECT 265.910 341.660 266.890 341.890 ;
        RECT 272.140 341.660 273.120 341.890 ;
        RECT 275.610 341.660 276.590 341.890 ;
        RECT 279.080 341.660 280.060 341.890 ;
        RECT 282.550 341.660 283.530 341.890 ;
        RECT 286.020 341.660 287.000 341.890 ;
        RECT 211.950 338.370 212.930 338.600 ;
        RECT 215.420 338.370 216.400 338.600 ;
        RECT 218.890 338.370 219.870 338.600 ;
        RECT 222.360 338.370 223.340 338.600 ;
        RECT 225.830 338.370 226.810 338.600 ;
        RECT 231.920 338.370 232.900 338.600 ;
        RECT 235.390 338.370 236.370 338.600 ;
        RECT 238.860 338.370 239.840 338.600 ;
        RECT 242.330 338.370 243.310 338.600 ;
        RECT 245.800 338.370 246.780 338.600 ;
        RECT 252.030 338.370 253.010 338.600 ;
        RECT 255.500 338.370 256.480 338.600 ;
        RECT 258.970 338.370 259.950 338.600 ;
        RECT 262.440 338.370 263.420 338.600 ;
        RECT 265.910 338.370 266.890 338.600 ;
        RECT 272.140 338.370 273.120 338.600 ;
        RECT 275.610 338.370 276.590 338.600 ;
        RECT 279.080 338.370 280.060 338.600 ;
        RECT 282.550 338.370 283.530 338.600 ;
        RECT 286.020 338.370 287.000 338.600 ;
        RECT 211.950 335.080 212.930 335.310 ;
        RECT 215.420 335.080 216.400 335.310 ;
        RECT 218.890 335.080 219.870 335.310 ;
        RECT 222.360 335.080 223.340 335.310 ;
        RECT 225.830 335.080 226.810 335.310 ;
        RECT 231.920 335.080 232.900 335.310 ;
        RECT 235.390 335.080 236.370 335.310 ;
        RECT 238.860 335.080 239.840 335.310 ;
        RECT 242.330 335.080 243.310 335.310 ;
        RECT 245.800 335.080 246.780 335.310 ;
        RECT 252.030 335.080 253.010 335.310 ;
        RECT 255.500 335.080 256.480 335.310 ;
        RECT 258.970 335.080 259.950 335.310 ;
        RECT 262.440 335.080 263.420 335.310 ;
        RECT 265.910 335.080 266.890 335.310 ;
        RECT 272.140 335.080 273.120 335.310 ;
        RECT 275.610 335.080 276.590 335.310 ;
        RECT 279.080 335.080 280.060 335.310 ;
        RECT 282.550 335.080 283.530 335.310 ;
        RECT 286.020 335.080 287.000 335.310 ;
        RECT 355.040 332.450 356.120 346.750 ;
        RECT 356.500 345.830 356.730 346.810 ;
        RECT 359.790 345.830 360.020 346.810 ;
        RECT 363.080 345.830 363.310 346.810 ;
        RECT 366.310 346.450 366.730 351.180 ;
        RECT 369.680 350.830 369.910 351.810 ;
        RECT 374.370 351.230 375.460 365.530 ;
        RECT 375.840 364.610 376.070 365.590 ;
        RECT 382.420 364.610 382.650 365.590 ;
        RECT 389.000 364.610 389.230 365.590 ;
        RECT 375.840 361.140 376.070 362.120 ;
        RECT 382.420 361.140 382.650 362.120 ;
        RECT 389.000 361.140 389.230 362.120 ;
        RECT 375.840 357.670 376.070 358.650 ;
        RECT 382.420 357.670 382.650 358.650 ;
        RECT 389.000 357.670 389.230 358.650 ;
        RECT 375.840 354.200 376.070 355.180 ;
        RECT 382.420 354.200 382.650 355.180 ;
        RECT 389.000 354.200 389.230 355.180 ;
        RECT 366.370 345.830 366.600 346.450 ;
        RECT 369.660 345.830 369.890 346.810 ;
        RECT 374.370 346.650 374.950 351.230 ;
        RECT 375.840 350.730 376.070 351.710 ;
        RECT 382.420 350.730 382.650 351.710 ;
        RECT 389.000 350.730 389.230 351.710 ;
        RECT 393.630 351.300 394.710 365.600 ;
        RECT 395.090 364.680 395.320 365.660 ;
        RECT 398.380 364.680 398.610 365.660 ;
        RECT 401.670 364.680 401.900 365.660 ;
        RECT 404.770 365.330 405.260 367.300 ;
        RECT 404.900 365.320 405.260 365.330 ;
        RECT 404.960 364.680 405.190 365.320 ;
        RECT 408.250 364.680 408.480 365.660 ;
        RECT 395.090 361.210 395.320 362.190 ;
        RECT 398.380 361.210 398.610 362.190 ;
        RECT 401.670 361.210 401.900 362.190 ;
        RECT 404.960 361.210 405.190 362.190 ;
        RECT 408.250 361.210 408.480 362.190 ;
        RECT 395.090 357.740 395.320 358.720 ;
        RECT 398.380 357.740 398.610 358.720 ;
        RECT 401.670 357.740 401.900 358.720 ;
        RECT 404.960 357.740 405.190 358.720 ;
        RECT 408.250 357.740 408.480 358.720 ;
        RECT 395.090 354.270 395.320 355.250 ;
        RECT 398.380 354.270 398.610 355.250 ;
        RECT 401.670 354.270 401.900 355.250 ;
        RECT 404.960 354.270 405.190 355.250 ;
        RECT 408.250 354.270 408.480 355.250 ;
        RECT 393.730 346.720 394.310 351.300 ;
        RECT 395.090 350.800 395.320 351.780 ;
        RECT 398.380 350.800 398.610 351.780 ;
        RECT 401.670 350.800 401.900 351.780 ;
        RECT 404.960 351.150 405.190 351.780 ;
        RECT 356.500 342.360 356.730 343.340 ;
        RECT 359.790 342.360 360.020 343.340 ;
        RECT 363.080 342.360 363.310 343.340 ;
        RECT 366.370 342.360 366.600 343.340 ;
        RECT 369.660 342.360 369.890 343.340 ;
        RECT 356.500 338.890 356.730 339.870 ;
        RECT 359.790 338.890 360.020 339.870 ;
        RECT 363.080 338.890 363.310 339.870 ;
        RECT 366.370 338.890 366.600 339.870 ;
        RECT 369.660 338.890 369.890 339.870 ;
        RECT 356.500 335.420 356.730 336.400 ;
        RECT 359.790 335.420 360.020 336.400 ;
        RECT 363.080 335.420 363.310 336.400 ;
        RECT 366.370 335.420 366.600 336.400 ;
        RECT 369.660 335.420 369.890 336.400 ;
        RECT 211.950 331.790 212.930 332.020 ;
        RECT 215.420 331.790 216.400 332.020 ;
        RECT 218.890 331.790 219.870 332.020 ;
        RECT 222.360 331.790 223.340 332.020 ;
        RECT 225.830 331.790 226.810 332.020 ;
        RECT 231.920 331.790 232.900 332.020 ;
        RECT 235.390 331.790 236.370 332.020 ;
        RECT 238.860 331.790 239.840 332.020 ;
        RECT 242.330 331.790 243.310 332.020 ;
        RECT 245.800 331.790 246.780 332.020 ;
        RECT 252.030 331.790 253.010 332.020 ;
        RECT 255.500 331.790 256.480 332.020 ;
        RECT 258.970 331.790 259.950 332.020 ;
        RECT 262.440 331.790 263.420 332.020 ;
        RECT 265.910 331.790 266.890 332.020 ;
        RECT 272.140 331.790 273.120 332.020 ;
        RECT 275.610 331.790 276.590 332.020 ;
        RECT 279.080 331.790 280.060 332.020 ;
        RECT 282.550 331.790 283.530 332.020 ;
        RECT 286.020 331.790 287.000 332.020 ;
        RECT 356.500 331.950 356.730 332.930 ;
        RECT 359.790 331.950 360.020 332.930 ;
        RECT 363.080 331.950 363.310 332.930 ;
        RECT 366.370 332.380 366.600 332.930 ;
        RECT 211.950 328.500 212.930 328.730 ;
        RECT 215.420 328.500 216.400 328.730 ;
        RECT 218.890 328.500 219.870 328.730 ;
        RECT 222.360 328.500 223.340 328.730 ;
        RECT 225.830 328.500 226.810 328.730 ;
        RECT 231.920 328.500 232.900 328.730 ;
        RECT 235.390 328.500 236.370 328.730 ;
        RECT 238.860 328.500 239.840 328.730 ;
        RECT 242.330 328.500 243.310 328.730 ;
        RECT 245.800 328.500 246.780 328.730 ;
        RECT 252.030 328.500 253.010 328.730 ;
        RECT 255.500 328.500 256.480 328.730 ;
        RECT 258.970 328.500 259.950 328.730 ;
        RECT 262.440 328.500 263.420 328.730 ;
        RECT 265.910 328.500 266.890 328.730 ;
        RECT 272.140 328.500 273.120 328.730 ;
        RECT 275.610 328.500 276.590 328.730 ;
        RECT 279.080 328.500 280.060 328.730 ;
        RECT 282.550 328.500 283.530 328.730 ;
        RECT 286.020 328.500 287.000 328.730 ;
        RECT 213.670 325.040 226.900 325.480 ;
        RECT 4.770 324.360 5.750 324.590 ;
        RECT 8.240 324.360 9.220 324.590 ;
        RECT 11.710 324.360 12.690 324.590 ;
        RECT 18.110 324.340 19.090 324.570 ;
        RECT 21.580 324.340 22.560 324.570 ;
        RECT 25.050 324.340 26.030 324.570 ;
        RECT 31.480 324.370 32.460 324.600 ;
        RECT 34.950 324.370 35.930 324.600 ;
        RECT 38.420 324.370 39.400 324.600 ;
        RECT 44.710 324.370 45.690 324.600 ;
        RECT 48.180 324.370 49.160 324.600 ;
        RECT 51.650 324.370 52.630 324.600 ;
        RECT 57.980 324.340 58.960 324.570 ;
        RECT 61.450 324.340 62.430 324.570 ;
        RECT 64.920 324.340 65.900 324.570 ;
        RECT 71.250 324.370 72.230 324.600 ;
        RECT 74.720 324.370 75.700 324.600 ;
        RECT 78.190 324.370 79.170 324.600 ;
        RECT 84.380 324.390 85.360 324.620 ;
        RECT 87.850 324.390 88.830 324.620 ;
        RECT 91.320 324.390 92.300 324.620 ;
        RECT 97.800 324.610 98.780 324.840 ;
        RECT 101.270 324.610 102.250 324.840 ;
        RECT 205.900 324.740 226.900 325.040 ;
        RECT 233.710 324.740 246.940 325.470 ;
        RECT 253.770 324.740 267.000 325.470 ;
        RECT 273.820 324.740 287.050 325.470 ;
        RECT 205.900 323.820 287.050 324.740 ;
        RECT 205.900 323.570 226.900 323.820 ;
        RECT 213.670 323.470 226.900 323.570 ;
        RECT 233.710 323.460 246.940 323.820 ;
        RECT 253.770 323.460 267.000 323.820 ;
        RECT 273.820 323.460 287.050 323.820 ;
        RECT 211.890 322.580 212.870 322.810 ;
        RECT 215.360 322.580 216.340 322.810 ;
        RECT 218.830 322.580 219.810 322.810 ;
        RECT 222.300 322.580 223.280 322.810 ;
        RECT 225.770 322.580 226.750 322.810 ;
        RECT 231.930 322.570 232.910 322.800 ;
        RECT 235.400 322.570 236.380 322.800 ;
        RECT 238.870 322.570 239.850 322.800 ;
        RECT 242.340 322.570 243.320 322.800 ;
        RECT 245.810 322.570 246.790 322.800 ;
        RECT 251.990 322.570 252.970 322.800 ;
        RECT 255.460 322.570 256.440 322.800 ;
        RECT 258.930 322.570 259.910 322.800 ;
        RECT 262.400 322.570 263.380 322.800 ;
        RECT 265.870 322.570 266.850 322.800 ;
        RECT 272.040 322.570 273.020 322.800 ;
        RECT 275.510 322.570 276.490 322.800 ;
        RECT 278.980 322.570 279.960 322.800 ;
        RECT 282.450 322.570 283.430 322.800 ;
        RECT 285.920 322.570 286.900 322.800 ;
        RECT 4.770 321.070 5.750 321.300 ;
        RECT 8.240 321.070 9.220 321.300 ;
        RECT 11.710 321.070 12.690 321.300 ;
        RECT 18.110 321.050 19.090 321.280 ;
        RECT 21.580 321.050 22.560 321.280 ;
        RECT 25.050 321.050 26.030 321.280 ;
        RECT 31.480 321.080 32.460 321.310 ;
        RECT 34.950 321.080 35.930 321.310 ;
        RECT 38.420 321.080 39.400 321.310 ;
        RECT 44.710 321.080 45.690 321.310 ;
        RECT 48.180 321.080 49.160 321.310 ;
        RECT 51.650 321.080 52.630 321.310 ;
        RECT 57.980 321.050 58.960 321.280 ;
        RECT 61.450 321.050 62.430 321.280 ;
        RECT 64.920 321.050 65.900 321.280 ;
        RECT 71.250 321.080 72.230 321.310 ;
        RECT 74.720 321.080 75.700 321.310 ;
        RECT 78.190 321.080 79.170 321.310 ;
        RECT 84.380 321.100 85.360 321.330 ;
        RECT 87.850 321.100 88.830 321.330 ;
        RECT 91.320 321.100 92.300 321.330 ;
        RECT 97.800 321.320 98.780 321.550 ;
        RECT 101.270 321.320 102.250 321.550 ;
        RECT 103.460 320.160 104.050 320.720 ;
        RECT 4.770 317.780 5.750 318.010 ;
        RECT 8.240 317.780 9.220 318.010 ;
        RECT 11.710 317.780 12.690 318.010 ;
        RECT 18.110 317.760 19.090 317.990 ;
        RECT 21.580 317.760 22.560 317.990 ;
        RECT 25.050 317.760 26.030 317.990 ;
        RECT 31.480 317.790 32.460 318.020 ;
        RECT 34.950 317.790 35.930 318.020 ;
        RECT 38.420 317.790 39.400 318.020 ;
        RECT 44.710 317.790 45.690 318.020 ;
        RECT 48.180 317.790 49.160 318.020 ;
        RECT 51.650 317.790 52.630 318.020 ;
        RECT 57.980 317.760 58.960 317.990 ;
        RECT 61.450 317.760 62.430 317.990 ;
        RECT 64.920 317.760 65.900 317.990 ;
        RECT 71.250 317.790 72.230 318.020 ;
        RECT 74.720 317.790 75.700 318.020 ;
        RECT 78.190 317.790 79.170 318.020 ;
        RECT 84.380 317.810 85.360 318.040 ;
        RECT 87.850 317.810 88.830 318.040 ;
        RECT 91.320 317.810 92.300 318.040 ;
        RECT 97.800 318.030 98.780 318.260 ;
        RECT 101.270 318.030 102.250 318.260 ;
        RECT 211.890 316.000 212.870 316.230 ;
        RECT 215.360 316.000 216.340 316.230 ;
        RECT 218.830 316.000 219.810 316.230 ;
        RECT 222.300 316.000 223.280 316.230 ;
        RECT 225.770 316.000 226.750 316.230 ;
        RECT 231.930 315.990 232.910 316.220 ;
        RECT 235.400 315.990 236.380 316.220 ;
        RECT 238.870 315.990 239.850 316.220 ;
        RECT 242.340 315.990 243.320 316.220 ;
        RECT 245.810 315.990 246.790 316.220 ;
        RECT 251.990 315.990 252.970 316.220 ;
        RECT 255.460 315.990 256.440 316.220 ;
        RECT 258.930 315.990 259.910 316.220 ;
        RECT 262.400 315.990 263.380 316.220 ;
        RECT 265.870 315.990 266.850 316.220 ;
        RECT 272.040 315.990 273.020 316.220 ;
        RECT 275.510 315.990 276.490 316.220 ;
        RECT 278.980 315.990 279.960 316.220 ;
        RECT 282.450 315.990 283.430 316.220 ;
        RECT 285.920 315.990 286.900 316.220 ;
        RECT 4.770 314.490 5.750 314.720 ;
        RECT 8.240 314.490 9.220 314.720 ;
        RECT 11.710 314.490 12.690 314.720 ;
        RECT 18.110 314.470 19.090 314.700 ;
        RECT 21.580 314.470 22.560 314.700 ;
        RECT 25.050 314.470 26.030 314.700 ;
        RECT 31.480 314.500 32.460 314.730 ;
        RECT 34.950 314.500 35.930 314.730 ;
        RECT 38.420 314.500 39.400 314.730 ;
        RECT 44.710 314.500 45.690 314.730 ;
        RECT 48.180 314.500 49.160 314.730 ;
        RECT 51.650 314.500 52.630 314.730 ;
        RECT 57.980 314.470 58.960 314.700 ;
        RECT 61.450 314.470 62.430 314.700 ;
        RECT 64.920 314.470 65.900 314.700 ;
        RECT 71.250 314.500 72.230 314.730 ;
        RECT 74.720 314.500 75.700 314.730 ;
        RECT 78.190 314.500 79.170 314.730 ;
        RECT 84.380 314.520 85.360 314.750 ;
        RECT 87.850 314.520 88.830 314.750 ;
        RECT 91.320 314.520 92.300 314.750 ;
        RECT 97.800 314.740 98.780 314.970 ;
        RECT 101.270 314.740 102.250 314.970 ;
        RECT 355.040 313.600 356.120 327.900 ;
        RECT 356.500 326.980 356.730 327.960 ;
        RECT 359.790 326.980 360.020 327.960 ;
        RECT 363.080 326.980 363.310 327.960 ;
        RECT 366.190 327.390 366.810 332.380 ;
        RECT 369.660 331.950 369.890 332.930 ;
        RECT 374.360 332.350 375.440 346.650 ;
        RECT 375.820 345.730 376.050 346.710 ;
        RECT 382.400 345.730 382.630 346.710 ;
        RECT 388.980 345.730 389.210 346.710 ;
        RECT 375.820 342.260 376.050 343.240 ;
        RECT 382.400 342.260 382.630 343.240 ;
        RECT 388.980 342.260 389.210 343.240 ;
        RECT 375.820 338.790 376.050 339.770 ;
        RECT 382.400 338.790 382.630 339.770 ;
        RECT 388.980 338.790 389.210 339.770 ;
        RECT 375.820 335.320 376.050 336.300 ;
        RECT 382.400 335.320 382.630 336.300 ;
        RECT 388.980 335.320 389.210 336.300 ;
        RECT 366.370 326.980 366.600 327.390 ;
        RECT 369.660 326.980 369.890 327.960 ;
        RECT 374.370 327.800 374.950 332.350 ;
        RECT 375.820 331.850 376.050 332.830 ;
        RECT 382.400 331.850 382.630 332.830 ;
        RECT 388.980 331.850 389.210 332.830 ;
        RECT 393.610 332.420 394.690 346.720 ;
        RECT 395.070 345.800 395.300 346.780 ;
        RECT 398.360 345.800 398.590 346.780 ;
        RECT 401.650 345.800 401.880 346.780 ;
        RECT 404.880 346.420 405.300 351.150 ;
        RECT 408.250 350.800 408.480 351.780 ;
        RECT 404.940 345.800 405.170 346.420 ;
        RECT 408.230 345.800 408.460 346.780 ;
        RECT 395.070 342.330 395.300 343.310 ;
        RECT 398.360 342.330 398.590 343.310 ;
        RECT 401.650 342.330 401.880 343.310 ;
        RECT 404.940 342.330 405.170 343.310 ;
        RECT 408.230 342.330 408.460 343.310 ;
        RECT 395.070 338.860 395.300 339.840 ;
        RECT 398.360 338.860 398.590 339.840 ;
        RECT 401.650 338.860 401.880 339.840 ;
        RECT 404.940 338.860 405.170 339.840 ;
        RECT 408.230 338.860 408.460 339.840 ;
        RECT 395.070 335.390 395.300 336.370 ;
        RECT 398.360 335.390 398.590 336.370 ;
        RECT 401.650 335.390 401.880 336.370 ;
        RECT 404.940 335.390 405.170 336.370 ;
        RECT 408.230 335.390 408.460 336.370 ;
        RECT 393.730 327.870 394.310 332.420 ;
        RECT 395.070 331.920 395.300 332.900 ;
        RECT 398.360 331.920 398.590 332.900 ;
        RECT 401.650 331.920 401.880 332.900 ;
        RECT 404.940 332.350 405.170 332.900 ;
        RECT 356.500 323.510 356.730 324.490 ;
        RECT 359.790 323.510 360.020 324.490 ;
        RECT 363.080 323.510 363.310 324.490 ;
        RECT 366.370 323.510 366.600 324.490 ;
        RECT 369.660 323.510 369.890 324.490 ;
        RECT 356.500 320.040 356.730 321.020 ;
        RECT 359.790 320.040 360.020 321.020 ;
        RECT 363.080 320.040 363.310 321.020 ;
        RECT 366.370 320.040 366.600 321.020 ;
        RECT 369.660 320.040 369.890 321.020 ;
        RECT 356.500 316.570 356.730 317.550 ;
        RECT 359.790 316.570 360.020 317.550 ;
        RECT 363.080 316.570 363.310 317.550 ;
        RECT 366.370 316.570 366.600 317.550 ;
        RECT 369.660 316.570 369.890 317.550 ;
        RECT 356.500 313.100 356.730 314.080 ;
        RECT 359.790 313.100 360.020 314.080 ;
        RECT 363.080 313.100 363.310 314.080 ;
        RECT 366.370 313.880 366.600 314.080 ;
        RECT 4.770 311.200 5.750 311.430 ;
        RECT 8.240 311.200 9.220 311.430 ;
        RECT 11.710 311.200 12.690 311.430 ;
        RECT 18.110 311.180 19.090 311.410 ;
        RECT 21.580 311.180 22.560 311.410 ;
        RECT 25.050 311.180 26.030 311.410 ;
        RECT 31.480 311.210 32.460 311.440 ;
        RECT 34.950 311.210 35.930 311.440 ;
        RECT 38.420 311.210 39.400 311.440 ;
        RECT 44.710 311.210 45.690 311.440 ;
        RECT 48.180 311.210 49.160 311.440 ;
        RECT 51.650 311.210 52.630 311.440 ;
        RECT 57.980 311.180 58.960 311.410 ;
        RECT 61.450 311.180 62.430 311.410 ;
        RECT 64.920 311.180 65.900 311.410 ;
        RECT 71.250 311.210 72.230 311.440 ;
        RECT 74.720 311.210 75.700 311.440 ;
        RECT 78.190 311.210 79.170 311.440 ;
        RECT 84.380 311.230 85.360 311.460 ;
        RECT 87.850 311.230 88.830 311.460 ;
        RECT 91.320 311.230 92.300 311.460 ;
        RECT 97.800 311.450 98.780 311.680 ;
        RECT 101.270 311.450 102.250 311.680 ;
        RECT 211.890 309.420 212.870 309.650 ;
        RECT 215.360 309.420 216.340 309.650 ;
        RECT 218.830 309.420 219.810 309.650 ;
        RECT 222.300 309.420 223.280 309.650 ;
        RECT 225.770 309.420 226.750 309.650 ;
        RECT 231.930 309.410 232.910 309.640 ;
        RECT 235.400 309.410 236.380 309.640 ;
        RECT 238.870 309.410 239.850 309.640 ;
        RECT 242.340 309.410 243.320 309.640 ;
        RECT 245.810 309.410 246.790 309.640 ;
        RECT 251.990 309.410 252.970 309.640 ;
        RECT 255.460 309.410 256.440 309.640 ;
        RECT 258.930 309.410 259.910 309.640 ;
        RECT 262.400 309.410 263.380 309.640 ;
        RECT 265.870 309.410 266.850 309.640 ;
        RECT 272.040 309.410 273.020 309.640 ;
        RECT 275.510 309.410 276.490 309.640 ;
        RECT 278.980 309.410 279.960 309.640 ;
        RECT 282.450 309.410 283.430 309.640 ;
        RECT 285.920 309.410 286.900 309.640 ;
        RECT 4.770 307.910 5.750 308.140 ;
        RECT 8.240 307.910 9.220 308.140 ;
        RECT 11.710 307.910 12.690 308.140 ;
        RECT 18.110 307.890 19.090 308.120 ;
        RECT 21.580 307.890 22.560 308.120 ;
        RECT 25.050 307.890 26.030 308.120 ;
        RECT 31.480 307.920 32.460 308.150 ;
        RECT 34.950 307.920 35.930 308.150 ;
        RECT 38.420 307.920 39.400 308.150 ;
        RECT 44.710 307.920 45.690 308.150 ;
        RECT 48.180 307.920 49.160 308.150 ;
        RECT 51.650 307.920 52.630 308.150 ;
        RECT 57.980 307.890 58.960 308.120 ;
        RECT 61.450 307.890 62.430 308.120 ;
        RECT 64.920 307.890 65.900 308.120 ;
        RECT 71.250 307.920 72.230 308.150 ;
        RECT 74.720 307.920 75.700 308.150 ;
        RECT 78.190 307.920 79.170 308.150 ;
        RECT 84.380 307.940 85.360 308.170 ;
        RECT 87.850 307.940 88.830 308.170 ;
        RECT 91.320 307.940 92.300 308.170 ;
        RECT 97.800 308.160 98.780 308.390 ;
        RECT 101.270 308.160 102.250 308.390 ;
        RECT 15.400 305.100 16.550 305.410 ;
        RECT 28.570 305.100 29.810 305.580 ;
        RECT 41.870 305.310 42.940 305.960 ;
        RECT 11.980 304.850 16.550 305.100 ;
        RECT 4.770 304.620 5.750 304.850 ;
        RECT 8.240 304.620 9.220 304.850 ;
        RECT 11.710 304.620 16.550 304.850 ;
        RECT 25.530 304.830 29.810 305.100 ;
        RECT 38.740 304.860 42.940 305.310 ;
        RECT 55.250 305.050 56.400 305.540 ;
        RECT 52.040 304.860 56.400 305.050 ;
        RECT 68.500 305.010 69.400 305.700 ;
        RECT 81.580 305.140 82.910 305.410 ;
        RECT 94.330 305.260 95.440 305.870 ;
        RECT 11.980 304.300 16.550 304.620 ;
        RECT 18.110 304.600 19.090 304.830 ;
        RECT 21.580 304.600 22.560 304.830 ;
        RECT 25.050 304.600 29.810 304.830 ;
        RECT 31.480 304.630 32.460 304.860 ;
        RECT 34.950 304.630 35.930 304.860 ;
        RECT 38.420 304.630 42.940 304.860 ;
        RECT 44.710 304.630 45.690 304.860 ;
        RECT 48.180 304.630 49.160 304.860 ;
        RECT 51.650 304.630 56.400 304.860 ;
        RECT 65.080 304.830 69.400 305.010 ;
        RECT 78.460 304.860 82.910 305.140 ;
        RECT 91.590 304.880 95.440 305.260 ;
        RECT 15.400 303.520 16.550 304.300 ;
        RECT 25.530 304.260 29.810 304.600 ;
        RECT 28.570 303.650 29.810 304.260 ;
        RECT 38.740 304.130 42.940 304.630 ;
        RECT 41.870 303.400 42.940 304.130 ;
        RECT 52.040 304.090 56.400 304.630 ;
        RECT 57.980 304.600 58.960 304.830 ;
        RECT 61.450 304.600 62.430 304.830 ;
        RECT 64.920 304.600 69.400 304.830 ;
        RECT 71.250 304.630 72.230 304.860 ;
        RECT 74.720 304.630 75.700 304.860 ;
        RECT 78.190 304.630 82.910 304.860 ;
        RECT 84.380 304.650 85.360 304.880 ;
        RECT 87.850 304.650 88.830 304.880 ;
        RECT 91.320 304.650 95.440 304.880 ;
        RECT 97.800 304.870 98.780 305.100 ;
        RECT 101.270 304.870 102.250 305.100 ;
        RECT 65.080 304.420 69.400 304.600 ;
        RECT 78.460 304.550 82.910 304.630 ;
        RECT 55.250 303.230 56.400 304.090 ;
        RECT 68.500 303.440 69.400 304.420 ;
        RECT 81.580 303.940 82.910 304.550 ;
        RECT 91.590 304.470 95.440 304.650 ;
        RECT 94.330 304.020 95.440 304.470 ;
        RECT 213.630 304.440 226.860 304.490 ;
        RECT 207.020 304.170 226.860 304.440 ;
        RECT 205.530 303.790 226.860 304.170 ;
        RECT 233.600 303.790 246.830 304.490 ;
        RECT 253.710 303.790 266.940 304.490 ;
        RECT 273.820 303.790 287.050 304.490 ;
        RECT 205.530 302.870 287.050 303.790 ;
        RECT 205.530 302.480 226.860 302.870 ;
        RECT 233.600 302.480 246.830 302.870 ;
        RECT 253.710 302.480 266.940 302.870 ;
        RECT 273.820 302.480 287.050 302.870 ;
        RECT 205.530 302.160 216.800 302.480 ;
        RECT 4.770 301.330 5.750 301.560 ;
        RECT 8.240 301.330 9.220 301.560 ;
        RECT 11.710 301.330 12.690 301.560 ;
        RECT 18.110 301.310 19.090 301.540 ;
        RECT 21.580 301.310 22.560 301.540 ;
        RECT 25.050 301.310 26.030 301.540 ;
        RECT 31.480 301.340 32.460 301.570 ;
        RECT 34.950 301.340 35.930 301.570 ;
        RECT 38.420 301.340 39.400 301.570 ;
        RECT 44.710 301.340 45.690 301.570 ;
        RECT 48.180 301.340 49.160 301.570 ;
        RECT 51.650 301.340 52.630 301.570 ;
        RECT 57.980 301.310 58.960 301.540 ;
        RECT 61.450 301.310 62.430 301.540 ;
        RECT 64.920 301.310 65.900 301.540 ;
        RECT 71.250 301.340 72.230 301.570 ;
        RECT 74.720 301.340 75.700 301.570 ;
        RECT 78.190 301.340 79.170 301.570 ;
        RECT 84.380 301.360 85.360 301.590 ;
        RECT 87.850 301.360 88.830 301.590 ;
        RECT 91.320 301.360 92.300 301.590 ;
        RECT 97.800 301.580 98.780 301.810 ;
        RECT 101.270 301.580 102.250 301.810 ;
        RECT 9.000 298.870 97.390 299.130 ;
        RECT 1.170 298.630 97.390 298.870 ;
        RECT 1.170 297.980 103.000 298.630 ;
        RECT 1.170 297.450 12.880 297.980 ;
        RECT 1.170 297.310 10.740 297.450 ;
        RECT 18.060 297.430 26.220 297.980 ;
        RECT 31.430 297.460 39.590 297.980 ;
        RECT 44.660 297.460 52.820 297.980 ;
        RECT 57.930 297.430 66.090 297.980 ;
        RECT 71.200 297.460 79.360 297.980 ;
        RECT 84.330 297.480 92.490 297.980 ;
        RECT 1.170 289.370 2.470 297.310 ;
        RECT 96.820 297.280 103.000 297.980 ;
        RECT 4.630 293.020 5.610 293.250 ;
        RECT 8.100 293.020 9.080 293.250 ;
        RECT 11.570 293.020 12.550 293.250 ;
        RECT 17.970 293.000 18.950 293.230 ;
        RECT 21.440 293.000 22.420 293.230 ;
        RECT 24.910 293.000 25.890 293.230 ;
        RECT 31.340 293.030 32.320 293.260 ;
        RECT 34.810 293.030 35.790 293.260 ;
        RECT 38.280 293.030 39.260 293.260 ;
        RECT 44.570 293.030 45.550 293.260 ;
        RECT 48.040 293.030 49.020 293.260 ;
        RECT 51.510 293.030 52.490 293.260 ;
        RECT 57.840 293.000 58.820 293.230 ;
        RECT 61.310 293.000 62.290 293.230 ;
        RECT 64.780 293.000 65.760 293.230 ;
        RECT 71.110 293.030 72.090 293.260 ;
        RECT 74.580 293.030 75.560 293.260 ;
        RECT 78.050 293.030 79.030 293.260 ;
        RECT 84.240 293.050 85.220 293.280 ;
        RECT 87.710 293.050 88.690 293.280 ;
        RECT 91.180 293.050 92.160 293.280 ;
        RECT 97.660 293.270 98.640 293.500 ;
        RECT 101.130 293.270 102.110 293.500 ;
        RECT 1.110 282.760 2.770 289.370 ;
        RECT 4.630 286.440 5.610 286.670 ;
        RECT 8.100 286.440 9.080 286.670 ;
        RECT 11.570 286.440 12.550 286.670 ;
        RECT 17.970 286.420 18.950 286.650 ;
        RECT 21.440 286.420 22.420 286.650 ;
        RECT 24.910 286.420 25.890 286.650 ;
        RECT 31.340 286.450 32.320 286.680 ;
        RECT 34.810 286.450 35.790 286.680 ;
        RECT 38.280 286.450 39.260 286.680 ;
        RECT 44.570 286.450 45.550 286.680 ;
        RECT 48.040 286.450 49.020 286.680 ;
        RECT 51.510 286.450 52.490 286.680 ;
        RECT 57.840 286.420 58.820 286.650 ;
        RECT 61.310 286.420 62.290 286.650 ;
        RECT 64.780 286.420 65.760 286.650 ;
        RECT 71.110 286.450 72.090 286.680 ;
        RECT 74.580 286.450 75.560 286.680 ;
        RECT 78.050 286.450 79.030 286.680 ;
        RECT 84.240 286.470 85.220 286.700 ;
        RECT 87.710 286.470 88.690 286.700 ;
        RECT 91.180 286.470 92.160 286.700 ;
        RECT 97.660 286.690 98.640 286.920 ;
        RECT 101.130 286.690 102.110 286.920 ;
        RECT 1.170 267.250 2.470 282.760 ;
        RECT 205.530 282.300 208.350 302.160 ;
        RECT 211.850 301.590 212.830 301.820 ;
        RECT 215.320 301.590 216.300 301.820 ;
        RECT 218.790 301.590 219.770 301.820 ;
        RECT 222.260 301.590 223.240 301.820 ;
        RECT 225.730 301.590 226.710 301.820 ;
        RECT 231.820 301.590 232.800 301.820 ;
        RECT 235.290 301.590 236.270 301.820 ;
        RECT 238.760 301.590 239.740 301.820 ;
        RECT 242.230 301.590 243.210 301.820 ;
        RECT 245.700 301.590 246.680 301.820 ;
        RECT 251.930 301.590 252.910 301.820 ;
        RECT 255.400 301.590 256.380 301.820 ;
        RECT 258.870 301.590 259.850 301.820 ;
        RECT 262.340 301.590 263.320 301.820 ;
        RECT 265.810 301.590 266.790 301.820 ;
        RECT 272.040 301.590 273.020 301.820 ;
        RECT 275.510 301.590 276.490 301.820 ;
        RECT 278.980 301.590 279.960 301.820 ;
        RECT 282.450 301.590 283.430 301.820 ;
        RECT 285.920 301.590 286.900 301.820 ;
        RECT 211.850 295.010 212.830 295.240 ;
        RECT 215.320 295.010 216.300 295.240 ;
        RECT 218.790 295.010 219.770 295.240 ;
        RECT 222.260 295.010 223.240 295.240 ;
        RECT 225.730 295.010 226.710 295.240 ;
        RECT 231.820 295.010 232.800 295.240 ;
        RECT 235.290 295.010 236.270 295.240 ;
        RECT 238.760 295.010 239.740 295.240 ;
        RECT 242.230 295.010 243.210 295.240 ;
        RECT 245.700 295.010 246.680 295.240 ;
        RECT 251.930 295.010 252.910 295.240 ;
        RECT 255.400 295.010 256.380 295.240 ;
        RECT 258.870 295.010 259.850 295.240 ;
        RECT 262.340 295.010 263.320 295.240 ;
        RECT 265.810 295.010 266.790 295.240 ;
        RECT 272.040 295.010 273.020 295.240 ;
        RECT 275.510 295.010 276.490 295.240 ;
        RECT 278.980 295.010 279.960 295.240 ;
        RECT 282.450 295.010 283.430 295.240 ;
        RECT 285.920 295.010 286.900 295.240 ;
        RECT 355.040 294.780 356.120 309.080 ;
        RECT 356.500 308.160 356.730 309.140 ;
        RECT 359.790 308.160 360.020 309.140 ;
        RECT 363.080 308.160 363.310 309.140 ;
        RECT 366.300 308.540 366.680 313.880 ;
        RECT 369.660 313.100 369.890 314.080 ;
        RECT 374.360 313.500 375.440 327.800 ;
        RECT 375.820 326.880 376.050 327.860 ;
        RECT 382.400 326.880 382.630 327.860 ;
        RECT 388.980 326.880 389.210 327.860 ;
        RECT 375.820 323.410 376.050 324.390 ;
        RECT 382.400 323.410 382.630 324.390 ;
        RECT 388.980 323.410 389.210 324.390 ;
        RECT 375.820 319.940 376.050 320.920 ;
        RECT 382.400 319.940 382.630 320.920 ;
        RECT 388.980 319.940 389.210 320.920 ;
        RECT 375.820 316.470 376.050 317.450 ;
        RECT 382.400 316.470 382.630 317.450 ;
        RECT 388.980 316.470 389.210 317.450 ;
        RECT 366.370 308.160 366.600 308.540 ;
        RECT 369.660 308.160 369.890 309.140 ;
        RECT 374.370 308.980 374.950 313.500 ;
        RECT 375.820 313.000 376.050 313.980 ;
        RECT 382.400 313.000 382.630 313.980 ;
        RECT 388.980 313.000 389.210 313.980 ;
        RECT 393.610 313.570 394.690 327.870 ;
        RECT 395.070 326.950 395.300 327.930 ;
        RECT 398.360 326.950 398.590 327.930 ;
        RECT 401.650 326.950 401.880 327.930 ;
        RECT 404.760 327.360 405.380 332.350 ;
        RECT 408.230 331.920 408.460 332.900 ;
        RECT 404.940 326.950 405.170 327.360 ;
        RECT 408.230 326.950 408.460 327.930 ;
        RECT 395.070 323.480 395.300 324.460 ;
        RECT 398.360 323.480 398.590 324.460 ;
        RECT 401.650 323.480 401.880 324.460 ;
        RECT 404.940 323.480 405.170 324.460 ;
        RECT 408.230 323.480 408.460 324.460 ;
        RECT 395.070 320.010 395.300 320.990 ;
        RECT 398.360 320.010 398.590 320.990 ;
        RECT 401.650 320.010 401.880 320.990 ;
        RECT 404.940 320.010 405.170 320.990 ;
        RECT 408.230 320.010 408.460 320.990 ;
        RECT 395.070 316.540 395.300 317.520 ;
        RECT 398.360 316.540 398.590 317.520 ;
        RECT 401.650 316.540 401.880 317.520 ;
        RECT 404.940 316.540 405.170 317.520 ;
        RECT 408.230 316.540 408.460 317.520 ;
        RECT 393.730 309.050 394.310 313.570 ;
        RECT 395.070 313.070 395.300 314.050 ;
        RECT 398.360 313.070 398.590 314.050 ;
        RECT 401.650 313.070 401.880 314.050 ;
        RECT 404.940 313.850 405.170 314.050 ;
        RECT 356.500 304.690 356.730 305.670 ;
        RECT 359.790 304.690 360.020 305.670 ;
        RECT 363.080 304.690 363.310 305.670 ;
        RECT 366.370 304.690 366.600 305.670 ;
        RECT 369.660 304.690 369.890 305.670 ;
        RECT 356.500 301.220 356.730 302.200 ;
        RECT 359.790 301.220 360.020 302.200 ;
        RECT 363.080 301.220 363.310 302.200 ;
        RECT 366.370 301.220 366.600 302.200 ;
        RECT 369.660 301.220 369.890 302.200 ;
        RECT 356.500 297.750 356.730 298.730 ;
        RECT 359.790 297.750 360.020 298.730 ;
        RECT 363.080 297.750 363.310 298.730 ;
        RECT 366.370 297.750 366.600 298.730 ;
        RECT 369.660 297.750 369.890 298.730 ;
        RECT 356.500 294.280 356.730 295.260 ;
        RECT 359.790 294.280 360.020 295.260 ;
        RECT 363.080 294.280 363.310 295.260 ;
        RECT 366.370 295.030 366.600 295.260 ;
        RECT 211.850 288.430 212.830 288.660 ;
        RECT 215.320 288.430 216.300 288.660 ;
        RECT 218.790 288.430 219.770 288.660 ;
        RECT 222.260 288.430 223.240 288.660 ;
        RECT 225.730 288.430 226.710 288.660 ;
        RECT 231.820 288.430 232.800 288.660 ;
        RECT 235.290 288.430 236.270 288.660 ;
        RECT 238.760 288.430 239.740 288.660 ;
        RECT 242.230 288.430 243.210 288.660 ;
        RECT 245.700 288.430 246.680 288.660 ;
        RECT 251.930 288.430 252.910 288.660 ;
        RECT 255.400 288.430 256.380 288.660 ;
        RECT 258.870 288.430 259.850 288.660 ;
        RECT 262.340 288.430 263.320 288.660 ;
        RECT 265.810 288.430 266.790 288.660 ;
        RECT 272.040 288.430 273.020 288.660 ;
        RECT 275.510 288.430 276.490 288.660 ;
        RECT 278.980 288.430 279.960 288.660 ;
        RECT 282.450 288.430 283.430 288.660 ;
        RECT 285.920 288.430 286.900 288.660 ;
        RECT 213.390 282.300 226.620 282.540 ;
        RECT 205.530 281.770 226.620 282.300 ;
        RECT 233.430 281.770 246.660 282.530 ;
        RECT 253.490 281.770 266.720 282.530 ;
        RECT 273.540 281.770 286.770 282.530 ;
        RECT 205.530 280.850 286.770 281.770 ;
        RECT 205.530 280.690 226.620 280.850 ;
        RECT 213.390 280.530 226.620 280.690 ;
        RECT 233.430 280.520 246.660 280.850 ;
        RECT 253.490 280.520 266.720 280.850 ;
        RECT 273.540 280.520 286.770 280.850 ;
        RECT 4.630 279.860 5.610 280.090 ;
        RECT 8.100 279.860 9.080 280.090 ;
        RECT 11.570 279.860 12.550 280.090 ;
        RECT 17.970 279.840 18.950 280.070 ;
        RECT 21.440 279.840 22.420 280.070 ;
        RECT 24.910 279.840 25.890 280.070 ;
        RECT 31.340 279.870 32.320 280.100 ;
        RECT 34.810 279.870 35.790 280.100 ;
        RECT 38.280 279.870 39.260 280.100 ;
        RECT 44.570 279.870 45.550 280.100 ;
        RECT 48.040 279.870 49.020 280.100 ;
        RECT 51.510 279.870 52.490 280.100 ;
        RECT 57.840 279.840 58.820 280.070 ;
        RECT 61.310 279.840 62.290 280.070 ;
        RECT 64.780 279.840 65.760 280.070 ;
        RECT 71.110 279.870 72.090 280.100 ;
        RECT 74.580 279.870 75.560 280.100 ;
        RECT 78.050 279.870 79.030 280.100 ;
        RECT 84.240 279.890 85.220 280.120 ;
        RECT 87.710 279.890 88.690 280.120 ;
        RECT 91.180 279.890 92.160 280.120 ;
        RECT 97.660 280.110 98.640 280.340 ;
        RECT 101.130 280.110 102.110 280.340 ;
        RECT 211.610 279.640 212.590 279.870 ;
        RECT 215.080 279.640 216.060 279.870 ;
        RECT 218.550 279.640 219.530 279.870 ;
        RECT 222.020 279.640 223.000 279.870 ;
        RECT 225.490 279.640 226.470 279.870 ;
        RECT 285.750 279.860 286.680 280.520 ;
        RECT 231.650 279.630 232.630 279.860 ;
        RECT 235.120 279.630 236.100 279.860 ;
        RECT 238.590 279.630 239.570 279.860 ;
        RECT 242.060 279.630 243.040 279.860 ;
        RECT 245.530 279.630 246.510 279.860 ;
        RECT 251.710 279.630 252.690 279.860 ;
        RECT 255.180 279.630 256.160 279.860 ;
        RECT 258.650 279.630 259.630 279.860 ;
        RECT 262.120 279.630 263.100 279.860 ;
        RECT 265.590 279.630 266.570 279.860 ;
        RECT 271.760 279.630 272.740 279.860 ;
        RECT 275.230 279.630 276.210 279.860 ;
        RECT 278.700 279.630 279.680 279.860 ;
        RECT 282.170 279.630 283.150 279.860 ;
        RECT 285.640 279.680 286.680 279.860 ;
        RECT 285.640 279.630 286.620 279.680 ;
        RECT 211.610 276.350 212.590 276.580 ;
        RECT 215.080 276.350 216.060 276.580 ;
        RECT 218.550 276.350 219.530 276.580 ;
        RECT 222.020 276.350 223.000 276.580 ;
        RECT 225.490 276.350 226.470 276.580 ;
        RECT 231.650 276.340 232.630 276.570 ;
        RECT 235.120 276.340 236.100 276.570 ;
        RECT 238.590 276.340 239.570 276.570 ;
        RECT 242.060 276.340 243.040 276.570 ;
        RECT 245.530 276.340 246.510 276.570 ;
        RECT 251.710 276.340 252.690 276.570 ;
        RECT 255.180 276.340 256.160 276.570 ;
        RECT 258.650 276.340 259.630 276.570 ;
        RECT 262.120 276.340 263.100 276.570 ;
        RECT 265.590 276.340 266.570 276.570 ;
        RECT 271.760 276.340 272.740 276.570 ;
        RECT 275.230 276.340 276.210 276.570 ;
        RECT 278.700 276.340 279.680 276.570 ;
        RECT 282.170 276.340 283.150 276.570 ;
        RECT 285.640 276.340 286.620 276.570 ;
        RECT 355.040 275.900 356.120 290.200 ;
        RECT 356.500 289.280 356.730 290.260 ;
        RECT 359.790 289.280 360.020 290.260 ;
        RECT 363.080 289.280 363.310 290.260 ;
        RECT 366.300 289.690 366.680 295.030 ;
        RECT 369.660 294.280 369.890 295.260 ;
        RECT 374.360 294.680 375.440 308.980 ;
        RECT 375.820 308.060 376.050 309.040 ;
        RECT 382.400 308.060 382.630 309.040 ;
        RECT 388.980 308.060 389.210 309.040 ;
        RECT 375.820 304.590 376.050 305.570 ;
        RECT 382.400 304.590 382.630 305.570 ;
        RECT 388.980 304.590 389.210 305.570 ;
        RECT 375.820 301.120 376.050 302.100 ;
        RECT 382.400 301.120 382.630 302.100 ;
        RECT 388.980 301.120 389.210 302.100 ;
        RECT 375.820 297.650 376.050 298.630 ;
        RECT 382.400 297.650 382.630 298.630 ;
        RECT 388.980 297.650 389.210 298.630 ;
        RECT 366.370 289.280 366.600 289.690 ;
        RECT 369.660 289.280 369.890 290.260 ;
        RECT 374.370 290.100 374.950 294.680 ;
        RECT 375.820 294.180 376.050 295.160 ;
        RECT 382.400 294.180 382.630 295.160 ;
        RECT 388.980 294.180 389.210 295.160 ;
        RECT 393.610 294.750 394.690 309.050 ;
        RECT 395.070 308.130 395.300 309.110 ;
        RECT 398.360 308.130 398.590 309.110 ;
        RECT 401.650 308.130 401.880 309.110 ;
        RECT 404.870 308.510 405.250 313.850 ;
        RECT 408.230 313.070 408.460 314.050 ;
        RECT 404.940 308.130 405.170 308.510 ;
        RECT 408.230 308.130 408.460 309.110 ;
        RECT 395.070 304.660 395.300 305.640 ;
        RECT 398.360 304.660 398.590 305.640 ;
        RECT 401.650 304.660 401.880 305.640 ;
        RECT 404.940 304.660 405.170 305.640 ;
        RECT 408.230 304.660 408.460 305.640 ;
        RECT 395.070 301.190 395.300 302.170 ;
        RECT 398.360 301.190 398.590 302.170 ;
        RECT 401.650 301.190 401.880 302.170 ;
        RECT 404.940 301.190 405.170 302.170 ;
        RECT 408.230 301.190 408.460 302.170 ;
        RECT 395.070 297.720 395.300 298.700 ;
        RECT 398.360 297.720 398.590 298.700 ;
        RECT 401.650 297.720 401.880 298.700 ;
        RECT 404.940 297.720 405.170 298.700 ;
        RECT 408.230 297.720 408.460 298.700 ;
        RECT 393.730 290.170 394.310 294.750 ;
        RECT 395.070 294.250 395.300 295.230 ;
        RECT 398.360 294.250 398.590 295.230 ;
        RECT 401.650 294.250 401.880 295.230 ;
        RECT 404.940 295.000 405.170 295.230 ;
        RECT 356.500 285.810 356.730 286.790 ;
        RECT 359.790 285.810 360.020 286.790 ;
        RECT 363.080 285.810 363.310 286.790 ;
        RECT 366.370 285.810 366.600 286.790 ;
        RECT 369.660 285.810 369.890 286.790 ;
        RECT 356.500 282.340 356.730 283.320 ;
        RECT 359.790 282.340 360.020 283.320 ;
        RECT 363.080 282.340 363.310 283.320 ;
        RECT 366.370 282.340 366.600 283.320 ;
        RECT 369.660 282.340 369.890 283.320 ;
        RECT 356.500 278.870 356.730 279.850 ;
        RECT 359.790 278.870 360.020 279.850 ;
        RECT 363.080 278.870 363.310 279.850 ;
        RECT 366.370 278.870 366.600 279.850 ;
        RECT 369.660 278.870 369.890 279.850 ;
        RECT 356.500 275.400 356.730 276.380 ;
        RECT 359.790 275.400 360.020 276.380 ;
        RECT 363.080 275.400 363.310 276.380 ;
        RECT 366.370 276.130 366.600 276.380 ;
        RECT 15.260 273.760 16.410 274.070 ;
        RECT 28.430 273.760 29.670 274.240 ;
        RECT 41.730 273.970 42.800 274.620 ;
        RECT 11.840 273.510 16.410 273.760 ;
        RECT 4.630 273.280 5.610 273.510 ;
        RECT 8.100 273.280 9.080 273.510 ;
        RECT 11.570 273.280 16.410 273.510 ;
        RECT 25.390 273.490 29.670 273.760 ;
        RECT 38.600 273.520 42.800 273.970 ;
        RECT 55.110 273.710 56.260 274.200 ;
        RECT 51.900 273.520 56.260 273.710 ;
        RECT 68.360 273.670 69.260 274.360 ;
        RECT 81.440 273.800 82.770 274.070 ;
        RECT 94.190 273.920 95.300 274.530 ;
        RECT 11.840 272.960 16.410 273.280 ;
        RECT 17.970 273.260 18.950 273.490 ;
        RECT 21.440 273.260 22.420 273.490 ;
        RECT 24.910 273.260 29.670 273.490 ;
        RECT 31.340 273.290 32.320 273.520 ;
        RECT 34.810 273.290 35.790 273.520 ;
        RECT 38.280 273.290 42.800 273.520 ;
        RECT 44.570 273.290 45.550 273.520 ;
        RECT 48.040 273.290 49.020 273.520 ;
        RECT 51.510 273.290 56.260 273.520 ;
        RECT 64.940 273.490 69.260 273.670 ;
        RECT 78.320 273.520 82.770 273.800 ;
        RECT 91.450 273.540 95.300 273.920 ;
        RECT 15.260 272.180 16.410 272.960 ;
        RECT 25.390 272.920 29.670 273.260 ;
        RECT 28.430 272.310 29.670 272.920 ;
        RECT 38.600 272.790 42.800 273.290 ;
        RECT 41.730 272.060 42.800 272.790 ;
        RECT 51.900 272.750 56.260 273.290 ;
        RECT 57.840 273.260 58.820 273.490 ;
        RECT 61.310 273.260 62.290 273.490 ;
        RECT 64.780 273.260 69.260 273.490 ;
        RECT 71.110 273.290 72.090 273.520 ;
        RECT 74.580 273.290 75.560 273.520 ;
        RECT 78.050 273.290 82.770 273.520 ;
        RECT 84.240 273.310 85.220 273.540 ;
        RECT 87.710 273.310 88.690 273.540 ;
        RECT 91.180 273.310 95.300 273.540 ;
        RECT 97.660 273.530 98.640 273.760 ;
        RECT 101.130 273.530 102.110 273.760 ;
        RECT 64.940 273.080 69.260 273.260 ;
        RECT 78.320 273.210 82.770 273.290 ;
        RECT 55.110 271.890 56.260 272.750 ;
        RECT 68.360 272.100 69.260 273.080 ;
        RECT 81.440 272.600 82.770 273.210 ;
        RECT 91.450 273.130 95.300 273.310 ;
        RECT 93.580 272.680 95.300 273.130 ;
        RECT 211.610 273.060 212.590 273.290 ;
        RECT 215.080 273.060 216.060 273.290 ;
        RECT 218.550 273.060 219.530 273.290 ;
        RECT 222.020 273.060 223.000 273.290 ;
        RECT 225.490 273.060 226.470 273.290 ;
        RECT 231.650 273.050 232.630 273.280 ;
        RECT 235.120 273.050 236.100 273.280 ;
        RECT 238.590 273.050 239.570 273.280 ;
        RECT 242.060 273.050 243.040 273.280 ;
        RECT 245.530 273.050 246.510 273.280 ;
        RECT 251.710 273.050 252.690 273.280 ;
        RECT 255.180 273.050 256.160 273.280 ;
        RECT 258.650 273.050 259.630 273.280 ;
        RECT 262.120 273.050 263.100 273.280 ;
        RECT 265.590 273.050 266.570 273.280 ;
        RECT 271.760 273.050 272.740 273.280 ;
        RECT 275.230 273.050 276.210 273.280 ;
        RECT 278.700 273.050 279.680 273.280 ;
        RECT 282.170 273.050 283.150 273.280 ;
        RECT 285.640 273.050 286.620 273.280 ;
        RECT 93.580 268.630 94.330 272.680 ;
        RECT 211.610 269.770 212.590 270.000 ;
        RECT 215.080 269.770 216.060 270.000 ;
        RECT 218.550 269.770 219.530 270.000 ;
        RECT 222.020 269.770 223.000 270.000 ;
        RECT 225.490 269.770 226.470 270.000 ;
        RECT 231.650 269.760 232.630 269.990 ;
        RECT 235.120 269.760 236.100 269.990 ;
        RECT 238.590 269.760 239.570 269.990 ;
        RECT 242.060 269.760 243.040 269.990 ;
        RECT 245.530 269.760 246.510 269.990 ;
        RECT 251.710 269.760 252.690 269.990 ;
        RECT 255.180 269.760 256.160 269.990 ;
        RECT 258.650 269.760 259.630 269.990 ;
        RECT 262.120 269.760 263.100 269.990 ;
        RECT 265.590 269.760 266.570 269.990 ;
        RECT 271.760 269.760 272.740 269.990 ;
        RECT 275.230 269.760 276.210 269.990 ;
        RECT 278.700 269.760 279.680 269.990 ;
        RECT 282.170 269.760 283.150 269.990 ;
        RECT 285.640 269.760 286.620 269.990 ;
        RECT 1.170 266.640 10.610 267.250 ;
        RECT 1.170 266.560 12.880 266.640 ;
        RECT 18.060 266.560 26.220 266.620 ;
        RECT 31.430 266.560 39.590 266.650 ;
        RECT 44.660 266.560 52.820 266.650 ;
        RECT 57.930 266.560 66.090 266.620 ;
        RECT 71.200 266.560 79.360 266.650 ;
        RECT 84.330 266.560 92.490 266.670 ;
        RECT 96.820 266.560 103.000 266.800 ;
        RECT 1.170 265.690 103.000 266.560 ;
        RECT 211.610 266.480 212.590 266.710 ;
        RECT 215.080 266.480 216.060 266.710 ;
        RECT 218.550 266.480 219.530 266.710 ;
        RECT 222.020 266.480 223.000 266.710 ;
        RECT 225.490 266.480 226.470 266.710 ;
        RECT 231.650 266.470 232.630 266.700 ;
        RECT 235.120 266.470 236.100 266.700 ;
        RECT 238.590 266.470 239.570 266.700 ;
        RECT 242.060 266.470 243.040 266.700 ;
        RECT 245.530 266.470 246.510 266.700 ;
        RECT 251.710 266.470 252.690 266.700 ;
        RECT 255.180 266.470 256.160 266.700 ;
        RECT 258.650 266.470 259.630 266.700 ;
        RECT 262.120 266.470 263.100 266.700 ;
        RECT 265.590 266.470 266.570 266.700 ;
        RECT 271.760 266.470 272.740 266.700 ;
        RECT 275.230 266.470 276.210 266.700 ;
        RECT 278.700 266.470 279.680 266.700 ;
        RECT 282.170 266.470 283.150 266.700 ;
        RECT 285.640 266.470 286.620 266.700 ;
        RECT -46.180 236.630 -32.570 239.310 ;
        RECT 1.170 237.320 2.470 265.690 ;
        RECT 4.720 265.620 103.000 265.690 ;
        RECT 9.840 265.450 103.000 265.620 ;
        RECT 9.840 265.410 98.230 265.450 ;
        RECT 4.630 264.480 5.610 264.710 ;
        RECT 8.100 264.480 9.080 264.710 ;
        RECT 11.570 264.480 12.550 264.710 ;
        RECT 17.970 264.460 18.950 264.690 ;
        RECT 21.440 264.460 22.420 264.690 ;
        RECT 24.910 264.460 25.890 264.690 ;
        RECT 31.340 264.490 32.320 264.720 ;
        RECT 34.810 264.490 35.790 264.720 ;
        RECT 38.280 264.490 39.260 264.720 ;
        RECT 44.570 264.490 45.550 264.720 ;
        RECT 48.040 264.490 49.020 264.720 ;
        RECT 51.510 264.490 52.490 264.720 ;
        RECT 57.840 264.460 58.820 264.690 ;
        RECT 61.310 264.460 62.290 264.690 ;
        RECT 64.780 264.460 65.760 264.690 ;
        RECT 71.110 264.490 72.090 264.720 ;
        RECT 74.580 264.490 75.560 264.720 ;
        RECT 78.050 264.490 79.030 264.720 ;
        RECT 84.240 264.510 85.220 264.740 ;
        RECT 87.710 264.510 88.690 264.740 ;
        RECT 91.180 264.510 92.160 264.740 ;
        RECT 97.660 264.730 98.640 264.960 ;
        RECT 101.130 264.730 102.110 264.960 ;
        RECT 211.610 263.190 212.590 263.420 ;
        RECT 215.080 263.190 216.060 263.420 ;
        RECT 218.550 263.190 219.530 263.420 ;
        RECT 222.020 263.190 223.000 263.420 ;
        RECT 225.490 263.190 226.470 263.420 ;
        RECT 231.650 263.180 232.630 263.410 ;
        RECT 235.120 263.180 236.100 263.410 ;
        RECT 238.590 263.180 239.570 263.410 ;
        RECT 242.060 263.180 243.040 263.410 ;
        RECT 245.530 263.180 246.510 263.410 ;
        RECT 251.710 263.180 252.690 263.410 ;
        RECT 255.180 263.180 256.160 263.410 ;
        RECT 258.650 263.180 259.630 263.410 ;
        RECT 262.120 263.180 263.100 263.410 ;
        RECT 265.590 263.180 266.570 263.410 ;
        RECT 271.760 263.180 272.740 263.410 ;
        RECT 275.230 263.180 276.210 263.410 ;
        RECT 278.700 263.180 279.680 263.410 ;
        RECT 282.170 263.180 283.150 263.410 ;
        RECT 285.640 263.180 286.620 263.410 ;
        RECT 4.630 261.190 5.610 261.420 ;
        RECT 8.100 261.190 9.080 261.420 ;
        RECT 11.570 261.190 12.550 261.420 ;
        RECT 17.970 261.170 18.950 261.400 ;
        RECT 21.440 261.170 22.420 261.400 ;
        RECT 24.910 261.170 25.890 261.400 ;
        RECT 31.340 261.200 32.320 261.430 ;
        RECT 34.810 261.200 35.790 261.430 ;
        RECT 38.280 261.200 39.260 261.430 ;
        RECT 44.570 261.200 45.550 261.430 ;
        RECT 48.040 261.200 49.020 261.430 ;
        RECT 51.510 261.200 52.490 261.430 ;
        RECT 57.840 261.170 58.820 261.400 ;
        RECT 61.310 261.170 62.290 261.400 ;
        RECT 64.780 261.170 65.760 261.400 ;
        RECT 71.110 261.200 72.090 261.430 ;
        RECT 74.580 261.200 75.560 261.430 ;
        RECT 78.050 261.200 79.030 261.430 ;
        RECT 84.240 261.220 85.220 261.450 ;
        RECT 87.710 261.220 88.690 261.450 ;
        RECT 91.180 261.220 92.160 261.450 ;
        RECT 97.660 261.440 98.640 261.670 ;
        RECT 101.130 261.440 102.110 261.670 ;
        RECT 213.350 261.340 226.580 261.550 ;
        RECT 233.320 261.340 246.550 261.550 ;
        RECT 253.430 261.340 266.660 261.550 ;
        RECT 273.540 261.340 286.770 261.550 ;
        RECT 213.350 260.900 286.770 261.340 ;
        RECT 288.050 260.900 289.000 262.250 ;
        RECT 213.350 260.420 289.000 260.900 ;
        RECT 213.350 259.540 226.580 260.420 ;
        RECT 233.320 259.540 246.550 260.420 ;
        RECT 253.430 259.540 266.660 260.420 ;
        RECT 273.540 260.300 289.000 260.420 ;
        RECT 273.540 259.540 286.770 260.300 ;
        RECT 288.050 259.540 289.000 260.300 ;
        RECT 211.570 258.650 212.550 258.880 ;
        RECT 215.040 258.650 216.020 258.880 ;
        RECT 218.510 258.650 219.490 258.880 ;
        RECT 221.980 258.650 222.960 258.880 ;
        RECT 225.450 258.650 226.430 258.880 ;
        RECT 231.540 258.650 232.520 258.880 ;
        RECT 235.010 258.650 235.990 258.880 ;
        RECT 238.480 258.650 239.460 258.880 ;
        RECT 241.950 258.650 242.930 258.880 ;
        RECT 245.420 258.650 246.400 258.880 ;
        RECT 251.650 258.650 252.630 258.880 ;
        RECT 255.120 258.650 256.100 258.880 ;
        RECT 258.590 258.650 259.570 258.880 ;
        RECT 262.060 258.650 263.040 258.880 ;
        RECT 265.530 258.650 266.510 258.880 ;
        RECT 271.760 258.650 272.740 258.880 ;
        RECT 275.230 258.650 276.210 258.880 ;
        RECT 278.700 258.650 279.680 258.880 ;
        RECT 282.170 258.650 283.150 258.880 ;
        RECT 285.640 258.650 286.620 258.880 ;
        RECT 4.630 257.900 5.610 258.130 ;
        RECT 8.100 257.900 9.080 258.130 ;
        RECT 11.570 257.900 12.550 258.130 ;
        RECT 17.970 257.880 18.950 258.110 ;
        RECT 21.440 257.880 22.420 258.110 ;
        RECT 24.910 257.880 25.890 258.110 ;
        RECT 31.340 257.910 32.320 258.140 ;
        RECT 34.810 257.910 35.790 258.140 ;
        RECT 38.280 257.910 39.260 258.140 ;
        RECT 44.570 257.910 45.550 258.140 ;
        RECT 48.040 257.910 49.020 258.140 ;
        RECT 51.510 257.910 52.490 258.140 ;
        RECT 57.840 257.880 58.820 258.110 ;
        RECT 61.310 257.880 62.290 258.110 ;
        RECT 64.780 257.880 65.760 258.110 ;
        RECT 71.110 257.910 72.090 258.140 ;
        RECT 74.580 257.910 75.560 258.140 ;
        RECT 78.050 257.910 79.030 258.140 ;
        RECT 84.240 257.930 85.220 258.160 ;
        RECT 87.710 257.930 88.690 258.160 ;
        RECT 91.180 257.930 92.160 258.160 ;
        RECT 97.660 258.150 98.640 258.380 ;
        RECT 101.130 258.150 102.110 258.380 ;
        RECT 355.060 257.040 356.140 271.340 ;
        RECT 356.520 270.420 356.750 271.400 ;
        RECT 359.810 270.420 360.040 271.400 ;
        RECT 363.100 270.420 363.330 271.400 ;
        RECT 366.300 270.790 366.680 276.130 ;
        RECT 369.660 275.400 369.890 276.380 ;
        RECT 374.360 275.800 375.440 290.100 ;
        RECT 375.820 289.180 376.050 290.160 ;
        RECT 382.400 289.180 382.630 290.160 ;
        RECT 388.980 289.180 389.210 290.160 ;
        RECT 375.820 285.710 376.050 286.690 ;
        RECT 382.400 285.710 382.630 286.690 ;
        RECT 388.980 285.710 389.210 286.690 ;
        RECT 375.820 282.240 376.050 283.220 ;
        RECT 382.400 282.240 382.630 283.220 ;
        RECT 388.980 282.240 389.210 283.220 ;
        RECT 375.820 278.770 376.050 279.750 ;
        RECT 382.400 278.770 382.630 279.750 ;
        RECT 388.980 278.770 389.210 279.750 ;
        RECT 366.390 270.420 366.620 270.790 ;
        RECT 369.680 270.420 369.910 271.400 ;
        RECT 374.370 271.240 374.950 275.800 ;
        RECT 375.820 275.300 376.050 276.280 ;
        RECT 382.400 275.300 382.630 276.280 ;
        RECT 388.980 275.300 389.210 276.280 ;
        RECT 393.610 275.870 394.690 290.170 ;
        RECT 395.070 289.250 395.300 290.230 ;
        RECT 398.360 289.250 398.590 290.230 ;
        RECT 401.650 289.250 401.880 290.230 ;
        RECT 404.870 289.660 405.250 295.000 ;
        RECT 408.230 294.250 408.460 295.230 ;
        RECT 404.940 289.250 405.170 289.660 ;
        RECT 408.230 289.250 408.460 290.230 ;
        RECT 395.070 285.780 395.300 286.760 ;
        RECT 398.360 285.780 398.590 286.760 ;
        RECT 401.650 285.780 401.880 286.760 ;
        RECT 404.940 285.780 405.170 286.760 ;
        RECT 408.230 285.780 408.460 286.760 ;
        RECT 395.070 282.310 395.300 283.290 ;
        RECT 398.360 282.310 398.590 283.290 ;
        RECT 401.650 282.310 401.880 283.290 ;
        RECT 404.940 282.310 405.170 283.290 ;
        RECT 408.230 282.310 408.460 283.290 ;
        RECT 395.070 278.840 395.300 279.820 ;
        RECT 398.360 278.840 398.590 279.820 ;
        RECT 401.650 278.840 401.880 279.820 ;
        RECT 404.940 278.840 405.170 279.820 ;
        RECT 408.230 278.840 408.460 279.820 ;
        RECT 393.730 271.310 394.310 275.870 ;
        RECT 395.070 275.370 395.300 276.350 ;
        RECT 398.360 275.370 398.590 276.350 ;
        RECT 401.650 275.370 401.880 276.350 ;
        RECT 404.940 276.100 405.170 276.350 ;
        RECT 374.370 268.500 375.460 271.240 ;
        RECT 375.840 270.320 376.070 271.300 ;
        RECT 382.420 270.320 382.650 271.300 ;
        RECT 389.000 270.320 389.230 271.300 ;
        RECT 356.520 266.950 356.750 267.930 ;
        RECT 359.810 266.950 360.040 267.930 ;
        RECT 363.100 266.950 363.330 267.930 ;
        RECT 366.390 266.950 366.620 267.930 ;
        RECT 369.680 266.950 369.910 267.930 ;
        RECT 356.520 263.480 356.750 264.460 ;
        RECT 359.810 263.480 360.040 264.460 ;
        RECT 363.100 263.480 363.330 264.460 ;
        RECT 366.390 263.480 366.620 264.460 ;
        RECT 369.680 263.480 369.910 264.460 ;
        RECT 356.520 260.010 356.750 260.990 ;
        RECT 359.810 260.010 360.040 260.990 ;
        RECT 363.100 260.010 363.330 260.990 ;
        RECT 366.390 260.010 366.620 260.990 ;
        RECT 369.680 260.010 369.910 260.990 ;
        RECT 356.520 256.540 356.750 257.520 ;
        RECT 359.810 256.540 360.040 257.520 ;
        RECT 363.100 256.540 363.330 257.520 ;
        RECT 366.390 256.540 366.620 257.520 ;
        RECT 369.680 256.540 369.910 257.520 ;
        RECT 374.380 256.940 375.460 268.500 ;
        RECT 375.840 266.850 376.070 267.830 ;
        RECT 382.420 266.850 382.650 267.830 ;
        RECT 389.000 266.850 389.230 267.830 ;
        RECT 375.840 263.380 376.070 264.360 ;
        RECT 382.420 263.380 382.650 264.360 ;
        RECT 389.000 263.380 389.230 264.360 ;
        RECT 375.840 259.910 376.070 260.890 ;
        RECT 382.420 259.910 382.650 260.890 ;
        RECT 389.000 259.910 389.230 260.890 ;
        RECT 375.840 256.440 376.070 257.420 ;
        RECT 382.420 256.440 382.650 257.420 ;
        RECT 389.000 256.440 389.230 257.420 ;
        RECT 393.630 257.010 394.710 271.310 ;
        RECT 395.090 270.390 395.320 271.370 ;
        RECT 398.380 270.390 398.610 271.370 ;
        RECT 401.670 270.390 401.900 271.370 ;
        RECT 404.870 270.760 405.250 276.100 ;
        RECT 408.230 275.370 408.460 276.350 ;
        RECT 409.480 274.770 410.430 379.560 ;
        RECT 470.680 379.360 1085.940 379.560 ;
        RECT 631.350 355.240 635.000 379.360 ;
        RECT 681.280 379.320 766.750 379.360 ;
        RECT 690.920 378.750 766.750 379.320 ;
        RECT 626.590 355.045 654.810 355.240 ;
        RECT 626.590 354.940 655.410 355.045 ;
        RECT 657.550 354.940 672.910 355.035 ;
        RECT 626.590 354.840 672.910 354.940 ;
        RECT 675.600 354.900 690.960 354.995 ;
        RECT 691.520 354.900 692.810 378.750 ;
        RECT 693.190 354.900 708.550 355.015 ;
        RECT 675.600 354.870 708.550 354.900 ;
        RECT 711.040 354.870 726.400 355.015 ;
        RECT 729.300 354.870 744.660 355.015 ;
        RECT 673.870 354.840 674.700 354.850 ;
        RECT 675.600 354.840 744.660 354.870 ;
        RECT 626.590 354.820 744.660 354.840 ;
        RECT 745.200 354.820 746.490 378.750 ;
        RECT 747.070 354.890 762.430 354.985 ;
        RECT 765.110 354.890 780.470 354.905 ;
        RECT 747.070 354.820 780.470 354.890 ;
        RECT 783.270 354.830 798.630 354.945 ;
        RECT 801.650 354.830 817.010 354.955 ;
        RECT 817.840 354.880 819.130 379.360 ;
        RECT 837.490 379.160 850.480 379.360 ;
        RECT 876.770 355.690 878.060 379.360 ;
        RECT 882.500 379.310 1085.940 379.360 ;
        RECT 882.500 378.910 944.550 379.310 ;
        RECT 1072.580 379.180 1085.940 379.310 ;
        RECT 626.590 354.810 780.470 354.820 ;
        RECT 781.260 354.810 782.430 354.820 ;
        RECT 783.270 354.810 817.010 354.830 ;
        RECT 626.590 354.805 817.010 354.810 ;
        RECT 626.590 354.665 658.090 354.805 ;
        RECT 671.510 354.790 817.010 354.805 ;
        RECT 817.790 354.790 819.140 354.880 ;
        RECT 820.450 354.790 835.810 354.935 ;
        RECT 671.510 354.785 835.810 354.790 ;
        RECT 671.510 354.765 694.270 354.785 ;
        RECT 671.510 354.665 676.150 354.765 ;
        RECT 626.590 354.625 676.150 354.665 ;
        RECT 689.630 354.645 694.270 354.765 ;
        RECT 706.730 354.645 711.370 354.785 ;
        RECT 725.580 354.645 730.220 354.785 ;
        RECT 742.870 354.780 835.810 354.785 ;
        RECT 836.990 354.780 837.920 354.840 ;
        RECT 838.920 354.820 840.360 354.915 ;
        RECT 841.420 354.820 878.500 355.690 ;
        RECT 838.920 354.780 878.500 354.820 ;
        RECT 742.870 354.755 878.500 354.780 ;
        RECT 742.870 354.645 747.510 354.755 ;
        RECT 689.630 354.625 747.510 354.645 ;
        RECT 626.590 354.615 747.510 354.625 ;
        RECT 761.210 354.725 878.500 354.755 ;
        RECT 761.210 354.715 802.110 354.725 ;
        RECT 761.210 354.675 784.160 354.715 ;
        RECT 761.210 354.615 765.850 354.675 ;
        RECT 626.590 354.535 765.850 354.615 ;
        RECT 779.520 354.575 784.160 354.675 ;
        RECT 797.470 354.585 802.110 354.715 ;
        RECT 816.400 354.705 878.500 354.725 ;
        RECT 816.400 354.585 821.040 354.705 ;
        RECT 797.470 354.575 821.040 354.585 ;
        RECT 779.520 354.565 821.040 354.575 ;
        RECT 832.110 354.565 832.710 354.705 ;
        RECT 834.830 354.565 878.500 354.705 ;
        RECT 779.520 354.535 878.500 354.565 ;
        RECT 626.590 354.490 878.500 354.535 ;
        RECT 626.590 354.470 655.410 354.490 ;
        RECT 590.450 336.010 591.550 336.270 ;
        RECT 590.450 335.980 601.090 336.010 ;
        RECT 626.600 335.980 627.400 354.470 ;
        RECT 631.350 354.230 635.000 354.470 ;
        RECT 653.970 354.305 655.410 354.470 ;
        RECT 655.990 354.130 656.950 354.490 ;
        RECT 657.550 354.430 690.960 354.490 ;
        RECT 691.520 354.440 692.810 354.490 ;
        RECT 693.190 354.480 878.500 354.490 ;
        RECT 693.190 354.460 762.430 354.480 ;
        RECT 657.550 354.295 672.910 354.430 ;
        RECT 673.870 354.120 674.700 354.430 ;
        RECT 675.600 354.255 690.960 354.430 ;
        RECT 691.530 354.150 692.780 354.440 ;
        RECT 693.190 354.275 708.550 354.460 ;
        RECT 709.230 354.020 710.310 354.460 ;
        RECT 711.040 354.275 726.400 354.460 ;
        RECT 727.330 353.910 728.290 354.460 ;
        RECT 729.300 354.410 762.430 354.460 ;
        RECT 729.300 354.275 744.660 354.410 ;
        RECT 745.200 354.320 746.490 354.410 ;
        RECT 745.210 354.140 746.480 354.320 ;
        RECT 747.070 354.245 762.430 354.410 ;
        RECT 763.250 354.070 764.080 354.480 ;
        RECT 765.110 354.420 878.500 354.480 ;
        RECT 765.110 354.400 798.630 354.420 ;
        RECT 765.110 354.165 780.470 354.400 ;
        RECT 781.260 354.020 782.430 354.400 ;
        RECT 783.270 354.205 798.630 354.400 ;
        RECT 799.490 353.740 800.420 354.420 ;
        RECT 801.650 354.380 878.500 354.420 ;
        RECT 801.650 354.215 817.010 354.380 ;
        RECT 817.790 354.110 819.140 354.380 ;
        RECT 820.450 354.370 878.500 354.380 ;
        RECT 820.450 354.195 835.810 354.370 ;
        RECT 836.990 353.750 837.920 354.370 ;
        RECT 838.920 354.290 878.500 354.370 ;
        RECT 838.920 354.175 840.360 354.290 ;
        RECT 841.420 354.180 878.500 354.290 ;
        RECT 832.020 351.980 832.450 352.350 ;
        RECT 832.090 351.950 832.370 351.980 ;
        RECT 783.830 346.730 787.190 346.775 ;
        RECT 790.390 346.730 791.830 346.805 ;
        RECT 793.850 346.750 809.210 346.865 ;
        RECT 813.210 346.750 828.570 346.775 ;
        RECT 793.850 346.730 828.570 346.750 ;
        RECT 783.830 346.690 828.570 346.730 ;
        RECT 841.630 346.690 841.970 354.180 ;
        RECT 876.770 353.680 878.340 354.180 ;
        RECT 783.830 346.635 842.030 346.690 ;
        RECT 783.830 346.545 794.840 346.635 ;
        RECT 785.340 346.495 794.840 346.545 ;
        RECT 808.120 346.545 842.030 346.635 ;
        RECT 808.120 346.495 813.980 346.545 ;
        RECT 785.340 346.405 813.980 346.495 ;
        RECT 827.570 346.405 842.030 346.545 ;
        RECT 783.830 346.290 842.030 346.405 ;
        RECT 783.830 346.280 809.210 346.290 ;
        RECT 783.830 346.270 791.900 346.280 ;
        RECT 792.440 346.270 809.210 346.280 ;
        RECT 783.830 346.035 787.190 346.270 ;
        RECT 788.280 346.140 789.060 346.270 ;
        RECT 790.390 346.065 791.830 346.270 ;
        RECT 792.440 346.080 793.190 346.270 ;
        RECT 793.850 346.125 809.210 346.270 ;
        RECT 810.590 346.010 811.400 346.290 ;
        RECT 813.210 346.220 842.030 346.290 ;
        RECT 813.210 346.035 828.570 346.220 ;
        RECT 829.180 345.820 829.950 346.220 ;
        RECT 877.150 339.780 878.340 353.680 ;
        RECT 856.860 337.790 878.340 339.780 ;
        RECT 857.280 337.730 878.340 337.790 ;
        RECT 648.630 335.980 649.200 336.040 ;
        RECT 590.450 335.970 631.990 335.980 ;
        RECT 647.740 335.970 653.970 335.980 ;
        RECT 590.450 335.290 656.780 335.970 ;
        RECT 590.450 335.060 591.550 335.290 ;
        RECT 600.500 335.160 656.780 335.290 ;
        RECT 601.180 332.860 601.890 335.160 ;
        RECT 601.180 331.070 601.920 332.860 ;
        RECT 602.590 332.780 602.840 335.160 ;
        RECT 610.280 332.790 610.530 335.160 ;
        RECT 602.590 332.620 606.000 332.780 ;
        RECT 607.140 332.630 610.530 332.790 ;
        RECT 602.590 332.310 602.840 332.620 ;
        RECT 604.200 332.450 604.370 332.620 ;
        RECT 605.800 332.450 605.970 332.620 ;
        RECT 607.150 332.460 607.320 332.630 ;
        RECT 608.720 332.460 608.890 332.630 ;
        RECT 602.600 332.070 602.830 332.310 ;
        RECT 604.180 332.070 604.410 332.450 ;
        RECT 605.760 332.070 605.990 332.450 ;
        RECT 607.120 332.080 607.350 332.460 ;
        RECT 608.700 332.080 608.930 332.460 ;
        RECT 610.280 332.320 610.530 332.630 ;
        RECT 611.640 332.790 611.890 335.160 ;
        RECT 611.640 332.630 615.040 332.790 ;
        RECT 619.220 332.770 619.460 335.160 ;
        RECT 620.440 332.780 620.690 335.160 ;
        RECT 610.280 332.080 610.510 332.320 ;
        RECT 611.640 332.210 611.890 332.630 ;
        RECT 613.240 332.460 613.410 332.630 ;
        RECT 614.840 332.460 615.010 332.630 ;
        RECT 616.090 332.610 619.470 332.770 ;
        RECT 620.440 332.620 623.850 332.780 ;
        RECT 627.940 332.770 628.190 335.160 ;
        RECT 629.020 333.150 629.730 335.160 ;
        RECT 631.350 335.150 656.780 335.160 ;
        RECT 647.740 335.110 653.970 335.150 ;
        RECT 656.010 333.930 656.740 335.150 ;
        RECT 611.640 332.080 611.870 332.210 ;
        RECT 613.220 332.080 613.450 332.460 ;
        RECT 614.800 332.080 615.030 332.460 ;
        RECT 616.100 332.440 616.270 332.610 ;
        RECT 617.670 332.440 617.840 332.610 ;
        RECT 596.510 330.895 601.920 331.070 ;
        RECT 602.630 330.980 602.810 332.070 ;
        RECT 604.200 330.980 604.380 332.070 ;
        RECT 605.770 330.980 605.950 332.070 ;
        RECT 607.150 330.990 607.330 332.080 ;
        RECT 608.720 330.990 608.900 332.080 ;
        RECT 610.290 330.990 610.470 332.080 ;
        RECT 611.670 330.990 611.850 332.080 ;
        RECT 613.240 330.990 613.420 332.080 ;
        RECT 614.810 330.990 614.990 332.080 ;
        RECT 616.070 332.060 616.300 332.440 ;
        RECT 617.650 332.060 617.880 332.440 ;
        RECT 619.220 332.260 619.460 332.610 ;
        RECT 620.440 332.310 620.690 332.620 ;
        RECT 622.050 332.450 622.220 332.620 ;
        RECT 623.650 332.450 623.820 332.620 ;
        RECT 624.790 332.610 628.190 332.770 ;
        RECT 619.230 332.060 619.460 332.260 ;
        RECT 620.450 332.070 620.680 332.310 ;
        RECT 622.030 332.070 622.260 332.450 ;
        RECT 623.610 332.070 623.840 332.450 ;
        RECT 624.800 332.440 624.970 332.610 ;
        RECT 626.370 332.440 626.540 332.610 ;
        RECT 627.940 332.440 628.190 332.610 ;
        RECT 595.370 330.720 601.920 330.895 ;
        RECT 595.370 330.665 596.810 330.720 ;
        RECT 596.490 330.525 596.630 330.665 ;
        RECT 595.370 330.155 596.810 330.525 ;
        RECT 601.180 330.000 601.920 330.720 ;
        RECT 602.600 330.600 602.830 330.980 ;
        RECT 604.180 330.600 604.410 330.980 ;
        RECT 605.760 330.600 605.990 330.980 ;
        RECT 607.120 330.610 607.350 330.990 ;
        RECT 608.700 330.610 608.930 330.990 ;
        RECT 610.280 330.610 610.510 330.990 ;
        RECT 611.640 330.610 611.870 330.990 ;
        RECT 613.220 330.610 613.450 330.990 ;
        RECT 614.800 330.610 615.030 330.990 ;
        RECT 616.100 330.970 616.280 332.060 ;
        RECT 617.670 330.970 617.850 332.060 ;
        RECT 619.240 330.970 619.420 332.060 ;
        RECT 620.480 330.980 620.660 332.070 ;
        RECT 622.050 330.980 622.230 332.070 ;
        RECT 623.620 330.980 623.800 332.070 ;
        RECT 624.770 332.060 625.000 332.440 ;
        RECT 626.350 332.060 626.580 332.440 ;
        RECT 627.930 332.280 628.190 332.440 ;
        RECT 627.930 332.060 628.160 332.280 ;
        RECT 616.070 330.590 616.300 330.970 ;
        RECT 617.650 330.590 617.880 330.970 ;
        RECT 619.230 330.590 619.460 330.970 ;
        RECT 620.450 330.600 620.680 330.980 ;
        RECT 622.030 330.600 622.260 330.980 ;
        RECT 623.610 330.600 623.840 330.980 ;
        RECT 624.800 330.970 624.980 332.060 ;
        RECT 626.370 330.970 626.550 332.060 ;
        RECT 627.940 330.970 628.120 332.060 ;
        RECT 628.880 331.420 629.750 333.150 ;
        RECT 655.270 332.260 657.570 333.930 ;
        RECT 663.190 332.455 666.550 332.685 ;
        RECT 668.820 332.455 672.180 332.685 ;
        RECT 664.750 332.315 665.490 332.455 ;
        RECT 670.050 332.315 670.940 332.455 ;
        RECT 674.580 332.355 677.940 332.585 ;
        RECT 681.610 332.395 685.450 332.625 ;
        RECT 687.470 332.405 690.830 332.635 ;
        RECT 663.190 331.945 666.550 332.315 ;
        RECT 668.820 331.945 672.180 332.315 ;
        RECT 675.480 332.215 676.430 332.355 ;
        RECT 683.000 332.255 683.970 332.395 ;
        RECT 688.750 332.265 689.550 332.405 ;
        RECT 674.580 332.080 677.940 332.215 ;
        RECT 674.580 332.070 678.660 332.080 ;
        RECT 674.580 331.870 678.700 332.070 ;
        RECT 681.610 331.885 685.450 332.255 ;
        RECT 687.470 331.895 690.830 332.265 ;
        RECT 674.580 331.845 677.940 331.870 ;
        RECT 678.370 331.840 678.700 331.870 ;
        RECT 636.380 331.435 639.870 331.450 ;
        RECT 640.650 331.435 645.360 331.490 ;
        RECT 628.880 331.345 635.540 331.420 ;
        RECT 636.380 331.345 645.360 331.435 ;
        RECT 628.880 331.280 645.360 331.345 ;
        RECT 628.880 331.240 640.890 331.280 ;
        RECT 643.090 331.260 644.990 331.280 ;
        RECT 628.880 331.140 636.700 331.240 ;
        RECT 639.450 331.205 640.890 331.240 ;
        RECT 624.770 330.590 625.000 330.970 ;
        RECT 626.350 330.590 626.580 330.970 ;
        RECT 627.930 330.590 628.160 330.970 ;
        RECT 628.880 329.830 629.750 331.140 ;
        RECT 635.260 331.115 636.700 331.140 ;
        RECT 635.390 330.975 635.570 331.115 ;
        RECT 639.580 331.065 639.820 331.205 ;
        RECT 643.550 331.185 644.990 331.260 ;
        RECT 635.260 330.605 636.700 330.975 ;
        RECT 639.450 330.695 640.890 331.065 ;
        RECT 644.670 331.045 644.910 331.185 ;
        RECT 643.550 330.980 644.990 331.045 ;
        RECT 643.550 330.900 645.660 330.980 ;
        RECT 678.370 330.930 679.130 331.840 ;
        RECT 643.550 330.710 645.980 330.900 ;
        RECT 643.550 330.675 644.990 330.710 ;
        RECT 645.340 329.590 645.980 330.710 ;
        RECT 857.280 329.200 858.140 337.730 ;
        RECT 862.790 331.120 863.180 337.730 ;
        RECT 864.640 337.700 864.870 337.730 ;
        RECT 869.210 337.700 869.450 337.730 ;
        RECT 877.150 337.590 878.340 337.730 ;
        RECT 857.280 328.980 858.380 329.200 ;
        RECT 862.390 329.040 863.760 331.120 ;
        RECT 857.890 328.110 858.380 328.980 ;
        RECT 857.890 327.960 860.950 328.110 ;
        RECT 857.890 327.610 858.380 327.960 ;
        RECT 858.110 327.590 858.380 327.610 ;
        RECT 860.710 327.590 860.950 327.960 ;
        RECT 858.110 327.440 858.370 327.590 ;
        RECT 860.710 327.540 860.970 327.590 ;
        RECT 591.380 325.100 592.640 326.180 ;
        RECT 658.760 326.155 660.200 326.385 ;
        RECT 659.210 326.015 659.680 326.155 ;
        RECT 663.660 326.115 665.100 326.345 ;
        RECT 668.250 326.145 669.690 326.375 ;
        RECT 679.700 326.365 682.080 326.500 ;
        RECT 685.060 326.365 687.750 326.520 ;
        RECT 690.460 326.385 693.150 326.540 ;
        RECT 690.460 326.365 696.110 326.385 ;
        RECT 658.760 325.645 660.200 326.015 ;
        RECT 664.070 325.975 664.560 326.115 ;
        RECT 668.790 326.005 669.260 326.145 ;
        RECT 672.790 326.125 674.230 326.355 ;
        RECT 676.220 326.240 696.110 326.365 ;
        RECT 676.220 326.220 690.800 326.240 ;
        RECT 676.220 326.135 680.060 326.220 ;
        RECT 681.990 326.135 685.350 326.220 ;
        RECT 687.440 326.135 690.800 326.220 ;
        RECT 668.250 326.000 669.690 326.005 ;
        RECT 663.660 325.605 665.100 325.975 ;
        RECT 668.250 325.780 671.180 326.000 ;
        RECT 673.250 325.985 673.740 326.125 ;
        RECT 676.840 325.995 677.620 326.135 ;
        RECT 684.090 325.995 684.360 326.135 ;
        RECT 688.910 325.995 689.180 326.135 ;
        RECT 668.250 325.680 671.340 325.780 ;
        RECT 668.250 325.635 669.690 325.680 ;
        RECT 591.880 323.495 592.130 325.100 ;
        RECT 670.660 324.700 671.340 325.680 ;
        RECT 672.790 325.615 674.230 325.985 ;
        RECT 676.220 325.625 680.060 325.995 ;
        RECT 681.990 325.625 685.350 325.995 ;
        RECT 687.440 325.625 690.800 325.995 ;
        RECT 691.370 325.670 691.690 326.240 ;
        RECT 692.750 326.155 696.110 326.240 ;
        RECT 858.110 326.350 858.360 327.440 ;
        RECT 694.310 326.015 694.580 326.155 ;
        RECT 691.280 324.570 692.030 325.670 ;
        RECT 692.750 325.645 696.110 326.015 ;
        RECT 858.110 325.970 858.370 326.350 ;
        RECT 858.110 324.880 858.360 325.970 ;
        RECT 858.110 324.500 858.370 324.880 ;
        RECT 858.110 323.410 858.360 324.500 ;
        RECT 858.110 323.030 858.370 323.410 ;
        RECT 858.110 321.940 858.360 323.030 ;
        RECT 858.110 321.560 858.370 321.940 ;
        RECT 670.240 320.525 673.380 320.630 ;
        RECT 675.700 320.525 678.840 320.650 ;
        RECT 681.040 320.525 684.180 320.610 ;
        RECT 684.800 320.525 685.070 320.550 ;
        RECT 686.310 320.525 689.450 320.650 ;
        RECT 670.240 320.515 689.450 320.525 ;
        RECT 667.220 320.505 689.450 320.515 ;
        RECT 691.200 320.505 691.340 320.660 ;
        RECT 661.400 320.275 665.240 320.505 ;
        RECT 667.220 320.400 691.550 320.505 ;
        RECT 667.220 320.380 676.020 320.400 ;
        RECT 667.220 320.285 670.580 320.380 ;
        RECT 672.660 320.295 676.020 320.380 ;
        RECT 677.980 320.360 686.690 320.400 ;
        RECT 677.980 320.295 681.340 320.360 ;
        RECT 683.330 320.295 686.690 320.360 ;
        RECT 661.400 320.135 662.260 320.275 ;
        RECT 663.540 320.135 664.300 320.275 ;
        RECT 667.250 320.145 667.910 320.285 ;
        RECT 668.920 320.145 669.190 320.285 ;
        RECT 661.400 319.765 665.240 320.135 ;
        RECT 667.220 320.130 670.580 320.145 ;
        RECT 671.050 320.130 672.200 320.230 ;
        RECT 674.380 320.155 674.650 320.295 ;
        RECT 679.290 320.155 680.580 320.295 ;
        RECT 684.800 320.155 685.070 320.295 ;
        RECT 689.150 320.275 691.550 320.400 ;
        RECT 667.220 319.790 672.200 320.130 ;
        RECT 667.220 319.775 670.580 319.790 ;
        RECT 671.050 319.500 672.200 319.790 ;
        RECT 672.660 319.785 676.020 320.155 ;
        RECT 677.980 320.040 681.340 320.155 ;
        RECT 677.980 320.020 682.060 320.040 ;
        RECT 677.980 319.785 682.660 320.020 ;
        RECT 683.330 319.785 686.690 320.155 ;
        RECT 690.300 320.135 690.570 320.275 ;
        RECT 689.150 320.130 691.550 320.135 ;
        RECT 691.930 320.130 693.110 320.460 ;
        RECT 693.550 320.275 695.950 320.505 ;
        RECT 858.110 320.470 858.360 321.560 ;
        RECT 860.720 320.520 860.970 327.540 ;
        RECT 864.660 321.160 867.480 321.190 ;
        RECT 868.600 321.160 871.420 321.180 ;
        RECT 864.660 321.150 871.420 321.160 ;
        RECT 871.900 321.150 872.230 321.300 ;
        RECT 864.660 321.000 872.230 321.150 ;
        RECT 864.680 320.850 864.920 321.000 ;
        RECT 867.200 320.990 872.230 321.000 ;
        RECT 867.200 320.950 868.970 320.990 ;
        RECT 867.280 320.930 868.970 320.950 ;
        RECT 864.680 320.710 864.940 320.850 ;
        RECT 867.280 320.750 867.520 320.930 ;
        RECT 864.680 320.590 864.960 320.710 ;
        RECT 867.280 320.590 867.570 320.750 ;
        RECT 694.750 320.135 695.020 320.275 ;
        RECT 681.260 319.750 682.660 319.785 ;
        RECT 689.150 319.780 693.110 320.130 ;
        RECT 689.150 319.765 691.550 319.780 ;
        RECT 681.830 319.140 682.660 319.750 ;
        RECT 691.930 319.730 693.110 319.780 ;
        RECT 693.550 319.765 695.950 320.135 ;
        RECT 858.110 320.090 858.370 320.470 ;
        RECT 858.110 319.000 858.360 320.090 ;
        RECT 860.610 319.780 861.190 320.520 ;
        RECT 864.620 319.920 865.060 320.590 ;
        RECT 867.290 320.470 867.570 320.590 ;
        RECT 868.620 320.660 868.970 320.930 ;
        RECT 871.220 320.740 871.460 320.990 ;
        RECT 871.760 320.840 872.230 320.990 ;
        RECT 868.620 320.580 868.900 320.660 ;
        RECT 871.220 320.580 871.510 320.740 ;
        RECT 858.110 318.620 858.370 319.000 ;
        RECT 590.390 317.750 591.490 318.050 ;
        RECT 600.350 317.750 631.840 317.810 ;
        RECT 590.390 317.030 631.840 317.750 ;
        RECT 590.390 316.840 591.490 317.030 ;
        RECT 600.350 316.990 631.840 317.030 ;
        RECT 858.110 317.530 858.360 318.620 ;
        RECT 858.110 317.150 858.370 317.530 ;
        RECT 601.030 314.690 601.740 316.990 ;
        RECT 601.030 312.900 601.770 314.690 ;
        RECT 602.440 314.610 602.690 316.990 ;
        RECT 610.130 314.620 610.380 316.990 ;
        RECT 602.440 314.450 605.850 314.610 ;
        RECT 606.990 314.460 610.380 314.620 ;
        RECT 602.440 314.140 602.690 314.450 ;
        RECT 604.050 314.280 604.220 314.450 ;
        RECT 605.650 314.280 605.820 314.450 ;
        RECT 607.000 314.290 607.170 314.460 ;
        RECT 608.570 314.290 608.740 314.460 ;
        RECT 602.450 313.900 602.680 314.140 ;
        RECT 604.030 313.900 604.260 314.280 ;
        RECT 605.610 313.900 605.840 314.280 ;
        RECT 606.970 313.910 607.200 314.290 ;
        RECT 608.550 313.910 608.780 314.290 ;
        RECT 610.130 314.150 610.380 314.460 ;
        RECT 611.490 314.620 611.740 316.990 ;
        RECT 611.490 314.460 614.890 314.620 ;
        RECT 619.070 314.600 619.310 316.990 ;
        RECT 620.290 314.610 620.540 316.990 ;
        RECT 610.130 313.910 610.360 314.150 ;
        RECT 611.490 314.040 611.740 314.460 ;
        RECT 613.090 314.290 613.260 314.460 ;
        RECT 614.690 314.290 614.860 314.460 ;
        RECT 615.940 314.440 619.320 314.600 ;
        RECT 620.290 314.450 623.700 314.610 ;
        RECT 627.790 314.600 628.040 316.990 ;
        RECT 628.870 314.980 629.580 316.990 ;
        RECT 858.110 316.060 858.360 317.150 ;
        RECT 858.110 315.680 858.370 316.060 ;
        RECT 611.490 313.910 611.720 314.040 ;
        RECT 613.070 313.910 613.300 314.290 ;
        RECT 614.650 313.910 614.880 314.290 ;
        RECT 615.950 314.270 616.120 314.440 ;
        RECT 617.520 314.270 617.690 314.440 ;
        RECT 596.360 312.725 601.770 312.900 ;
        RECT 602.480 312.810 602.660 313.900 ;
        RECT 604.050 312.810 604.230 313.900 ;
        RECT 605.620 312.810 605.800 313.900 ;
        RECT 607.000 312.820 607.180 313.910 ;
        RECT 608.570 312.820 608.750 313.910 ;
        RECT 610.140 312.820 610.320 313.910 ;
        RECT 611.520 312.820 611.700 313.910 ;
        RECT 613.090 312.820 613.270 313.910 ;
        RECT 614.660 312.820 614.840 313.910 ;
        RECT 615.920 313.890 616.150 314.270 ;
        RECT 617.500 313.890 617.730 314.270 ;
        RECT 619.070 314.090 619.310 314.440 ;
        RECT 620.290 314.140 620.540 314.450 ;
        RECT 621.900 314.280 622.070 314.450 ;
        RECT 623.500 314.280 623.670 314.450 ;
        RECT 624.640 314.440 628.040 314.600 ;
        RECT 619.080 313.890 619.310 314.090 ;
        RECT 620.300 313.900 620.530 314.140 ;
        RECT 621.880 313.900 622.110 314.280 ;
        RECT 623.460 313.900 623.690 314.280 ;
        RECT 624.650 314.270 624.820 314.440 ;
        RECT 626.220 314.270 626.390 314.440 ;
        RECT 627.790 314.270 628.040 314.440 ;
        RECT 595.220 312.550 601.770 312.725 ;
        RECT 595.220 312.495 596.660 312.550 ;
        RECT 596.340 312.355 596.480 312.495 ;
        RECT 595.220 311.985 596.660 312.355 ;
        RECT 601.030 311.830 601.770 312.550 ;
        RECT 602.450 312.430 602.680 312.810 ;
        RECT 604.030 312.430 604.260 312.810 ;
        RECT 605.610 312.430 605.840 312.810 ;
        RECT 606.970 312.440 607.200 312.820 ;
        RECT 608.550 312.440 608.780 312.820 ;
        RECT 610.130 312.440 610.360 312.820 ;
        RECT 611.490 312.440 611.720 312.820 ;
        RECT 613.070 312.440 613.300 312.820 ;
        RECT 614.650 312.440 614.880 312.820 ;
        RECT 615.950 312.800 616.130 313.890 ;
        RECT 617.520 312.800 617.700 313.890 ;
        RECT 619.090 312.800 619.270 313.890 ;
        RECT 620.330 312.810 620.510 313.900 ;
        RECT 621.900 312.810 622.080 313.900 ;
        RECT 623.470 312.810 623.650 313.900 ;
        RECT 624.620 313.890 624.850 314.270 ;
        RECT 626.200 313.890 626.430 314.270 ;
        RECT 627.780 314.110 628.040 314.270 ;
        RECT 627.780 313.890 628.010 314.110 ;
        RECT 615.920 312.420 616.150 312.800 ;
        RECT 617.500 312.420 617.730 312.800 ;
        RECT 619.080 312.420 619.310 312.800 ;
        RECT 620.300 312.430 620.530 312.810 ;
        RECT 621.880 312.430 622.110 312.810 ;
        RECT 623.460 312.430 623.690 312.810 ;
        RECT 624.650 312.800 624.830 313.890 ;
        RECT 626.220 312.800 626.400 313.890 ;
        RECT 627.790 312.800 627.970 313.890 ;
        RECT 628.730 313.250 629.600 314.980 ;
        RECT 680.050 314.580 680.720 315.030 ;
        RECT 858.110 314.590 858.360 315.680 ;
        RECT 636.230 313.265 639.720 313.280 ;
        RECT 640.500 313.265 645.210 313.320 ;
        RECT 628.730 313.175 635.390 313.250 ;
        RECT 636.230 313.175 645.210 313.265 ;
        RECT 628.730 313.110 645.210 313.175 ;
        RECT 628.730 313.070 640.740 313.110 ;
        RECT 642.940 313.090 644.840 313.110 ;
        RECT 628.730 312.970 636.550 313.070 ;
        RECT 639.300 313.035 640.740 313.070 ;
        RECT 624.620 312.420 624.850 312.800 ;
        RECT 626.200 312.420 626.430 312.800 ;
        RECT 627.780 312.420 628.010 312.800 ;
        RECT 628.730 311.660 629.600 312.970 ;
        RECT 635.110 312.945 636.550 312.970 ;
        RECT 635.240 312.805 635.420 312.945 ;
        RECT 639.430 312.895 639.670 313.035 ;
        RECT 643.400 313.015 644.840 313.090 ;
        RECT 635.110 312.435 636.550 312.805 ;
        RECT 639.300 312.525 640.740 312.895 ;
        RECT 644.520 312.875 644.760 313.015 ;
        RECT 643.400 312.820 644.840 312.875 ;
        RECT 645.240 312.820 645.880 312.920 ;
        RECT 643.400 312.550 645.880 312.820 ;
        RECT 643.400 312.505 644.840 312.550 ;
        RECT 645.240 311.610 645.880 312.550 ;
        RECT 680.290 303.370 680.480 314.580 ;
        RECT 858.110 314.330 858.370 314.590 ;
        RECT 858.140 314.210 858.370 314.330 ;
        RECT 860.720 314.310 860.970 319.780 ;
        RECT 864.690 314.750 864.960 319.920 ;
        RECT 867.300 319.380 867.570 320.470 ;
        RECT 867.290 319.000 867.570 319.380 ;
        RECT 867.300 317.910 867.570 319.000 ;
        RECT 867.290 317.530 867.570 317.910 ;
        RECT 867.300 316.440 867.570 317.530 ;
        RECT 867.290 316.060 867.570 316.440 ;
        RECT 867.300 314.970 867.570 316.060 ;
        RECT 867.290 314.790 867.570 314.970 ;
        RECT 864.710 314.590 864.940 314.750 ;
        RECT 867.290 314.590 867.520 314.790 ;
        RECT 868.630 314.740 868.900 320.580 ;
        RECT 871.230 320.460 871.510 320.580 ;
        RECT 871.240 319.370 871.510 320.460 ;
        RECT 871.230 318.990 871.510 319.370 ;
        RECT 871.900 319.010 872.230 320.840 ;
        RECT 871.240 317.900 871.510 318.990 ;
        RECT 871.230 317.520 871.510 317.900 ;
        RECT 871.240 316.430 871.510 317.520 ;
        RECT 871.230 316.050 871.510 316.430 ;
        RECT 871.240 314.960 871.510 316.050 ;
        RECT 871.830 315.090 872.310 319.010 ;
        RECT 871.230 314.780 871.510 314.960 ;
        RECT 868.650 314.580 868.880 314.740 ;
        RECT 871.230 314.580 871.460 314.780 ;
        RECT 860.720 314.210 860.950 314.310 ;
        RECT 796.480 308.170 811.840 308.215 ;
        RECT 814.240 308.170 829.600 308.215 ;
        RECT 831.780 308.170 833.220 308.185 ;
        RECT 796.480 308.150 833.220 308.170 ;
        RECT 835.420 308.180 840.700 308.245 ;
        RECT 842.690 308.180 844.130 308.245 ;
        RECT 835.420 308.150 844.130 308.180 ;
        RECT 796.480 308.120 844.130 308.150 ;
        RECT 854.330 308.120 856.310 308.140 ;
        RECT 796.480 308.015 856.310 308.120 ;
        RECT 796.480 307.985 836.410 308.015 ;
        RECT 810.950 307.845 814.710 307.985 ;
        RECT 828.660 307.875 836.410 307.985 ;
        RECT 840.370 307.875 856.310 308.015 ;
        RECT 828.660 307.845 856.310 307.875 ;
        RECT 796.480 307.720 856.310 307.845 ;
        RECT 796.480 307.650 840.700 307.720 ;
        RECT 796.480 307.475 811.840 307.650 ;
        RECT 812.180 307.320 813.390 307.650 ;
        RECT 814.240 307.475 829.600 307.650 ;
        RECT 830.070 307.320 831.280 307.650 ;
        RECT 831.780 307.630 840.700 307.650 ;
        RECT 831.780 307.445 833.220 307.630 ;
        RECT 835.420 307.505 840.700 307.630 ;
        RECT 841.170 307.300 842.380 307.720 ;
        RECT 842.690 307.650 856.310 307.720 ;
        RECT 842.690 307.505 844.130 307.650 ;
        RECT 854.330 307.610 856.310 307.650 ;
        RECT 680.260 302.100 680.510 303.370 ;
        RECT 680.290 299.700 680.480 302.100 ;
        RECT 679.810 299.155 680.760 299.700 ;
        RECT 679.810 299.100 695.420 299.155 ;
        RECT 715.160 299.140 730.520 299.175 ;
        RECT 711.410 299.115 730.520 299.140 ;
        RECT 680.060 299.070 695.420 299.100 ;
        RECT 697.550 299.080 730.520 299.115 ;
        RECT 732.860 299.080 748.220 299.125 ;
        RECT 750.600 299.080 765.960 299.115 ;
        RECT 697.550 299.070 765.960 299.080 ;
        RECT 680.060 298.945 765.960 299.070 ;
        RECT 680.060 298.925 715.660 298.945 ;
        RECT 590.490 298.580 591.590 298.890 ;
        RECT 680.290 298.785 680.480 298.925 ;
        RECT 694.250 298.885 715.660 298.925 ;
        RECT 694.250 298.785 698.500 298.885 ;
        RECT 680.060 298.745 698.500 298.785 ;
        RECT 711.410 298.805 715.660 298.885 ;
        RECT 729.390 298.895 765.960 298.945 ;
        RECT 729.390 298.805 733.640 298.895 ;
        RECT 711.410 298.755 733.640 298.805 ;
        RECT 747.120 298.885 765.960 298.895 ;
        RECT 747.120 298.755 751.370 298.885 ;
        RECT 711.410 298.745 751.370 298.755 ;
        RECT 600.300 298.580 631.790 298.630 ;
        RECT 590.490 297.860 631.790 298.580 ;
        RECT 680.060 298.620 765.960 298.745 ;
        RECT 680.060 298.550 712.910 298.620 ;
        RECT 680.060 298.415 695.420 298.550 ;
        RECT 695.850 297.880 696.860 298.550 ;
        RECT 697.550 298.375 712.910 298.550 ;
        RECT 713.500 298.240 714.440 298.620 ;
        RECT 715.160 298.560 765.960 298.620 ;
        RECT 715.160 298.435 730.520 298.560 ;
        RECT 731.130 298.080 732.050 298.560 ;
        RECT 732.860 298.385 748.220 298.560 ;
        RECT 748.900 298.060 749.740 298.560 ;
        RECT 750.600 298.375 765.960 298.560 ;
        RECT 855.880 298.475 856.300 307.610 ;
        RECT 855.800 298.245 859.160 298.475 ;
        RECT 855.880 298.105 856.300 298.245 ;
        RECT 858.260 298.105 858.690 298.245 ;
        RECT 855.800 298.060 859.160 298.105 ;
        RECT 859.720 298.060 860.310 298.420 ;
        RECT 590.490 297.680 591.590 297.860 ;
        RECT 600.300 297.810 631.790 297.860 ;
        RECT 855.800 297.840 860.310 298.060 ;
        RECT 600.980 295.510 601.690 297.810 ;
        RECT 600.980 293.720 601.720 295.510 ;
        RECT 602.390 295.430 602.640 297.810 ;
        RECT 610.080 295.440 610.330 297.810 ;
        RECT 602.390 295.270 605.800 295.430 ;
        RECT 606.940 295.280 610.330 295.440 ;
        RECT 602.390 294.960 602.640 295.270 ;
        RECT 604.000 295.100 604.170 295.270 ;
        RECT 605.600 295.100 605.770 295.270 ;
        RECT 606.950 295.110 607.120 295.280 ;
        RECT 608.520 295.110 608.690 295.280 ;
        RECT 602.400 294.720 602.630 294.960 ;
        RECT 603.980 294.720 604.210 295.100 ;
        RECT 605.560 294.720 605.790 295.100 ;
        RECT 606.920 294.730 607.150 295.110 ;
        RECT 608.500 294.730 608.730 295.110 ;
        RECT 610.080 294.970 610.330 295.280 ;
        RECT 611.440 295.440 611.690 297.810 ;
        RECT 611.440 295.280 614.840 295.440 ;
        RECT 619.020 295.420 619.260 297.810 ;
        RECT 620.240 295.430 620.490 297.810 ;
        RECT 610.080 294.730 610.310 294.970 ;
        RECT 611.440 294.860 611.690 295.280 ;
        RECT 613.040 295.110 613.210 295.280 ;
        RECT 614.640 295.110 614.810 295.280 ;
        RECT 615.890 295.260 619.270 295.420 ;
        RECT 620.240 295.270 623.650 295.430 ;
        RECT 627.740 295.420 627.990 297.810 ;
        RECT 628.820 295.800 629.530 297.810 ;
        RECT 855.800 297.735 859.160 297.840 ;
        RECT 859.720 297.680 860.310 297.840 ;
        RECT 834.860 296.520 839.720 296.540 ;
        RECT 844.890 296.530 845.320 296.540 ;
        RECT 834.840 296.495 839.720 296.520 ;
        RECT 842.500 296.495 845.320 296.530 ;
        RECT 834.840 296.370 845.320 296.495 ;
        RECT 611.440 294.730 611.670 294.860 ;
        RECT 613.020 294.730 613.250 295.110 ;
        RECT 614.600 294.730 614.830 295.110 ;
        RECT 615.900 295.090 616.070 295.260 ;
        RECT 617.470 295.090 617.640 295.260 ;
        RECT 596.310 293.545 601.720 293.720 ;
        RECT 602.430 293.630 602.610 294.720 ;
        RECT 604.000 293.630 604.180 294.720 ;
        RECT 605.570 293.630 605.750 294.720 ;
        RECT 606.950 293.640 607.130 294.730 ;
        RECT 608.520 293.640 608.700 294.730 ;
        RECT 610.090 293.640 610.270 294.730 ;
        RECT 611.470 293.640 611.650 294.730 ;
        RECT 613.040 293.640 613.220 294.730 ;
        RECT 614.610 293.640 614.790 294.730 ;
        RECT 615.870 294.710 616.100 295.090 ;
        RECT 617.450 294.710 617.680 295.090 ;
        RECT 619.020 294.910 619.260 295.260 ;
        RECT 620.240 294.960 620.490 295.270 ;
        RECT 621.850 295.100 622.020 295.270 ;
        RECT 623.450 295.100 623.620 295.270 ;
        RECT 624.590 295.260 627.990 295.420 ;
        RECT 619.030 294.710 619.260 294.910 ;
        RECT 620.250 294.720 620.480 294.960 ;
        RECT 621.830 294.720 622.060 295.100 ;
        RECT 623.410 294.720 623.640 295.100 ;
        RECT 624.600 295.090 624.770 295.260 ;
        RECT 626.170 295.090 626.340 295.260 ;
        RECT 627.740 295.090 627.990 295.260 ;
        RECT 595.170 293.370 601.720 293.545 ;
        RECT 595.170 293.315 596.610 293.370 ;
        RECT 596.290 293.175 596.430 293.315 ;
        RECT 595.170 292.805 596.610 293.175 ;
        RECT 600.980 292.650 601.720 293.370 ;
        RECT 602.400 293.250 602.630 293.630 ;
        RECT 603.980 293.250 604.210 293.630 ;
        RECT 605.560 293.250 605.790 293.630 ;
        RECT 606.920 293.260 607.150 293.640 ;
        RECT 608.500 293.260 608.730 293.640 ;
        RECT 610.080 293.260 610.310 293.640 ;
        RECT 611.440 293.260 611.670 293.640 ;
        RECT 613.020 293.260 613.250 293.640 ;
        RECT 614.600 293.260 614.830 293.640 ;
        RECT 615.900 293.620 616.080 294.710 ;
        RECT 617.470 293.620 617.650 294.710 ;
        RECT 619.040 293.620 619.220 294.710 ;
        RECT 620.280 293.630 620.460 294.720 ;
        RECT 621.850 293.630 622.030 294.720 ;
        RECT 623.420 293.630 623.600 294.720 ;
        RECT 624.570 294.710 624.800 295.090 ;
        RECT 626.150 294.710 626.380 295.090 ;
        RECT 627.730 294.930 627.990 295.090 ;
        RECT 627.730 294.710 627.960 294.930 ;
        RECT 615.870 293.240 616.100 293.620 ;
        RECT 617.450 293.240 617.680 293.620 ;
        RECT 619.030 293.240 619.260 293.620 ;
        RECT 620.250 293.250 620.480 293.630 ;
        RECT 621.830 293.250 622.060 293.630 ;
        RECT 623.410 293.250 623.640 293.630 ;
        RECT 624.600 293.620 624.780 294.710 ;
        RECT 626.170 293.620 626.350 294.710 ;
        RECT 627.740 293.620 627.920 294.710 ;
        RECT 628.680 294.070 629.550 295.800 ;
        RECT 636.180 294.085 639.670 294.100 ;
        RECT 640.450 294.085 645.160 294.140 ;
        RECT 628.680 293.995 635.340 294.070 ;
        RECT 636.180 293.995 645.160 294.085 ;
        RECT 628.680 293.930 645.160 293.995 ;
        RECT 628.680 293.890 640.690 293.930 ;
        RECT 642.890 293.910 644.790 293.930 ;
        RECT 628.680 293.790 636.500 293.890 ;
        RECT 639.250 293.855 640.690 293.890 ;
        RECT 624.570 293.240 624.800 293.620 ;
        RECT 626.150 293.240 626.380 293.620 ;
        RECT 627.730 293.240 627.960 293.620 ;
        RECT 628.680 292.480 629.550 293.790 ;
        RECT 635.060 293.765 636.500 293.790 ;
        RECT 635.190 293.625 635.370 293.765 ;
        RECT 639.380 293.715 639.620 293.855 ;
        RECT 643.350 293.835 644.790 293.910 ;
        RECT 635.060 293.255 636.500 293.625 ;
        RECT 639.250 293.345 640.690 293.715 ;
        RECT 644.470 293.695 644.710 293.835 ;
        RECT 643.350 293.650 644.790 293.695 ;
        RECT 643.350 293.380 645.950 293.650 ;
        RECT 643.350 293.325 644.790 293.380 ;
        RECT 645.310 292.340 645.950 293.380 ;
        RECT 818.940 293.255 822.300 293.485 ;
        RECT 820.430 293.115 820.650 293.255 ;
        RECT 818.940 293.010 822.300 293.115 ;
        RECT 818.940 292.760 824.550 293.010 ;
        RECT 818.940 292.745 822.300 292.760 ;
        RECT 819.460 292.510 819.860 292.745 ;
        RECT 822.770 292.210 823.750 292.760 ;
        RECT 824.370 291.315 824.550 292.760 ;
        RECT 827.430 291.335 830.270 291.370 ;
        RECT 834.840 291.335 835.100 296.370 ;
        RECT 839.390 296.360 845.310 296.370 ;
        RECT 839.390 296.265 842.750 296.360 ;
        RECT 841.470 296.125 841.690 296.265 ;
        RECT 839.390 295.755 842.750 296.125 ;
        RECT 843.310 295.390 844.180 296.360 ;
        RECT 844.870 296.200 845.310 296.360 ;
        RECT 845.150 294.845 845.310 296.200 ;
        RECT 846.750 294.845 846.970 294.850 ;
        RECT 845.090 294.615 848.450 294.845 ;
        RECT 846.750 294.475 846.970 294.615 ;
        RECT 845.090 294.105 848.450 294.475 ;
        RECT 861.180 294.345 864.540 294.575 ;
        RECT 862.170 294.205 862.390 294.345 ;
        RECT 863.680 294.205 864.140 294.345 ;
        RECT 861.180 293.835 864.540 294.205 ;
        RECT 858.330 292.945 858.760 293.250 ;
        RECT 855.840 292.715 859.200 292.945 ;
        RECT 858.060 292.575 858.280 292.715 ;
        RECT 855.840 292.205 859.200 292.575 ;
        RECT 827.430 291.315 835.210 291.335 ;
        RECT 824.370 291.200 835.210 291.315 ;
        RECT 824.370 291.110 827.750 291.200 ;
        RECT 824.390 291.085 827.750 291.110 ;
        RECT 825.780 290.945 826.000 291.085 ;
        RECT 824.390 290.575 827.750 290.945 ;
        RECT 828.220 290.410 828.930 291.200 ;
        RECT 829.930 291.105 835.210 291.200 ;
        RECT 839.400 291.145 842.760 291.375 ;
        RECT 831.650 290.965 831.870 291.105 ;
        RECT 833.280 290.965 833.500 291.105 ;
        RECT 841.190 291.005 841.810 291.145 ;
        RECT 829.930 290.595 835.210 290.965 ;
        RECT 839.400 290.635 842.760 291.005 ;
        RECT 819.400 288.325 819.850 288.610 ;
        RECT 818.910 288.095 822.270 288.325 ;
        RECT 820.430 287.955 820.650 288.095 ;
        RECT 818.910 287.585 822.270 287.955 ;
        RECT 858.350 287.545 858.910 288.010 ;
        RECT 855.910 287.315 859.270 287.545 ;
        RECT 856.080 287.175 856.780 287.315 ;
        RECT 857.970 287.175 858.190 287.315 ;
        RECT 855.910 286.805 859.270 287.175 ;
        RECT 860.060 285.720 860.940 286.160 ;
        RECT 860.060 285.525 861.590 285.720 ;
        RECT 860.060 285.340 864.620 285.525 ;
        RECT 860.060 285.200 860.940 285.340 ;
        RECT 861.260 285.295 864.620 285.340 ;
        RECT 862.910 285.155 864.170 285.295 ;
        RECT 861.260 284.785 864.620 285.155 ;
        RECT 799.530 283.405 800.970 283.635 ;
        RECT 800.040 283.265 800.550 283.405 ;
        RECT 819.490 283.295 819.890 283.680 ;
        RECT 799.530 282.895 800.970 283.265 ;
        RECT 819.350 283.065 824.630 283.295 ;
        RECT 828.120 283.205 828.620 283.660 ;
        RECT 831.110 283.205 833.320 283.290 ;
        RECT 838.220 283.205 840.710 283.230 ;
        RECT 841.830 283.205 842.270 283.490 ;
        RECT 843.990 283.205 846.580 283.220 ;
        RECT 827.960 283.070 851.580 283.205 ;
        RECT 821.720 282.925 822.030 283.065 ;
        RECT 827.960 282.975 831.320 283.070 ;
        RECT 684.390 282.425 696.960 282.640 ;
        RECT 710.120 282.590 710.720 282.600 ;
        RECT 701.660 282.425 714.860 282.590 ;
        RECT 719.380 282.425 732.580 282.570 ;
        RECT 736.600 282.435 749.800 282.570 ;
        RECT 819.350 282.555 824.630 282.925 ;
        RECT 829.540 282.835 829.850 282.975 ;
        RECT 827.960 282.465 831.320 282.835 ;
        RECT 736.600 282.425 754.440 282.435 ;
        RECT 684.390 282.415 754.440 282.425 ;
        RECT 679.390 282.300 754.440 282.415 ;
        RECT 679.390 282.280 701.950 282.300 ;
        RECT 679.390 282.270 690.240 282.280 ;
        RECT 690.800 282.270 701.950 282.280 ;
        RECT 679.390 282.185 684.670 282.270 ;
        RECT 679.760 282.045 680.400 282.185 ;
        RECT 681.680 282.045 681.860 282.185 ;
        RECT 679.390 281.675 684.670 282.045 ;
        RECT 685.190 281.630 685.940 282.270 ;
        RECT 589.960 280.120 591.060 280.350 ;
        RECT 682.190 280.320 682.640 280.380 ;
        RECT 690.810 280.320 691.120 282.270 ;
        RECT 696.670 282.195 701.950 282.270 ;
        RECT 698.290 282.055 698.470 282.195 ;
        RECT 699.840 282.055 700.140 282.195 ;
        RECT 696.670 281.685 701.950 282.055 ;
        RECT 702.800 281.400 703.490 282.300 ;
        RECT 710.120 281.890 710.720 282.300 ;
        RECT 714.440 282.280 754.440 282.300 ;
        RECT 714.440 282.195 719.720 282.280 ;
        RECT 717.230 282.055 717.530 282.195 ;
        RECT 714.440 281.685 719.720 282.055 ;
        RECT 720.220 281.450 721.180 282.280 ;
        RECT 731.680 282.195 736.960 282.280 ;
        RECT 734.170 282.055 734.430 282.195 ;
        RECT 731.680 281.685 736.960 282.055 ;
        RECT 737.630 281.300 738.670 282.280 ;
        RECT 749.160 282.205 754.440 282.280 ;
        RECT 752.140 282.065 753.660 282.205 ;
        RECT 749.160 282.020 754.440 282.065 ;
        RECT 754.830 282.020 755.580 282.390 ;
        RECT 831.640 282.250 832.740 283.070 ;
        RECT 833.250 282.975 838.530 283.070 ;
        RECT 835.660 282.835 835.970 282.975 ;
        RECT 833.250 282.465 838.530 282.835 ;
        RECT 838.950 282.390 839.860 283.070 ;
        RECT 840.460 283.050 851.580 283.070 ;
        RECT 840.460 282.975 844.300 283.050 ;
        RECT 846.300 282.975 851.580 283.050 ;
        RECT 842.920 282.835 843.650 282.975 ;
        RECT 850.520 282.835 850.680 282.975 ;
        RECT 840.460 282.465 844.300 282.835 ;
        RECT 846.300 282.810 851.580 282.835 ;
        RECT 851.880 282.810 852.500 283.150 ;
        RECT 846.300 282.600 852.500 282.810 ;
        RECT 846.300 282.465 851.580 282.600 ;
        RECT 851.880 282.530 852.500 282.600 ;
        RECT 858.350 282.085 858.910 282.600 ;
        RECT 749.160 281.790 755.580 282.020 ;
        RECT 855.930 281.855 859.290 282.085 ;
        RECT 749.160 281.695 754.440 281.790 ;
        RECT 754.830 281.640 755.580 281.790 ;
        RECT 857.410 281.715 857.630 281.855 ;
        RECT 855.930 281.345 859.290 281.715 ;
        RECT 699.490 280.320 699.940 280.430 ;
        RECT 717.280 280.320 717.730 280.470 ;
        RECT 734.540 280.320 734.990 280.500 ;
        RECT 752.010 280.410 752.460 280.490 ;
        RECT 756.350 280.410 757.010 280.560 ;
        RECT 752.010 280.320 757.010 280.410 ;
        RECT 682.190 280.230 757.010 280.320 ;
        RECT 682.190 280.180 752.460 280.230 ;
        RECT 600.220 280.120 631.710 280.160 ;
        RECT 589.960 279.400 631.710 280.120 ;
        RECT 682.190 280.040 682.640 280.180 ;
        RECT 699.490 280.090 699.940 280.180 ;
        RECT 717.280 280.130 717.730 280.180 ;
        RECT 734.540 280.160 734.990 280.180 ;
        RECT 752.010 280.150 752.460 280.180 ;
        RECT 756.350 279.950 757.010 280.230 ;
        RECT 589.960 279.140 591.060 279.400 ;
        RECT 600.220 279.340 631.710 279.400 ;
        RECT 600.900 277.040 601.610 279.340 ;
        RECT 600.900 275.250 601.640 277.040 ;
        RECT 602.310 276.960 602.560 279.340 ;
        RECT 610.000 276.970 610.250 279.340 ;
        RECT 602.310 276.800 605.720 276.960 ;
        RECT 606.860 276.810 610.250 276.970 ;
        RECT 602.310 276.490 602.560 276.800 ;
        RECT 603.920 276.630 604.090 276.800 ;
        RECT 605.520 276.630 605.690 276.800 ;
        RECT 606.870 276.640 607.040 276.810 ;
        RECT 608.440 276.640 608.610 276.810 ;
        RECT 602.320 276.250 602.550 276.490 ;
        RECT 603.900 276.250 604.130 276.630 ;
        RECT 605.480 276.250 605.710 276.630 ;
        RECT 606.840 276.260 607.070 276.640 ;
        RECT 608.420 276.260 608.650 276.640 ;
        RECT 610.000 276.500 610.250 276.810 ;
        RECT 611.360 276.970 611.610 279.340 ;
        RECT 611.360 276.810 614.760 276.970 ;
        RECT 618.940 276.950 619.180 279.340 ;
        RECT 620.160 276.960 620.410 279.340 ;
        RECT 610.000 276.260 610.230 276.500 ;
        RECT 611.360 276.390 611.610 276.810 ;
        RECT 612.960 276.640 613.130 276.810 ;
        RECT 614.560 276.640 614.730 276.810 ;
        RECT 615.810 276.790 619.190 276.950 ;
        RECT 620.160 276.800 623.570 276.960 ;
        RECT 627.660 276.950 627.910 279.340 ;
        RECT 628.740 277.330 629.450 279.340 ;
        RECT 611.360 276.260 611.590 276.390 ;
        RECT 612.940 276.260 613.170 276.640 ;
        RECT 614.520 276.260 614.750 276.640 ;
        RECT 615.820 276.620 615.990 276.790 ;
        RECT 617.390 276.620 617.560 276.790 ;
        RECT 596.230 275.075 601.640 275.250 ;
        RECT 602.350 275.160 602.530 276.250 ;
        RECT 603.920 275.160 604.100 276.250 ;
        RECT 605.490 275.160 605.670 276.250 ;
        RECT 606.870 275.170 607.050 276.260 ;
        RECT 608.440 275.170 608.620 276.260 ;
        RECT 610.010 275.170 610.190 276.260 ;
        RECT 611.390 275.170 611.570 276.260 ;
        RECT 612.960 275.170 613.140 276.260 ;
        RECT 614.530 275.170 614.710 276.260 ;
        RECT 615.790 276.240 616.020 276.620 ;
        RECT 617.370 276.240 617.600 276.620 ;
        RECT 618.940 276.440 619.180 276.790 ;
        RECT 620.160 276.490 620.410 276.800 ;
        RECT 621.770 276.630 621.940 276.800 ;
        RECT 623.370 276.630 623.540 276.800 ;
        RECT 624.510 276.790 627.910 276.950 ;
        RECT 618.950 276.240 619.180 276.440 ;
        RECT 620.170 276.250 620.400 276.490 ;
        RECT 621.750 276.250 621.980 276.630 ;
        RECT 623.330 276.250 623.560 276.630 ;
        RECT 624.520 276.620 624.690 276.790 ;
        RECT 626.090 276.620 626.260 276.790 ;
        RECT 627.660 276.620 627.910 276.790 ;
        RECT 595.090 274.900 601.640 275.075 ;
        RECT 595.090 274.845 596.530 274.900 ;
        RECT 409.470 274.730 410.430 274.770 ;
        RECT 409.470 274.590 410.640 274.730 ;
        RECT 596.210 274.705 596.350 274.845 ;
        RECT 409.480 271.470 410.640 274.590 ;
        RECT 595.090 274.335 596.530 274.705 ;
        RECT 600.900 274.180 601.640 274.900 ;
        RECT 602.320 274.780 602.550 275.160 ;
        RECT 603.900 274.780 604.130 275.160 ;
        RECT 605.480 274.780 605.710 275.160 ;
        RECT 606.840 274.790 607.070 275.170 ;
        RECT 608.420 274.790 608.650 275.170 ;
        RECT 610.000 274.790 610.230 275.170 ;
        RECT 611.360 274.790 611.590 275.170 ;
        RECT 612.940 274.790 613.170 275.170 ;
        RECT 614.520 274.790 614.750 275.170 ;
        RECT 615.820 275.150 616.000 276.240 ;
        RECT 617.390 275.150 617.570 276.240 ;
        RECT 618.960 275.150 619.140 276.240 ;
        RECT 620.200 275.160 620.380 276.250 ;
        RECT 621.770 275.160 621.950 276.250 ;
        RECT 623.340 275.160 623.520 276.250 ;
        RECT 624.490 276.240 624.720 276.620 ;
        RECT 626.070 276.240 626.300 276.620 ;
        RECT 627.650 276.460 627.910 276.620 ;
        RECT 627.650 276.240 627.880 276.460 ;
        RECT 615.790 274.770 616.020 275.150 ;
        RECT 617.370 274.770 617.600 275.150 ;
        RECT 618.950 274.770 619.180 275.150 ;
        RECT 620.170 274.780 620.400 275.160 ;
        RECT 621.750 274.780 621.980 275.160 ;
        RECT 623.330 274.780 623.560 275.160 ;
        RECT 624.520 275.150 624.700 276.240 ;
        RECT 626.090 275.150 626.270 276.240 ;
        RECT 627.660 275.150 627.840 276.240 ;
        RECT 628.600 275.600 629.470 277.330 ;
        RECT 710.350 277.050 710.950 277.350 ;
        RECT 709.300 276.875 715.130 277.050 ;
        RECT 719.200 276.875 722.420 276.960 ;
        RECT 684.400 276.755 687.620 276.840 ;
        RECT 679.800 276.715 687.620 276.755 ;
        RECT 692.060 276.775 697.670 276.790 ;
        RECT 701.630 276.775 704.850 276.860 ;
        RECT 692.060 276.735 704.850 276.775 ;
        RECT 709.300 276.835 722.420 276.875 ;
        RECT 726.730 276.905 732.190 277.070 ;
        RECT 736.370 276.905 739.590 276.990 ;
        RECT 726.730 276.865 739.590 276.905 ;
        RECT 743.920 276.965 749.840 277.230 ;
        RECT 754.180 276.965 757.400 277.050 ;
        RECT 743.920 276.925 757.400 276.965 ;
        RECT 743.920 276.865 762.100 276.925 ;
        RECT 726.730 276.850 762.100 276.865 ;
        RECT 726.730 276.835 754.860 276.850 ;
        RECT 709.300 276.790 754.860 276.835 ;
        RECT 709.300 276.760 737.050 276.790 ;
        RECT 709.300 276.735 719.880 276.760 ;
        RECT 692.060 276.715 719.880 276.735 ;
        RECT 679.800 276.670 719.880 276.715 ;
        RECT 679.800 276.660 709.550 276.670 ;
        RECT 679.800 276.640 702.310 276.660 ;
        RECT 679.800 276.525 685.080 276.640 ;
        RECT 682.490 276.385 683.150 276.525 ;
        RECT 679.800 276.015 685.080 276.385 ;
        RECT 685.600 276.010 686.200 276.640 ;
        RECT 687.040 276.570 702.310 276.640 ;
        RECT 687.040 276.485 692.320 276.570 ;
        RECT 697.030 276.545 702.310 276.570 ;
        RECT 688.120 276.345 688.340 276.485 ;
        RECT 699.720 276.405 700.380 276.545 ;
        RECT 687.040 275.975 692.320 276.345 ;
        RECT 697.030 276.035 702.310 276.405 ;
        RECT 702.880 275.940 703.450 276.660 ;
        RECT 704.270 276.505 709.550 276.660 ;
        RECT 710.350 276.640 710.950 276.670 ;
        RECT 714.600 276.645 719.880 276.670 ;
        RECT 717.290 276.505 717.950 276.645 ;
        RECT 705.350 276.365 705.570 276.505 ;
        RECT 704.270 275.995 709.550 276.365 ;
        RECT 714.600 276.135 719.880 276.505 ;
        RECT 720.410 276.070 721.030 276.760 ;
        RECT 721.840 276.720 737.050 276.760 ;
        RECT 721.840 276.605 727.120 276.720 ;
        RECT 731.770 276.675 737.050 276.720 ;
        RECT 722.920 276.465 723.140 276.605 ;
        RECT 734.460 276.535 735.120 276.675 ;
        RECT 721.840 276.095 727.120 276.465 ;
        RECT 731.770 276.165 737.050 276.535 ;
        RECT 737.530 275.930 738.320 276.790 ;
        RECT 739.010 276.635 744.290 276.790 ;
        RECT 749.580 276.735 754.860 276.790 ;
        RECT 740.090 276.495 740.310 276.635 ;
        RECT 752.270 276.595 752.930 276.735 ;
        RECT 739.010 276.125 744.290 276.495 ;
        RECT 749.580 276.225 754.860 276.595 ;
        RECT 755.500 276.300 756.070 276.850 ;
        RECT 756.820 276.695 762.100 276.850 ;
        RECT 757.900 276.555 758.120 276.695 ;
        RECT 761.450 276.555 762.030 276.695 ;
        RECT 756.820 276.185 762.100 276.555 ;
        RECT 778.550 275.680 779.490 277.090 ;
        RECT 636.100 275.615 639.590 275.630 ;
        RECT 640.370 275.615 645.080 275.670 ;
        RECT 628.600 275.525 635.260 275.600 ;
        RECT 636.100 275.525 645.080 275.615 ;
        RECT 628.600 275.460 645.080 275.525 ;
        RECT 778.550 275.595 781.260 275.680 ;
        RECT 800.080 275.650 800.590 275.930 ;
        RECT 796.030 275.595 800.590 275.650 ;
        RECT 778.550 275.585 800.590 275.595 ;
        RECT 814.860 275.585 818.940 275.650 ;
        RECT 778.550 275.555 818.940 275.585 ;
        RECT 833.750 275.595 838.580 275.670 ;
        RECT 841.500 275.610 842.230 275.620 ;
        RECT 842.930 275.610 843.670 275.980 ;
        RECT 844.290 275.610 844.950 275.630 ;
        RECT 841.500 275.595 844.950 275.610 ;
        RECT 833.750 275.555 844.950 275.595 ;
        RECT 778.550 275.460 844.950 275.555 ;
        RECT 858.410 275.545 858.970 276.060 ;
        RECT 628.600 275.420 640.610 275.460 ;
        RECT 642.810 275.440 644.710 275.460 ;
        RECT 628.600 275.320 636.420 275.420 ;
        RECT 639.170 275.385 640.610 275.420 ;
        RECT 624.490 274.770 624.720 275.150 ;
        RECT 626.070 274.770 626.300 275.150 ;
        RECT 627.650 274.770 627.880 275.150 ;
        RECT 628.600 274.010 629.470 275.320 ;
        RECT 634.980 275.295 636.420 275.320 ;
        RECT 635.110 275.155 635.290 275.295 ;
        RECT 639.300 275.245 639.540 275.385 ;
        RECT 643.270 275.365 644.710 275.440 ;
        RECT 778.550 275.450 844.490 275.460 ;
        RECT 634.980 274.785 636.420 275.155 ;
        RECT 639.170 274.875 640.610 275.245 ;
        RECT 644.390 275.225 644.630 275.365 ;
        RECT 778.550 275.270 779.490 275.450 ;
        RECT 780.960 275.440 834.060 275.450 ;
        RECT 780.960 275.365 796.320 275.440 ;
        RECT 643.270 275.170 644.710 275.225 ;
        RECT 645.290 275.170 645.930 275.210 ;
        RECT 643.270 274.900 645.930 275.170 ;
        RECT 643.270 274.855 644.710 274.900 ;
        RECT 645.290 273.900 645.930 274.900 ;
        RECT 756.300 274.370 756.890 274.470 ;
        RECT 760.280 274.370 760.520 274.590 ;
        RECT 756.160 274.240 760.520 274.370 ;
        RECT 756.160 274.180 760.490 274.240 ;
        RECT 756.300 273.650 756.890 274.180 ;
        RECT 404.960 270.390 405.190 270.760 ;
        RECT 408.250 270.390 408.480 271.370 ;
        RECT 409.480 270.730 411.160 271.470 ;
        RECT 682.870 271.085 686.090 271.120 ;
        RECT 688.590 271.105 691.350 271.220 ;
        RECT 700.100 271.105 703.320 271.140 ;
        RECT 705.820 271.125 708.580 271.240 ;
        RECT 717.670 271.205 720.890 271.240 ;
        RECT 723.390 271.225 726.150 271.340 ;
        RECT 734.840 271.235 738.060 271.270 ;
        RECT 740.560 271.255 743.320 271.370 ;
        RECT 745.800 271.285 749.910 271.320 ;
        RECT 752.650 271.295 755.870 271.330 ;
        RECT 758.370 271.315 761.130 271.430 ;
        RECT 758.370 271.295 764.070 271.315 ;
        RECT 752.650 271.285 764.070 271.295 ;
        RECT 745.800 271.255 764.070 271.285 ;
        RECT 740.560 271.235 764.070 271.255 ;
        RECT 734.840 271.225 764.070 271.235 ;
        RECT 723.390 271.205 729.090 271.225 ;
        RECT 717.670 271.200 729.090 271.205 ;
        RECT 731.890 271.200 764.070 271.225 ;
        RECT 768.270 271.200 768.840 271.260 ;
        RECT 717.670 271.195 768.840 271.200 ;
        RECT 714.720 271.170 768.840 271.195 ;
        RECT 714.720 271.130 758.720 271.170 ;
        RECT 705.820 271.105 711.520 271.125 ;
        RECT 688.590 271.085 694.290 271.105 ;
        RECT 700.100 271.095 711.520 271.105 ;
        RECT 682.870 271.075 694.290 271.085 ;
        RECT 679.920 270.960 694.290 271.075 ;
        RECT 679.920 270.920 688.940 270.960 ;
        RECT 679.920 270.845 683.280 270.920 ;
        RECT 685.580 270.855 688.940 270.920 ;
        RECT 409.480 270.540 410.640 270.730 ;
        RECT 682.050 270.705 682.680 270.845 ;
        RECT 687.710 270.715 687.950 270.855 ;
        RECT 679.920 270.335 683.280 270.705 ;
        RECT 685.580 270.345 688.940 270.715 ;
        RECT 689.580 270.120 690.280 270.960 ;
        RECT 690.930 270.875 694.290 270.960 ;
        RECT 697.150 270.980 711.520 271.095 ;
        RECT 697.150 270.940 706.170 270.980 ;
        RECT 692.920 270.735 693.160 270.875 ;
        RECT 697.150 270.865 700.510 270.940 ;
        RECT 690.930 270.365 694.290 270.735 ;
        RECT 699.280 270.725 699.910 270.865 ;
        RECT 697.150 270.355 700.510 270.725 ;
        RECT 701.020 270.120 701.720 270.940 ;
        RECT 702.810 270.875 706.170 270.940 ;
        RECT 708.160 270.895 711.520 270.980 ;
        RECT 714.720 271.110 753.060 271.130 ;
        RECT 714.720 271.080 740.910 271.110 ;
        RECT 714.720 271.040 723.740 271.080 ;
        RECT 714.720 270.965 718.080 271.040 ;
        RECT 704.940 270.735 705.180 270.875 ;
        RECT 710.150 270.755 710.390 270.895 ;
        RECT 716.850 270.825 717.480 270.965 ;
        RECT 702.810 270.365 706.170 270.735 ;
        RECT 708.160 270.385 711.520 270.755 ;
        RECT 714.720 270.455 718.080 270.825 ;
        RECT 718.600 270.360 719.300 271.040 ;
        RECT 720.380 270.975 723.740 271.040 ;
        RECT 725.730 271.070 740.910 271.080 ;
        RECT 725.730 271.020 735.250 271.070 ;
        RECT 725.730 270.995 729.090 271.020 ;
        RECT 722.510 270.835 722.750 270.975 ;
        RECT 727.720 270.855 727.960 270.995 ;
        RECT 729.270 270.990 731.650 271.020 ;
        RECT 731.890 270.995 735.250 271.020 ;
        RECT 734.020 270.855 734.650 270.995 ;
        RECT 720.380 270.465 723.740 270.835 ;
        RECT 725.730 270.485 729.090 270.855 ;
        RECT 731.890 270.485 735.250 270.855 ;
        RECT 735.930 270.260 736.630 271.070 ;
        RECT 737.550 271.005 740.910 271.070 ;
        RECT 742.900 271.080 753.060 271.110 ;
        RECT 742.900 271.025 746.260 271.080 ;
        RECT 749.700 271.055 753.060 271.080 ;
        RECT 739.680 270.865 739.920 271.005 ;
        RECT 744.890 270.885 745.130 271.025 ;
        RECT 751.830 270.915 752.460 271.055 ;
        RECT 737.550 270.495 740.910 270.865 ;
        RECT 742.900 270.515 746.260 270.885 ;
        RECT 749.700 270.545 753.060 270.915 ;
        RECT 753.870 270.300 754.490 271.130 ;
        RECT 755.360 271.065 758.720 271.130 ;
        RECT 760.710 271.085 768.840 271.170 ;
        RECT 757.490 270.925 757.730 271.065 ;
        RECT 762.700 270.945 768.840 271.085 ;
        RECT 755.360 270.555 758.720 270.925 ;
        RECT 760.710 270.720 768.840 270.945 ;
        RECT 760.710 270.575 764.070 270.720 ;
        RECT 756.430 268.640 756.850 268.700 ;
        RECT 756.410 268.060 756.870 268.640 ;
        RECT 756.430 268.000 756.850 268.060 ;
        RECT 395.090 266.920 395.320 267.900 ;
        RECT 398.380 266.920 398.610 267.900 ;
        RECT 401.670 266.920 401.900 267.900 ;
        RECT 404.960 266.920 405.190 267.900 ;
        RECT 408.250 266.920 408.480 267.900 ;
        RECT 395.090 263.450 395.320 264.430 ;
        RECT 398.380 263.450 398.610 264.430 ;
        RECT 401.670 263.450 401.900 264.430 ;
        RECT 404.960 263.450 405.190 264.430 ;
        RECT 408.250 263.450 408.480 264.430 ;
        RECT 589.860 262.380 590.960 262.690 ;
        RECT 600.070 262.380 631.560 262.430 ;
        RECT 589.860 261.660 631.560 262.380 ;
        RECT 589.860 261.480 590.960 261.660 ;
        RECT 600.070 261.610 631.560 261.660 ;
        RECT 395.090 259.980 395.320 260.960 ;
        RECT 398.380 259.980 398.610 260.960 ;
        RECT 401.670 259.980 401.900 260.960 ;
        RECT 404.960 259.980 405.190 260.960 ;
        RECT 408.250 259.980 408.480 260.960 ;
        RECT 600.750 259.310 601.460 261.610 ;
        RECT 600.750 257.520 601.490 259.310 ;
        RECT 602.160 259.230 602.410 261.610 ;
        RECT 609.850 259.240 610.100 261.610 ;
        RECT 602.160 259.070 605.570 259.230 ;
        RECT 606.710 259.080 610.100 259.240 ;
        RECT 602.160 258.760 602.410 259.070 ;
        RECT 603.770 258.900 603.940 259.070 ;
        RECT 605.370 258.900 605.540 259.070 ;
        RECT 606.720 258.910 606.890 259.080 ;
        RECT 608.290 258.910 608.460 259.080 ;
        RECT 602.170 258.520 602.400 258.760 ;
        RECT 603.750 258.520 603.980 258.900 ;
        RECT 605.330 258.520 605.560 258.900 ;
        RECT 606.690 258.530 606.920 258.910 ;
        RECT 608.270 258.530 608.500 258.910 ;
        RECT 609.850 258.770 610.100 259.080 ;
        RECT 611.210 259.240 611.460 261.610 ;
        RECT 611.210 259.080 614.610 259.240 ;
        RECT 618.790 259.220 619.030 261.610 ;
        RECT 620.010 259.230 620.260 261.610 ;
        RECT 609.850 258.530 610.080 258.770 ;
        RECT 611.210 258.660 611.460 259.080 ;
        RECT 612.810 258.910 612.980 259.080 ;
        RECT 614.410 258.910 614.580 259.080 ;
        RECT 615.660 259.060 619.040 259.220 ;
        RECT 620.010 259.070 623.420 259.230 ;
        RECT 627.510 259.220 627.760 261.610 ;
        RECT 628.590 259.600 629.300 261.610 ;
        RECT 684.370 260.895 696.940 261.110 ;
        RECT 710.100 261.060 710.700 261.070 ;
        RECT 701.640 260.895 714.840 261.060 ;
        RECT 719.360 260.895 732.560 261.040 ;
        RECT 736.580 260.905 749.780 261.040 ;
        RECT 736.580 260.895 754.420 260.905 ;
        RECT 684.370 260.885 754.420 260.895 ;
        RECT 679.370 260.840 754.420 260.885 ;
        RECT 768.270 260.840 768.840 270.720 ;
        RECT 778.760 268.050 779.000 275.270 ;
        RECT 784.020 275.225 784.190 275.365 ;
        RECT 780.960 274.855 796.320 275.225 ;
        RECT 796.690 274.920 797.460 275.440 ;
        RECT 799.850 275.355 815.210 275.440 ;
        RECT 802.890 275.215 803.060 275.355 ;
        RECT 799.850 274.845 815.210 275.215 ;
        RECT 815.690 274.980 816.640 275.440 ;
        RECT 818.700 275.325 834.060 275.440 ;
        RECT 821.750 275.185 821.920 275.325 ;
        RECT 818.700 274.815 834.060 275.185 ;
        RECT 837.120 274.930 837.810 275.450 ;
        RECT 838.420 275.365 842.260 275.450 ;
        RECT 841.370 275.225 842.230 275.365 ;
        RECT 838.420 274.855 842.260 275.225 ;
        RECT 844.770 273.335 844.910 275.460 ;
        RECT 855.930 275.315 859.290 275.545 ;
        RECT 858.330 275.175 858.550 275.315 ;
        RECT 855.930 274.805 859.290 275.175 ;
        RECT 847.650 273.345 850.160 273.370 ;
        RECT 847.650 273.335 851.520 273.345 ;
        RECT 844.670 273.210 851.520 273.335 ;
        RECT 844.670 273.105 848.030 273.210 ;
        RECT 850.080 273.115 851.520 273.210 ;
        RECT 846.220 272.965 846.410 273.105 ;
        RECT 850.220 272.975 850.410 273.115 ;
        RECT 844.670 272.595 848.030 272.965 ;
        RECT 850.080 272.605 851.520 272.975 ;
        RECT 860.810 272.690 861.830 273.700 ;
        RECT 861.380 272.155 861.620 272.690 ;
        RECT 863.500 272.155 864.350 272.380 ;
        RECT 861.250 271.925 864.610 272.155 ;
        RECT 862.670 271.785 864.350 271.925 ;
        RECT 861.250 271.415 864.610 271.785 ;
        RECT 841.370 270.035 841.860 270.460 ;
        RECT 838.430 269.890 841.860 270.035 ;
        RECT 838.430 269.805 841.790 269.890 ;
        RECT 841.020 269.665 841.200 269.805 ;
        RECT 838.430 269.295 841.790 269.665 ;
        RECT 858.570 268.875 859.130 269.350 ;
        RECT 856.010 268.645 859.370 268.875 ;
        RECT 858.040 268.505 858.260 268.645 ;
        RECT 795.950 268.095 799.790 268.140 ;
        RECT 856.010 268.135 859.370 268.505 ;
        RECT 778.760 268.035 781.280 268.050 ;
        RECT 795.950 268.035 814.860 268.095 ;
        RECT 778.760 267.930 814.860 268.035 ;
        RECT 778.760 267.890 796.330 267.930 ;
        RECT 778.760 267.880 779.000 267.890 ;
        RECT 780.970 267.805 796.330 267.890 ;
        RECT 793.610 267.665 793.780 267.805 ;
        RECT 780.970 267.295 796.330 267.665 ;
        RECT 796.670 267.460 797.240 267.930 ;
        RECT 799.500 267.865 814.860 267.930 ;
        RECT 802.550 267.725 802.720 267.865 ;
        RECT 799.500 267.670 814.860 267.725 ;
        RECT 815.170 267.670 815.620 268.020 ;
        RECT 799.500 267.520 815.620 267.670 ;
        RECT 799.500 267.355 814.860 267.520 ;
        RECT 815.170 267.430 815.620 267.520 ;
        RECT 679.370 260.770 768.840 260.840 ;
        RECT 679.370 260.750 701.930 260.770 ;
        RECT 679.370 260.740 690.220 260.750 ;
        RECT 690.780 260.740 701.930 260.750 ;
        RECT 679.370 260.655 684.650 260.740 ;
        RECT 681.660 260.515 681.840 260.655 ;
        RECT 679.370 260.145 684.650 260.515 ;
        RECT 685.180 260.060 685.760 260.740 ;
        RECT 696.650 260.665 701.930 260.740 ;
        RECT 698.270 260.525 698.450 260.665 ;
        RECT 699.820 260.525 700.120 260.665 ;
        RECT 696.650 260.155 701.930 260.525 ;
        RECT 702.370 260.200 703.050 260.770 ;
        RECT 710.100 260.360 710.700 260.770 ;
        RECT 714.420 260.750 768.840 260.770 ;
        RECT 714.420 260.665 719.700 260.750 ;
        RECT 717.210 260.525 717.510 260.665 ;
        RECT 714.420 260.155 719.700 260.525 ;
        RECT 720.250 260.210 720.730 260.750 ;
        RECT 731.660 260.665 736.940 260.750 ;
        RECT 734.150 260.525 734.410 260.665 ;
        RECT 731.660 260.155 736.940 260.525 ;
        RECT 737.360 260.390 737.870 260.750 ;
        RECT 749.140 260.675 768.840 260.750 ;
        RECT 752.120 260.535 768.840 260.675 ;
        RECT 749.140 260.270 768.840 260.535 ;
        RECT 749.140 260.165 754.420 260.270 ;
        RECT 755.010 259.840 755.580 260.270 ;
        RECT 768.270 260.240 768.840 260.270 ;
        RECT 611.210 258.530 611.440 258.660 ;
        RECT 612.790 258.530 613.020 258.910 ;
        RECT 614.370 258.530 614.600 258.910 ;
        RECT 615.670 258.890 615.840 259.060 ;
        RECT 617.240 258.890 617.410 259.060 ;
        RECT 395.090 256.510 395.320 257.490 ;
        RECT 398.380 256.510 398.610 257.490 ;
        RECT 401.670 256.510 401.900 257.490 ;
        RECT 404.960 256.510 405.190 257.490 ;
        RECT 408.250 256.510 408.480 257.490 ;
        RECT 596.080 257.345 601.490 257.520 ;
        RECT 602.200 257.430 602.380 258.520 ;
        RECT 603.770 257.430 603.950 258.520 ;
        RECT 605.340 257.430 605.520 258.520 ;
        RECT 606.720 257.440 606.900 258.530 ;
        RECT 608.290 257.440 608.470 258.530 ;
        RECT 609.860 257.440 610.040 258.530 ;
        RECT 611.240 257.440 611.420 258.530 ;
        RECT 612.810 257.440 612.990 258.530 ;
        RECT 614.380 257.440 614.560 258.530 ;
        RECT 615.640 258.510 615.870 258.890 ;
        RECT 617.220 258.510 617.450 258.890 ;
        RECT 618.790 258.710 619.030 259.060 ;
        RECT 620.010 258.760 620.260 259.070 ;
        RECT 621.620 258.900 621.790 259.070 ;
        RECT 623.220 258.900 623.390 259.070 ;
        RECT 624.360 259.060 627.760 259.220 ;
        RECT 618.800 258.510 619.030 258.710 ;
        RECT 620.020 258.520 620.250 258.760 ;
        RECT 621.600 258.520 621.830 258.900 ;
        RECT 623.180 258.520 623.410 258.900 ;
        RECT 624.370 258.890 624.540 259.060 ;
        RECT 625.940 258.890 626.110 259.060 ;
        RECT 627.510 258.890 627.760 259.060 ;
        RECT 594.940 257.170 601.490 257.345 ;
        RECT 594.940 257.115 596.380 257.170 ;
        RECT 596.060 256.975 596.200 257.115 ;
        RECT 594.940 256.605 596.380 256.975 ;
        RECT 600.750 256.450 601.490 257.170 ;
        RECT 602.170 257.050 602.400 257.430 ;
        RECT 603.750 257.050 603.980 257.430 ;
        RECT 605.330 257.050 605.560 257.430 ;
        RECT 606.690 257.060 606.920 257.440 ;
        RECT 608.270 257.060 608.500 257.440 ;
        RECT 609.850 257.060 610.080 257.440 ;
        RECT 611.210 257.060 611.440 257.440 ;
        RECT 612.790 257.060 613.020 257.440 ;
        RECT 614.370 257.060 614.600 257.440 ;
        RECT 615.670 257.420 615.850 258.510 ;
        RECT 617.240 257.420 617.420 258.510 ;
        RECT 618.810 257.420 618.990 258.510 ;
        RECT 620.050 257.430 620.230 258.520 ;
        RECT 621.620 257.430 621.800 258.520 ;
        RECT 623.190 257.430 623.370 258.520 ;
        RECT 624.340 258.510 624.570 258.890 ;
        RECT 625.920 258.510 626.150 258.890 ;
        RECT 627.500 258.730 627.760 258.890 ;
        RECT 627.500 258.510 627.730 258.730 ;
        RECT 615.640 257.040 615.870 257.420 ;
        RECT 617.220 257.040 617.450 257.420 ;
        RECT 618.800 257.040 619.030 257.420 ;
        RECT 620.020 257.050 620.250 257.430 ;
        RECT 621.600 257.050 621.830 257.430 ;
        RECT 623.180 257.050 623.410 257.430 ;
        RECT 624.370 257.420 624.550 258.510 ;
        RECT 625.940 257.420 626.120 258.510 ;
        RECT 627.510 257.420 627.690 258.510 ;
        RECT 628.450 257.870 629.320 259.600 ;
        RECT 858.390 259.565 858.950 260.060 ;
        RECT 855.880 259.540 859.240 259.565 ;
        RECT 860.790 259.540 861.530 259.580 ;
        RECT 855.880 259.410 861.530 259.540 ;
        RECT 855.880 259.400 860.870 259.410 ;
        RECT 855.880 259.335 859.240 259.400 ;
        RECT 857.750 259.195 857.970 259.335 ;
        RECT 855.880 258.825 859.240 259.195 ;
        RECT 860.300 257.990 861.080 258.270 ;
        RECT 861.380 257.990 861.530 259.410 ;
        RECT 635.950 257.885 639.440 257.900 ;
        RECT 640.220 257.885 644.930 257.940 ;
        RECT 628.450 257.795 635.110 257.870 ;
        RECT 635.950 257.795 644.930 257.885 ;
        RECT 628.450 257.730 644.930 257.795 ;
        RECT 860.300 257.750 861.530 257.990 ;
        RECT 628.450 257.690 640.460 257.730 ;
        RECT 642.660 257.710 644.560 257.730 ;
        RECT 628.450 257.590 636.270 257.690 ;
        RECT 639.020 257.655 640.460 257.690 ;
        RECT 624.340 257.040 624.570 257.420 ;
        RECT 625.920 257.040 626.150 257.420 ;
        RECT 627.500 257.040 627.730 257.420 ;
        RECT 628.450 256.280 629.320 257.590 ;
        RECT 634.830 257.565 636.270 257.590 ;
        RECT 634.960 257.425 635.140 257.565 ;
        RECT 639.150 257.515 639.390 257.655 ;
        RECT 643.120 257.635 644.560 257.710 ;
        RECT 634.830 257.055 636.270 257.425 ;
        RECT 639.020 257.145 640.460 257.515 ;
        RECT 644.240 257.495 644.480 257.635 ;
        RECT 643.120 257.380 644.560 257.495 ;
        RECT 860.300 257.450 861.080 257.750 ;
        RECT 643.120 257.370 645.310 257.380 ;
        RECT 643.120 257.125 645.690 257.370 ;
        RECT 644.200 257.110 645.690 257.125 ;
        RECT 645.050 256.060 645.690 257.110 ;
        RECT 861.380 257.075 861.530 257.750 ;
        RECT 863.550 257.075 864.260 257.270 ;
        RECT 861.190 256.845 864.550 257.075 ;
        RECT 862.360 256.705 864.260 256.845 ;
        RECT 861.190 256.335 864.550 256.705 ;
        RECT 211.570 255.360 212.550 255.590 ;
        RECT 215.040 255.360 216.020 255.590 ;
        RECT 218.510 255.360 219.490 255.590 ;
        RECT 221.980 255.360 222.960 255.590 ;
        RECT 225.450 255.360 226.430 255.590 ;
        RECT 231.540 255.360 232.520 255.590 ;
        RECT 235.010 255.360 235.990 255.590 ;
        RECT 238.480 255.360 239.460 255.590 ;
        RECT 241.950 255.360 242.930 255.590 ;
        RECT 245.420 255.360 246.400 255.590 ;
        RECT 251.650 255.360 252.630 255.590 ;
        RECT 255.120 255.360 256.100 255.590 ;
        RECT 258.590 255.360 259.570 255.590 ;
        RECT 262.060 255.360 263.040 255.590 ;
        RECT 265.530 255.360 266.510 255.590 ;
        RECT 271.760 255.360 272.740 255.590 ;
        RECT 275.230 255.360 276.210 255.590 ;
        RECT 278.700 255.360 279.680 255.590 ;
        RECT 282.170 255.360 283.150 255.590 ;
        RECT 285.640 255.360 286.620 255.590 ;
        RECT 710.330 255.520 710.930 255.820 ;
        RECT 709.280 255.345 715.110 255.520 ;
        RECT 719.180 255.345 722.400 255.430 ;
        RECT 684.380 255.225 687.600 255.310 ;
        RECT 679.780 255.185 687.600 255.225 ;
        RECT 692.040 255.245 697.650 255.260 ;
        RECT 701.610 255.245 704.830 255.330 ;
        RECT 692.040 255.205 704.830 255.245 ;
        RECT 709.280 255.305 722.400 255.345 ;
        RECT 726.710 255.375 732.170 255.540 ;
        RECT 736.350 255.375 739.570 255.460 ;
        RECT 726.710 255.335 739.570 255.375 ;
        RECT 743.900 255.435 749.820 255.700 ;
        RECT 754.160 255.435 757.380 255.520 ;
        RECT 743.900 255.395 757.380 255.435 ;
        RECT 743.900 255.335 762.080 255.395 ;
        RECT 726.710 255.320 762.080 255.335 ;
        RECT 726.710 255.305 754.840 255.320 ;
        RECT 709.280 255.260 754.840 255.305 ;
        RECT 709.280 255.230 737.030 255.260 ;
        RECT 709.280 255.205 719.860 255.230 ;
        RECT 692.040 255.185 719.860 255.205 ;
        RECT 679.780 255.140 719.860 255.185 ;
        RECT 679.780 255.130 709.530 255.140 ;
        RECT 679.780 255.110 702.290 255.130 ;
        RECT 4.630 254.610 5.610 254.840 ;
        RECT 8.100 254.610 9.080 254.840 ;
        RECT 11.570 254.610 12.550 254.840 ;
        RECT 17.970 254.590 18.950 254.820 ;
        RECT 21.440 254.590 22.420 254.820 ;
        RECT 24.910 254.590 25.890 254.820 ;
        RECT 31.340 254.620 32.320 254.850 ;
        RECT 34.810 254.620 35.790 254.850 ;
        RECT 38.280 254.620 39.260 254.850 ;
        RECT 44.570 254.620 45.550 254.850 ;
        RECT 48.040 254.620 49.020 254.850 ;
        RECT 51.510 254.620 52.490 254.850 ;
        RECT 57.840 254.590 58.820 254.820 ;
        RECT 61.310 254.590 62.290 254.820 ;
        RECT 64.780 254.590 65.760 254.820 ;
        RECT 71.110 254.620 72.090 254.850 ;
        RECT 74.580 254.620 75.560 254.850 ;
        RECT 78.050 254.620 79.030 254.850 ;
        RECT 84.240 254.640 85.220 254.870 ;
        RECT 87.710 254.640 88.690 254.870 ;
        RECT 91.180 254.640 92.160 254.870 ;
        RECT 97.660 254.860 98.640 255.090 ;
        RECT 101.130 254.860 102.110 255.090 ;
        RECT 679.780 254.995 685.060 255.110 ;
        RECT 682.470 254.855 683.130 254.995 ;
        RECT 679.780 254.485 685.060 254.855 ;
        RECT 685.550 254.350 686.110 255.110 ;
        RECT 687.020 255.040 702.290 255.110 ;
        RECT 687.020 254.955 692.300 255.040 ;
        RECT 688.100 254.815 688.320 254.955 ;
        RECT 687.020 254.445 692.300 254.815 ;
        RECT 695.880 253.140 696.150 255.040 ;
        RECT 697.010 255.015 702.290 255.040 ;
        RECT 699.700 254.875 700.360 255.015 ;
        RECT 697.010 254.505 702.290 254.875 ;
        RECT 702.800 254.410 703.440 255.130 ;
        RECT 704.250 254.975 709.530 255.130 ;
        RECT 710.330 255.110 710.930 255.140 ;
        RECT 714.580 255.115 719.860 255.140 ;
        RECT 717.270 254.975 717.930 255.115 ;
        RECT 705.330 254.835 705.550 254.975 ;
        RECT 704.250 254.465 709.530 254.835 ;
        RECT 714.580 254.605 719.860 254.975 ;
        RECT 720.340 254.470 720.850 255.230 ;
        RECT 721.820 255.190 737.030 255.230 ;
        RECT 721.820 255.075 727.100 255.190 ;
        RECT 731.750 255.145 737.030 255.190 ;
        RECT 722.900 254.935 723.120 255.075 ;
        RECT 734.440 255.005 735.100 255.145 ;
        RECT 721.820 254.565 727.100 254.935 ;
        RECT 731.750 254.635 737.030 255.005 ;
        RECT 737.520 254.580 738.160 255.260 ;
        RECT 738.990 255.105 744.270 255.260 ;
        RECT 749.560 255.205 754.840 255.260 ;
        RECT 740.070 254.965 740.290 255.105 ;
        RECT 752.250 255.065 752.910 255.205 ;
        RECT 738.990 254.595 744.270 254.965 ;
        RECT 749.560 254.695 754.840 255.065 ;
        RECT 755.280 254.720 755.850 255.320 ;
        RECT 756.800 255.165 762.080 255.320 ;
        RECT 757.880 255.025 758.100 255.165 ;
        RECT 756.800 254.655 762.080 255.025 ;
        RECT 858.480 253.795 859.040 254.280 ;
        RECT 855.940 253.565 859.300 253.795 ;
        RECT 857.990 253.425 858.210 253.565 ;
        RECT 697.000 253.140 697.560 253.380 ;
        RECT 699.050 253.140 699.310 253.270 ;
        RECT 695.880 252.970 699.310 253.140 ;
        RECT 855.940 253.055 859.300 253.425 ;
        RECT 695.880 252.960 696.430 252.970 ;
        RECT 695.920 252.940 696.430 252.960 ;
        RECT 697.000 252.880 697.560 252.970 ;
        RECT 699.050 252.900 699.310 252.970 ;
        RECT 211.570 252.070 212.550 252.300 ;
        RECT 215.040 252.070 216.020 252.300 ;
        RECT 218.510 252.070 219.490 252.300 ;
        RECT 221.980 252.070 222.960 252.300 ;
        RECT 225.450 252.070 226.430 252.300 ;
        RECT 231.540 252.070 232.520 252.300 ;
        RECT 235.010 252.070 235.990 252.300 ;
        RECT 238.480 252.070 239.460 252.300 ;
        RECT 241.950 252.070 242.930 252.300 ;
        RECT 245.420 252.070 246.400 252.300 ;
        RECT 251.650 252.070 252.630 252.300 ;
        RECT 255.120 252.070 256.100 252.300 ;
        RECT 258.590 252.070 259.570 252.300 ;
        RECT 262.060 252.070 263.040 252.300 ;
        RECT 265.530 252.070 266.510 252.300 ;
        RECT 271.760 252.070 272.740 252.300 ;
        RECT 275.230 252.070 276.210 252.300 ;
        RECT 278.700 252.070 279.680 252.300 ;
        RECT 282.170 252.070 283.150 252.300 ;
        RECT 285.640 252.070 286.620 252.300 ;
        RECT 4.630 251.320 5.610 251.550 ;
        RECT 8.100 251.320 9.080 251.550 ;
        RECT 11.570 251.320 12.550 251.550 ;
        RECT 17.970 251.300 18.950 251.530 ;
        RECT 21.440 251.300 22.420 251.530 ;
        RECT 24.910 251.300 25.890 251.530 ;
        RECT 31.340 251.330 32.320 251.560 ;
        RECT 34.810 251.330 35.790 251.560 ;
        RECT 38.280 251.330 39.260 251.560 ;
        RECT 44.570 251.330 45.550 251.560 ;
        RECT 48.040 251.330 49.020 251.560 ;
        RECT 51.510 251.330 52.490 251.560 ;
        RECT 57.840 251.300 58.820 251.530 ;
        RECT 61.310 251.300 62.290 251.530 ;
        RECT 64.780 251.300 65.760 251.530 ;
        RECT 71.110 251.330 72.090 251.560 ;
        RECT 74.580 251.330 75.560 251.560 ;
        RECT 78.050 251.330 79.030 251.560 ;
        RECT 84.240 251.350 85.220 251.580 ;
        RECT 87.710 251.350 88.690 251.580 ;
        RECT 91.180 251.350 92.160 251.580 ;
        RECT 97.660 251.570 98.640 251.800 ;
        RECT 101.130 251.570 102.110 251.800 ;
        RECT 682.850 249.555 686.070 249.590 ;
        RECT 688.570 249.575 691.330 249.690 ;
        RECT 700.080 249.575 703.300 249.610 ;
        RECT 705.800 249.595 708.560 249.710 ;
        RECT 717.650 249.675 720.870 249.710 ;
        RECT 723.370 249.695 726.130 249.810 ;
        RECT 734.820 249.705 738.040 249.740 ;
        RECT 740.540 249.725 743.300 249.840 ;
        RECT 745.780 249.755 749.890 249.790 ;
        RECT 752.630 249.765 755.850 249.800 ;
        RECT 758.350 249.785 761.110 249.900 ;
        RECT 758.350 249.765 764.050 249.785 ;
        RECT 752.630 249.755 764.050 249.765 ;
        RECT 745.780 249.725 764.050 249.755 ;
        RECT 740.540 249.705 764.050 249.725 ;
        RECT 734.820 249.695 764.050 249.705 ;
        RECT 723.370 249.675 729.070 249.695 ;
        RECT 717.650 249.670 729.070 249.675 ;
        RECT 731.870 249.670 764.050 249.695 ;
        RECT 717.650 249.665 764.050 249.670 ;
        RECT 714.700 249.640 764.050 249.665 ;
        RECT 714.700 249.600 758.700 249.640 ;
        RECT 705.800 249.575 711.500 249.595 ;
        RECT 688.570 249.555 694.270 249.575 ;
        RECT 700.080 249.565 711.500 249.575 ;
        RECT 682.850 249.545 694.270 249.555 ;
        RECT 679.900 249.430 694.270 249.545 ;
        RECT 679.900 249.390 688.920 249.430 ;
        RECT 679.900 249.315 683.260 249.390 ;
        RECT 682.030 249.175 682.660 249.315 ;
        RECT 211.570 248.780 212.550 249.010 ;
        RECT 215.040 248.780 216.020 249.010 ;
        RECT 218.510 248.780 219.490 249.010 ;
        RECT 221.980 248.780 222.960 249.010 ;
        RECT 225.450 248.780 226.430 249.010 ;
        RECT 231.540 248.780 232.520 249.010 ;
        RECT 235.010 248.780 235.990 249.010 ;
        RECT 238.480 248.780 239.460 249.010 ;
        RECT 241.950 248.780 242.930 249.010 ;
        RECT 245.420 248.780 246.400 249.010 ;
        RECT 251.650 248.780 252.630 249.010 ;
        RECT 255.120 248.780 256.100 249.010 ;
        RECT 258.590 248.780 259.570 249.010 ;
        RECT 262.060 248.780 263.040 249.010 ;
        RECT 265.530 248.780 266.510 249.010 ;
        RECT 271.760 248.780 272.740 249.010 ;
        RECT 275.230 248.780 276.210 249.010 ;
        RECT 278.700 248.780 279.680 249.010 ;
        RECT 282.170 248.780 283.150 249.010 ;
        RECT 285.640 248.780 286.620 249.010 ;
        RECT 679.900 248.805 683.260 249.175 ;
        RECT 684.000 248.700 684.510 249.390 ;
        RECT 685.560 249.325 688.920 249.390 ;
        RECT 690.910 249.345 694.270 249.430 ;
        RECT 697.130 249.450 711.500 249.565 ;
        RECT 697.130 249.410 706.150 249.450 ;
        RECT 687.690 249.185 687.930 249.325 ;
        RECT 692.900 249.205 693.140 249.345 ;
        RECT 697.130 249.335 700.490 249.410 ;
        RECT 685.560 248.815 688.920 249.185 ;
        RECT 690.910 248.835 694.270 249.205 ;
        RECT 699.260 249.195 699.890 249.335 ;
        RECT 697.130 248.825 700.490 249.195 ;
        RECT 701.140 248.610 701.830 249.410 ;
        RECT 702.790 249.345 706.150 249.410 ;
        RECT 708.140 249.365 711.500 249.450 ;
        RECT 714.700 249.580 753.040 249.600 ;
        RECT 714.700 249.550 740.890 249.580 ;
        RECT 714.700 249.510 723.720 249.550 ;
        RECT 714.700 249.435 718.060 249.510 ;
        RECT 704.920 249.205 705.160 249.345 ;
        RECT 710.130 249.225 710.370 249.365 ;
        RECT 716.830 249.295 717.460 249.435 ;
        RECT 702.790 248.835 706.150 249.205 ;
        RECT 708.140 248.855 711.500 249.225 ;
        RECT 714.700 248.925 718.060 249.295 ;
        RECT 718.370 248.710 719.290 249.510 ;
        RECT 720.360 249.445 723.720 249.510 ;
        RECT 725.710 249.540 740.890 249.550 ;
        RECT 725.710 249.490 735.230 249.540 ;
        RECT 725.710 249.465 729.070 249.490 ;
        RECT 722.490 249.305 722.730 249.445 ;
        RECT 727.700 249.325 727.940 249.465 ;
        RECT 729.250 249.460 731.630 249.490 ;
        RECT 731.870 249.465 735.230 249.490 ;
        RECT 734.000 249.325 734.630 249.465 ;
        RECT 720.360 248.935 723.720 249.305 ;
        RECT 725.710 248.955 729.070 249.325 ;
        RECT 731.870 248.955 735.230 249.325 ;
        RECT 735.890 248.750 736.560 249.540 ;
        RECT 737.530 249.475 740.890 249.540 ;
        RECT 742.880 249.550 753.040 249.580 ;
        RECT 742.880 249.495 746.240 249.550 ;
        RECT 749.680 249.525 753.040 249.550 ;
        RECT 739.660 249.335 739.900 249.475 ;
        RECT 744.870 249.355 745.110 249.495 ;
        RECT 751.810 249.385 752.440 249.525 ;
        RECT 737.530 248.965 740.890 249.335 ;
        RECT 742.880 248.985 746.240 249.355 ;
        RECT 749.680 249.015 753.040 249.385 ;
        RECT 753.730 248.830 754.360 249.600 ;
        RECT 755.340 249.535 758.700 249.600 ;
        RECT 760.690 249.555 764.050 249.640 ;
        RECT 757.470 249.395 757.710 249.535 ;
        RECT 762.680 249.415 762.920 249.555 ;
        RECT 755.340 249.025 758.700 249.395 ;
        RECT 760.690 249.045 764.050 249.415 ;
        RECT 4.630 248.030 5.610 248.260 ;
        RECT 8.100 248.030 9.080 248.260 ;
        RECT 11.570 248.030 12.550 248.260 ;
        RECT 17.970 248.010 18.950 248.240 ;
        RECT 21.440 248.010 22.420 248.240 ;
        RECT 24.910 248.010 25.890 248.240 ;
        RECT 31.340 248.040 32.320 248.270 ;
        RECT 34.810 248.040 35.790 248.270 ;
        RECT 38.280 248.040 39.260 248.270 ;
        RECT 44.570 248.040 45.550 248.270 ;
        RECT 48.040 248.040 49.020 248.270 ;
        RECT 51.510 248.040 52.490 248.270 ;
        RECT 57.840 248.010 58.820 248.240 ;
        RECT 61.310 248.010 62.290 248.240 ;
        RECT 64.780 248.010 65.760 248.240 ;
        RECT 71.110 248.040 72.090 248.270 ;
        RECT 74.580 248.040 75.560 248.270 ;
        RECT 78.050 248.040 79.030 248.270 ;
        RECT 84.240 248.060 85.220 248.290 ;
        RECT 87.710 248.060 88.690 248.290 ;
        RECT 91.180 248.060 92.160 248.290 ;
        RECT 97.660 248.280 98.640 248.510 ;
        RECT 101.130 248.280 102.110 248.510 ;
        RECT 697.190 246.710 697.700 247.150 ;
        RECT 697.260 246.690 697.620 246.710 ;
        RECT 211.570 245.490 212.550 245.720 ;
        RECT 215.040 245.490 216.020 245.720 ;
        RECT 218.510 245.490 219.490 245.720 ;
        RECT 221.980 245.490 222.960 245.720 ;
        RECT 225.450 245.490 226.430 245.720 ;
        RECT 231.540 245.490 232.520 245.720 ;
        RECT 235.010 245.490 235.990 245.720 ;
        RECT 238.480 245.490 239.460 245.720 ;
        RECT 241.950 245.490 242.930 245.720 ;
        RECT 245.420 245.490 246.400 245.720 ;
        RECT 251.650 245.490 252.630 245.720 ;
        RECT 255.120 245.490 256.100 245.720 ;
        RECT 258.590 245.490 259.570 245.720 ;
        RECT 262.060 245.490 263.040 245.720 ;
        RECT 265.530 245.490 266.510 245.720 ;
        RECT 271.760 245.490 272.740 245.720 ;
        RECT 275.230 245.490 276.210 245.720 ;
        RECT 278.700 245.490 279.680 245.720 ;
        RECT 282.170 245.490 283.150 245.720 ;
        RECT 285.640 245.490 286.620 245.720 ;
        RECT 4.630 244.740 5.610 244.970 ;
        RECT 8.100 244.740 9.080 244.970 ;
        RECT 11.570 244.740 12.550 244.970 ;
        RECT 17.970 244.720 18.950 244.950 ;
        RECT 21.440 244.720 22.420 244.950 ;
        RECT 24.910 244.720 25.890 244.950 ;
        RECT 31.340 244.750 32.320 244.980 ;
        RECT 34.810 244.750 35.790 244.980 ;
        RECT 38.280 244.750 39.260 244.980 ;
        RECT 44.570 244.750 45.550 244.980 ;
        RECT 48.040 244.750 49.020 244.980 ;
        RECT 51.510 244.750 52.490 244.980 ;
        RECT 57.840 244.720 58.820 244.950 ;
        RECT 61.310 244.720 62.290 244.950 ;
        RECT 64.780 244.720 65.760 244.950 ;
        RECT 71.110 244.750 72.090 244.980 ;
        RECT 74.580 244.750 75.560 244.980 ;
        RECT 78.050 244.750 79.030 244.980 ;
        RECT 84.240 244.770 85.220 245.000 ;
        RECT 87.710 244.770 88.690 245.000 ;
        RECT 91.180 244.770 92.160 245.000 ;
        RECT 97.660 244.990 98.640 245.220 ;
        RECT 101.130 244.990 102.110 245.220 ;
        RECT 103.270 243.330 103.830 243.790 ;
        RECT 15.260 241.930 16.410 242.240 ;
        RECT 28.430 241.930 29.670 242.410 ;
        RECT 41.730 242.140 42.800 242.790 ;
        RECT 11.840 241.680 16.410 241.930 ;
        RECT 4.630 241.450 5.610 241.680 ;
        RECT 8.100 241.450 9.080 241.680 ;
        RECT 11.570 241.450 16.410 241.680 ;
        RECT 25.390 241.660 29.670 241.930 ;
        RECT 38.600 241.690 42.800 242.140 ;
        RECT 55.110 241.880 56.260 242.370 ;
        RECT 51.900 241.690 56.260 241.880 ;
        RECT 68.360 241.840 69.260 242.530 ;
        RECT 81.440 241.970 82.770 242.240 ;
        RECT 94.190 242.090 95.300 242.700 ;
        RECT 211.570 242.200 212.550 242.430 ;
        RECT 215.040 242.200 216.020 242.430 ;
        RECT 218.510 242.200 219.490 242.430 ;
        RECT 221.980 242.200 222.960 242.430 ;
        RECT 225.450 242.200 226.430 242.430 ;
        RECT 231.540 242.200 232.520 242.430 ;
        RECT 235.010 242.200 235.990 242.430 ;
        RECT 238.480 242.200 239.460 242.430 ;
        RECT 241.950 242.200 242.930 242.430 ;
        RECT 245.420 242.200 246.400 242.430 ;
        RECT 251.650 242.200 252.630 242.430 ;
        RECT 255.120 242.200 256.100 242.430 ;
        RECT 258.590 242.200 259.570 242.430 ;
        RECT 262.060 242.200 263.040 242.430 ;
        RECT 265.530 242.200 266.510 242.430 ;
        RECT 271.760 242.200 272.740 242.430 ;
        RECT 275.230 242.200 276.210 242.430 ;
        RECT 278.700 242.200 279.680 242.430 ;
        RECT 282.170 242.200 283.150 242.430 ;
        RECT 285.640 242.200 286.620 242.430 ;
        RECT 11.840 241.130 16.410 241.450 ;
        RECT 17.970 241.430 18.950 241.660 ;
        RECT 21.440 241.430 22.420 241.660 ;
        RECT 24.910 241.430 29.670 241.660 ;
        RECT 31.340 241.460 32.320 241.690 ;
        RECT 34.810 241.460 35.790 241.690 ;
        RECT 38.280 241.460 42.800 241.690 ;
        RECT 44.570 241.460 45.550 241.690 ;
        RECT 48.040 241.460 49.020 241.690 ;
        RECT 51.510 241.460 56.260 241.690 ;
        RECT 64.940 241.660 69.260 241.840 ;
        RECT 78.320 241.690 82.770 241.970 ;
        RECT 91.450 241.710 95.300 242.090 ;
        RECT 15.260 240.350 16.410 241.130 ;
        RECT 25.390 241.090 29.670 241.430 ;
        RECT 28.430 240.480 29.670 241.090 ;
        RECT 38.600 240.960 42.800 241.460 ;
        RECT 41.730 240.230 42.800 240.960 ;
        RECT 51.900 240.920 56.260 241.460 ;
        RECT 57.840 241.430 58.820 241.660 ;
        RECT 61.310 241.430 62.290 241.660 ;
        RECT 64.780 241.430 69.260 241.660 ;
        RECT 71.110 241.460 72.090 241.690 ;
        RECT 74.580 241.460 75.560 241.690 ;
        RECT 78.050 241.460 82.770 241.690 ;
        RECT 84.240 241.480 85.220 241.710 ;
        RECT 87.710 241.480 88.690 241.710 ;
        RECT 91.180 241.480 95.300 241.710 ;
        RECT 97.660 241.700 98.640 241.930 ;
        RECT 101.130 241.700 102.110 241.930 ;
        RECT 64.940 241.250 69.260 241.430 ;
        RECT 78.320 241.380 82.770 241.460 ;
        RECT 55.110 240.060 56.260 240.920 ;
        RECT 68.360 240.270 69.260 241.250 ;
        RECT 81.440 240.770 82.770 241.380 ;
        RECT 91.450 241.300 95.300 241.480 ;
        RECT 94.190 240.850 95.300 241.300 ;
        RECT 213.100 240.380 224.920 241.290 ;
        RECT 232.640 240.380 247.090 241.090 ;
        RECT 253.030 240.380 267.220 241.030 ;
        RECT 271.770 240.380 286.360 241.090 ;
        RECT 213.100 239.460 286.360 240.380 ;
        RECT 213.100 239.180 224.920 239.460 ;
        RECT 232.640 239.310 247.090 239.460 ;
        RECT 253.030 239.240 267.220 239.460 ;
        RECT 271.770 239.310 286.360 239.460 ;
        RECT 4.630 238.160 5.610 238.390 ;
        RECT 8.100 238.160 9.080 238.390 ;
        RECT 11.570 238.160 12.550 238.390 ;
        RECT 17.970 238.140 18.950 238.370 ;
        RECT 21.440 238.140 22.420 238.370 ;
        RECT 24.910 238.140 25.890 238.370 ;
        RECT 31.340 238.170 32.320 238.400 ;
        RECT 34.810 238.170 35.790 238.400 ;
        RECT 38.280 238.170 39.260 238.400 ;
        RECT 44.570 238.170 45.550 238.400 ;
        RECT 48.040 238.170 49.020 238.400 ;
        RECT 51.510 238.170 52.490 238.400 ;
        RECT 57.840 238.140 58.820 238.370 ;
        RECT 61.310 238.140 62.290 238.370 ;
        RECT 64.780 238.140 65.760 238.370 ;
        RECT 71.110 238.170 72.090 238.400 ;
        RECT 74.580 238.170 75.560 238.400 ;
        RECT 78.050 238.170 79.030 238.400 ;
        RECT 84.240 238.190 85.220 238.420 ;
        RECT 87.710 238.190 88.690 238.420 ;
        RECT 91.180 238.190 92.160 238.420 ;
        RECT 97.660 238.410 98.640 238.640 ;
        RECT 101.130 238.410 102.110 238.640 ;
        RECT 1.170 237.000 13.740 237.320 ;
        RECT 1.170 236.760 22.080 237.000 ;
        RECT 45.190 236.760 53.170 237.150 ;
        RECT 70.820 236.760 78.480 237.080 ;
        RECT 84.810 236.760 92.070 237.170 ;
        RECT 97.030 236.760 102.620 237.060 ;
        RECT -51.950 236.050 -51.410 236.280 ;
        RECT -50.660 236.050 -50.120 236.280 ;
        RECT -49.370 236.050 -48.830 236.280 ;
        RECT -48.080 236.050 -47.540 236.280 ;
        RECT -46.790 236.050 -46.250 236.280 ;
        RECT -45.500 236.050 -44.960 236.280 ;
        RECT -44.210 236.050 -43.670 236.280 ;
        RECT -42.920 236.050 -42.380 236.280 ;
        RECT -41.630 236.050 -41.090 236.280 ;
        RECT -40.340 236.050 -39.800 236.280 ;
        RECT -39.050 236.050 -38.510 236.280 ;
        RECT -37.760 236.050 -37.220 236.280 ;
        RECT -36.470 236.050 -35.930 236.280 ;
        RECT -35.180 236.050 -34.640 236.280 ;
        RECT -33.890 236.050 -33.350 236.280 ;
        RECT -32.600 236.050 -32.060 236.280 ;
        RECT -31.310 236.050 -30.770 236.280 ;
        RECT -30.020 236.050 -29.480 236.280 ;
        RECT -28.730 236.050 -28.190 236.280 ;
        RECT -27.440 236.050 -26.900 236.280 ;
        RECT 1.170 236.050 102.620 236.760 ;
        RECT -52.475 235.390 -52.205 235.410 ;
        RECT -44.035 235.390 -43.885 236.050 ;
        RECT 1.170 236.020 13.740 236.050 ;
        RECT 1.170 235.920 2.470 236.020 ;
        RECT 20.900 235.950 102.620 236.050 ;
        RECT 20.900 235.800 97.760 235.950 ;
        RECT -52.545 235.050 -26.295 235.390 ;
        RECT -52.475 233.930 -52.205 235.050 ;
        RECT -49.835 234.135 -49.565 235.050 ;
        RECT -52.440 232.555 -52.210 233.930 ;
        RECT -49.860 233.890 -49.565 234.135 ;
        RECT -49.860 232.555 -49.630 233.890 ;
        RECT -47.305 233.870 -47.035 235.050 ;
        RECT -47.280 232.555 -47.050 233.870 ;
        RECT -44.715 233.810 -44.445 235.050 ;
        RECT -42.135 233.810 -41.865 235.050 ;
        RECT -44.700 232.555 -44.470 233.810 ;
        RECT -42.120 232.555 -41.890 233.810 ;
        RECT -39.565 233.750 -39.295 235.050 ;
        RECT -39.540 232.555 -39.310 233.750 ;
        RECT -36.975 233.730 -36.705 235.050 ;
        RECT -34.395 233.870 -34.125 235.050 ;
        RECT -36.960 232.555 -36.730 233.730 ;
        RECT -34.380 232.555 -34.150 233.870 ;
        RECT -31.825 233.850 -31.555 235.050 ;
        RECT -29.225 233.850 -28.955 235.050 ;
        RECT -26.635 234.135 -26.365 235.050 ;
        RECT -31.800 232.555 -31.570 233.850 ;
        RECT -29.220 232.555 -28.990 233.850 ;
        RECT -26.640 233.810 -26.365 234.135 ;
        RECT -26.640 232.555 -26.410 233.810 ;
        RECT -46.070 224.520 -32.460 227.200 ;
        RECT -51.840 223.900 -51.300 224.130 ;
        RECT -50.550 223.900 -50.010 224.130 ;
        RECT -49.260 223.900 -48.720 224.130 ;
        RECT -47.970 223.900 -47.430 224.130 ;
        RECT -46.680 223.900 -46.140 224.130 ;
        RECT -45.390 223.900 -44.850 224.130 ;
        RECT -44.100 223.900 -43.560 224.130 ;
        RECT -42.810 223.900 -42.270 224.130 ;
        RECT -41.520 223.900 -40.980 224.130 ;
        RECT -40.230 223.900 -39.690 224.130 ;
        RECT -38.940 223.900 -38.400 224.130 ;
        RECT -37.650 223.900 -37.110 224.130 ;
        RECT -36.360 223.900 -35.820 224.130 ;
        RECT -35.070 223.900 -34.530 224.130 ;
        RECT -33.780 223.900 -33.240 224.130 ;
        RECT -32.490 223.900 -31.950 224.130 ;
        RECT -31.200 223.900 -30.660 224.130 ;
        RECT -29.910 223.900 -29.370 224.130 ;
        RECT -28.620 223.900 -28.080 224.130 ;
        RECT -27.330 223.900 -26.790 224.130 ;
        RECT -52.365 223.240 -52.095 223.260 ;
        RECT -43.925 223.240 -43.775 223.900 ;
        RECT -52.435 222.900 -26.185 223.240 ;
        RECT -52.365 221.780 -52.095 222.900 ;
        RECT -49.725 221.985 -49.455 222.900 ;
        RECT -52.330 220.405 -52.100 221.780 ;
        RECT -49.750 221.740 -49.455 221.985 ;
        RECT -49.750 220.405 -49.520 221.740 ;
        RECT -47.195 221.720 -46.925 222.900 ;
        RECT -47.170 220.405 -46.940 221.720 ;
        RECT -44.605 221.660 -44.335 222.900 ;
        RECT -42.025 221.660 -41.755 222.900 ;
        RECT -44.590 220.405 -44.360 221.660 ;
        RECT -42.010 220.405 -41.780 221.660 ;
        RECT -39.455 221.600 -39.185 222.900 ;
        RECT -39.430 220.405 -39.200 221.600 ;
        RECT -36.865 221.580 -36.595 222.900 ;
        RECT -34.285 221.720 -34.015 222.900 ;
        RECT -36.850 220.405 -36.620 221.580 ;
        RECT -34.270 220.405 -34.040 221.720 ;
        RECT -31.715 221.700 -31.445 222.900 ;
        RECT -29.115 221.700 -28.845 222.900 ;
        RECT -26.525 221.985 -26.255 222.900 ;
        RECT -31.690 220.405 -31.460 221.700 ;
        RECT -29.110 220.405 -28.880 221.700 ;
        RECT -26.530 221.660 -26.255 221.985 ;
        RECT -26.530 220.405 -26.300 221.660 ;
        RECT -46.070 136.910 -32.460 139.590 ;
        RECT -51.880 136.250 -51.340 136.480 ;
        RECT -50.590 136.250 -50.050 136.480 ;
        RECT -49.300 136.250 -48.760 136.480 ;
        RECT -48.010 136.250 -47.470 136.480 ;
        RECT -46.720 136.250 -46.180 136.480 ;
        RECT -45.430 136.250 -44.890 136.480 ;
        RECT -44.140 136.250 -43.600 136.480 ;
        RECT -42.850 136.250 -42.310 136.480 ;
        RECT -41.560 136.250 -41.020 136.480 ;
        RECT -40.270 136.250 -39.730 136.480 ;
        RECT -38.980 136.250 -38.440 136.480 ;
        RECT -37.690 136.250 -37.150 136.480 ;
        RECT -36.400 136.250 -35.860 136.480 ;
        RECT -35.110 136.250 -34.570 136.480 ;
        RECT -33.820 136.250 -33.280 136.480 ;
        RECT -32.530 136.250 -31.990 136.480 ;
        RECT -31.240 136.250 -30.700 136.480 ;
        RECT -29.950 136.250 -29.410 136.480 ;
        RECT -28.660 136.250 -28.120 136.480 ;
        RECT -27.370 136.250 -26.830 136.480 ;
        RECT -52.405 135.590 -52.135 135.610 ;
        RECT -43.965 135.590 -43.815 136.250 ;
        RECT -52.475 135.250 -26.225 135.590 ;
        RECT -52.405 134.130 -52.135 135.250 ;
        RECT -49.765 134.335 -49.495 135.250 ;
        RECT -52.370 132.755 -52.140 134.130 ;
        RECT -49.790 134.090 -49.495 134.335 ;
        RECT -49.790 132.755 -49.560 134.090 ;
        RECT -47.235 134.070 -46.965 135.250 ;
        RECT -47.210 132.755 -46.980 134.070 ;
        RECT -44.645 134.010 -44.375 135.250 ;
        RECT -42.065 134.010 -41.795 135.250 ;
        RECT -44.630 132.755 -44.400 134.010 ;
        RECT -42.050 132.755 -41.820 134.010 ;
        RECT -39.495 133.950 -39.225 135.250 ;
        RECT -39.470 132.755 -39.240 133.950 ;
        RECT -36.905 133.930 -36.635 135.250 ;
        RECT -34.325 134.070 -34.055 135.250 ;
        RECT -36.890 132.755 -36.660 133.930 ;
        RECT -34.310 132.755 -34.080 134.070 ;
        RECT -31.755 134.050 -31.485 135.250 ;
        RECT -29.155 134.050 -28.885 135.250 ;
        RECT -26.565 134.335 -26.295 135.250 ;
        RECT -31.730 132.755 -31.500 134.050 ;
        RECT -29.150 132.755 -28.920 134.050 ;
        RECT -26.570 134.010 -26.295 134.335 ;
        RECT -26.570 132.755 -26.340 134.010 ;
        RECT -45.950 17.470 -32.340 20.150 ;
        RECT -51.760 16.810 -51.220 17.040 ;
        RECT -50.470 16.810 -49.930 17.040 ;
        RECT -49.180 16.810 -48.640 17.040 ;
        RECT -47.890 16.810 -47.350 17.040 ;
        RECT -46.600 16.810 -46.060 17.040 ;
        RECT -45.310 16.810 -44.770 17.040 ;
        RECT -44.020 16.810 -43.480 17.040 ;
        RECT -42.730 16.810 -42.190 17.040 ;
        RECT -41.440 16.810 -40.900 17.040 ;
        RECT -40.150 16.810 -39.610 17.040 ;
        RECT -38.860 16.810 -38.320 17.040 ;
        RECT -37.570 16.810 -37.030 17.040 ;
        RECT -36.280 16.810 -35.740 17.040 ;
        RECT -34.990 16.810 -34.450 17.040 ;
        RECT -33.700 16.810 -33.160 17.040 ;
        RECT -32.410 16.810 -31.870 17.040 ;
        RECT -31.120 16.810 -30.580 17.040 ;
        RECT -29.830 16.810 -29.290 17.040 ;
        RECT -28.540 16.810 -28.000 17.040 ;
        RECT -27.250 16.810 -26.710 17.040 ;
        RECT -52.285 16.150 -52.015 16.170 ;
        RECT -43.845 16.150 -43.695 16.810 ;
        RECT -52.355 15.810 -26.105 16.150 ;
        RECT -52.285 14.690 -52.015 15.810 ;
        RECT -49.645 14.895 -49.375 15.810 ;
        RECT -52.250 13.315 -52.020 14.690 ;
        RECT -49.670 14.650 -49.375 14.895 ;
        RECT -49.670 13.315 -49.440 14.650 ;
        RECT -47.115 14.630 -46.845 15.810 ;
        RECT -47.090 13.315 -46.860 14.630 ;
        RECT -44.525 14.570 -44.255 15.810 ;
        RECT -41.945 14.570 -41.675 15.810 ;
        RECT -44.510 13.315 -44.280 14.570 ;
        RECT -41.930 13.315 -41.700 14.570 ;
        RECT -39.375 14.510 -39.105 15.810 ;
        RECT -39.350 13.315 -39.120 14.510 ;
        RECT -36.785 14.490 -36.515 15.810 ;
        RECT -34.205 14.630 -33.935 15.810 ;
        RECT -36.770 13.315 -36.540 14.490 ;
        RECT -34.190 13.315 -33.960 14.630 ;
        RECT -31.635 14.610 -31.365 15.810 ;
        RECT -29.035 14.610 -28.765 15.810 ;
        RECT -26.445 14.895 -26.175 15.810 ;
        RECT -31.610 13.315 -31.380 14.610 ;
        RECT -29.030 13.315 -28.800 14.610 ;
        RECT -26.450 14.570 -26.175 14.895 ;
        RECT -26.450 13.315 -26.220 14.570 ;
      LAYER via ;
        RECT -34.695 378.580 29.565 410.840 ;
        RECT 1086.970 380.290 1130.750 409.670 ;
        RECT -44.565 358.040 -34.385 359.580 ;
        RECT -46.065 236.720 -32.685 239.220 ;
        RECT 590.550 335.215 591.450 336.115 ;
        RECT 832.280 354.465 832.540 354.725 ;
        RECT 832.105 352.035 832.365 352.295 ;
        RECT 655.330 332.325 657.510 333.865 ;
        RECT 664.830 332.150 665.090 332.410 ;
        RECT 665.150 332.150 665.410 332.410 ;
        RECT 670.130 332.260 670.390 332.520 ;
        RECT 670.450 332.260 670.710 332.520 ;
        RECT 675.770 332.130 676.030 332.390 ;
        RECT 676.090 332.130 676.350 332.390 ;
        RECT 683.080 332.090 683.340 332.350 ;
        RECT 683.400 332.090 683.660 332.350 ;
        RECT 688.830 332.130 689.090 332.390 ;
        RECT 689.150 332.130 689.410 332.390 ;
        RECT 591.560 325.190 592.460 326.090 ;
        RECT 659.315 326.040 659.575 326.300 ;
        RECT 664.195 326.060 664.455 326.320 ;
        RECT 659.315 325.720 659.575 325.980 ;
        RECT 668.895 326.020 669.155 326.280 ;
        RECT 673.355 326.060 673.615 326.320 ;
        RECT 664.195 325.740 664.455 326.000 ;
        RECT 668.895 325.700 669.155 325.960 ;
        RECT 673.355 325.740 673.615 326.000 ;
        RECT 676.940 325.880 677.200 326.140 ;
        RECT 677.260 325.880 677.520 326.140 ;
        RECT 661.540 319.845 662.120 320.425 ;
        RECT 663.630 319.985 663.890 320.245 ;
        RECT 663.950 319.985 664.210 320.245 ;
        RECT 667.450 319.995 667.710 320.255 ;
        RECT 680.210 320.030 680.470 320.290 ;
        RECT 860.770 320.180 861.030 320.440 ;
        RECT 860.770 319.860 861.030 320.120 ;
        RECT 864.710 320.285 864.970 320.545 ;
        RECT 864.710 319.965 864.970 320.225 ;
        RECT 590.490 316.995 591.390 317.895 ;
        RECT 680.255 314.675 680.515 314.935 ;
        RECT 679.995 299.110 680.575 299.690 ;
        RECT 590.590 297.835 591.490 298.735 ;
        RECT 858.345 298.045 858.605 298.305 ;
        RECT 819.530 292.640 819.790 292.900 ;
        RECT 863.780 294.115 864.040 294.375 ;
        RECT 858.415 292.865 858.675 293.125 ;
        RECT 841.460 290.995 841.720 291.255 ;
        RECT 819.495 288.240 819.755 288.500 ;
        RECT 858.500 287.730 858.760 287.990 ;
        RECT 858.500 287.410 858.760 287.670 ;
        RECT 856.140 287.075 856.400 287.335 ;
        RECT 856.460 287.075 856.720 287.335 ;
        RECT 863.810 285.145 864.070 285.405 ;
        RECT 800.165 283.190 800.425 283.450 ;
        RECT 819.560 283.290 819.820 283.550 ;
        RECT 828.240 283.385 828.500 283.645 ;
        RECT 828.240 283.065 828.500 283.325 ;
        RECT 841.920 283.135 842.180 283.395 ;
        RECT 679.950 281.915 680.210 282.175 ;
        RECT 590.060 279.295 590.960 280.195 ;
        RECT 710.290 282.275 710.550 282.535 ;
        RECT 710.290 281.955 710.550 282.215 ;
        RECT 842.995 282.570 843.575 283.150 ;
        RECT 858.500 282.320 858.760 282.580 ;
        RECT 858.500 282.000 858.760 282.260 ;
        RECT 756.550 280.285 756.810 280.545 ;
        RECT 756.550 279.965 756.810 280.225 ;
        RECT 710.520 277.025 710.780 277.285 ;
        RECT 710.520 276.705 710.780 276.965 ;
        RECT 682.600 276.425 682.860 276.685 ;
        RECT 682.600 276.105 682.860 276.365 ;
        RECT 699.830 276.445 700.090 276.705 ;
        RECT 699.830 276.125 700.090 276.385 ;
        RECT 717.400 276.545 717.660 276.805 ;
        RECT 717.400 276.225 717.660 276.485 ;
        RECT 734.570 276.575 734.830 276.835 ;
        RECT 734.570 276.255 734.830 276.515 ;
        RECT 752.380 276.635 752.640 276.895 ;
        RECT 752.380 276.315 752.640 276.575 ;
        RECT 761.610 276.620 761.870 276.880 ;
        RECT 761.610 276.300 761.870 276.560 ;
        RECT 778.730 275.410 779.310 276.950 ;
        RECT 800.205 275.560 800.465 275.820 ;
        RECT 756.465 274.090 756.725 274.350 ;
        RECT 756.465 273.770 756.725 274.030 ;
        RECT 682.310 270.755 682.570 271.015 ;
        RECT 682.310 270.435 682.570 270.695 ;
        RECT 699.540 270.775 699.800 271.035 ;
        RECT 699.540 270.455 699.800 270.715 ;
        RECT 717.110 270.875 717.370 271.135 ;
        RECT 717.110 270.555 717.370 270.815 ;
        RECT 734.280 270.905 734.540 271.165 ;
        RECT 734.280 270.585 734.540 270.845 ;
        RECT 752.090 270.965 752.350 271.225 ;
        RECT 752.090 270.645 752.350 270.905 ;
        RECT 756.510 268.380 756.770 268.640 ;
        RECT 756.510 268.060 756.770 268.320 ;
        RECT 589.960 261.635 590.860 262.535 ;
        RECT 710.270 260.745 710.530 261.005 ;
        RECT 841.575 275.010 842.155 275.590 ;
        RECT 843.010 275.585 843.270 275.845 ;
        RECT 843.330 275.585 843.590 275.845 ;
        RECT 858.560 275.780 858.820 276.040 ;
        RECT 858.560 275.460 858.820 275.720 ;
        RECT 863.635 271.695 864.215 272.275 ;
        RECT 841.485 270.045 841.745 270.305 ;
        RECT 858.720 269.070 858.980 269.330 ;
        RECT 858.720 268.750 858.980 269.010 ;
        RECT 710.270 260.425 710.530 260.685 ;
        RECT 858.540 259.780 858.800 260.040 ;
        RECT 858.540 259.460 858.800 259.720 ;
        RECT 863.615 256.570 864.195 257.150 ;
        RECT 710.500 255.495 710.760 255.755 ;
        RECT 710.500 255.175 710.760 255.435 ;
        RECT 682.580 254.895 682.840 255.155 ;
        RECT 682.580 254.575 682.840 254.835 ;
        RECT 699.810 254.915 700.070 255.175 ;
        RECT 699.810 254.595 700.070 254.855 ;
        RECT 717.380 255.015 717.640 255.275 ;
        RECT 717.380 254.695 717.640 254.955 ;
        RECT 734.550 255.045 734.810 255.305 ;
        RECT 734.550 254.725 734.810 254.985 ;
        RECT 752.360 255.105 752.620 255.365 ;
        RECT 752.360 254.785 752.620 255.045 ;
        RECT 858.630 254.000 858.890 254.260 ;
        RECT 858.630 253.680 858.890 253.940 ;
        RECT 697.150 253.000 697.410 253.260 ;
        RECT 682.290 249.225 682.550 249.485 ;
        RECT 682.290 248.905 682.550 249.165 ;
        RECT 699.520 249.245 699.780 249.505 ;
        RECT 699.520 248.925 699.780 249.185 ;
        RECT 717.090 249.345 717.350 249.605 ;
        RECT 717.090 249.025 717.350 249.285 ;
        RECT 734.260 249.375 734.520 249.635 ;
        RECT 734.260 249.055 734.520 249.315 ;
        RECT 752.070 249.435 752.330 249.695 ;
        RECT 752.070 249.115 752.330 249.375 ;
        RECT 697.315 246.800 697.575 247.060 ;
        RECT -45.955 224.610 -32.575 227.110 ;
        RECT -45.955 137.000 -32.575 139.500 ;
        RECT -45.835 17.560 -32.455 20.060 ;
      LAYER met2 ;
        RECT -34.700 378.420 29.570 411.000 ;
        RECT 1086.970 380.100 1130.750 409.860 ;
        RECT -44.590 357.940 -34.360 359.680 ;
        RECT 832.160 354.320 832.660 354.870 ;
        RECT 832.160 352.400 832.350 354.320 ;
        RECT 832.070 351.930 832.400 352.400 ;
        RECT 590.500 336.130 591.500 336.320 ;
        RECT 589.990 335.010 591.500 336.130 ;
        RECT 589.990 326.040 590.700 335.010 ;
        RECT 655.320 332.620 657.520 333.980 ;
        RECT 655.320 332.610 665.250 332.620 ;
        RECT 655.320 332.420 665.440 332.610 ;
        RECT 670.100 332.420 670.740 332.720 ;
        RECT 675.740 332.420 676.380 332.590 ;
        RECT 683.050 332.420 683.690 332.550 ;
        RECT 688.800 332.420 689.440 332.590 ;
        RECT 655.320 332.290 689.440 332.420 ;
        RECT 655.320 332.210 657.520 332.290 ;
        RECT 591.430 326.040 592.590 326.230 ;
        RECT 589.990 325.570 592.590 326.040 ;
        RECT 589.990 319.940 590.700 325.570 ;
        RECT 591.430 325.050 592.590 325.570 ;
        RECT 656.060 326.150 656.570 332.210 ;
        RECT 664.800 332.130 689.440 332.290 ;
        RECT 664.800 331.950 665.440 332.130 ;
        RECT 670.100 332.060 670.740 332.130 ;
        RECT 675.740 331.930 676.380 332.130 ;
        RECT 683.050 331.890 683.690 332.130 ;
        RECT 688.800 331.930 689.440 332.130 ;
        RECT 659.260 326.150 659.630 326.370 ;
        RECT 656.060 326.090 659.630 326.150 ;
        RECT 664.140 326.090 664.510 326.390 ;
        RECT 668.840 326.090 669.210 326.350 ;
        RECT 673.300 326.090 673.670 326.390 ;
        RECT 656.060 325.990 673.670 326.090 ;
        RECT 676.890 325.990 677.570 326.330 ;
        RECT 656.060 325.810 677.570 325.990 ;
        RECT 656.060 320.710 656.490 325.810 ;
        RECT 659.260 325.740 677.570 325.810 ;
        RECT 659.260 325.650 659.630 325.740 ;
        RECT 664.140 325.670 664.510 325.740 ;
        RECT 668.840 325.630 669.210 325.740 ;
        RECT 673.300 325.700 677.570 325.740 ;
        RECT 673.300 325.670 673.670 325.700 ;
        RECT 676.890 325.690 677.570 325.700 ;
        RECT 656.060 320.240 656.530 320.710 ;
        RECT 661.450 320.280 662.210 320.490 ;
        RECT 659.050 320.240 662.210 320.280 ;
        RECT 589.970 319.590 590.710 319.940 ;
        RECT 656.060 319.790 662.210 320.240 ;
        RECT 656.060 319.750 658.700 319.790 ;
        RECT 661.450 319.780 662.210 319.790 ;
        RECT 663.590 320.300 664.250 320.450 ;
        RECT 667.300 320.300 667.860 320.410 ;
        RECT 663.590 320.050 667.860 320.300 ;
        RECT 663.590 319.780 664.250 320.050 ;
        RECT 667.300 319.840 667.860 320.050 ;
        RECT 680.150 319.830 680.530 320.490 ;
        RECT 860.660 320.330 861.140 320.570 ;
        RECT 864.670 320.330 865.010 320.640 ;
        RECT 860.660 320.100 865.010 320.330 ;
        RECT 860.660 319.730 861.140 320.100 ;
        RECT 864.670 319.870 865.010 320.100 ;
        RECT 589.990 318.100 590.700 319.590 ;
        RECT 589.990 316.790 591.440 318.100 ;
        RECT 589.990 300.710 590.700 316.790 ;
        RECT 680.100 314.530 680.670 315.080 ;
        RECT 589.990 299.970 590.650 300.710 ;
        RECT 589.990 298.940 590.700 299.970 ;
        RECT 679.860 299.050 680.710 299.750 ;
        RECT 589.990 297.630 591.540 298.940 ;
        RECT 589.990 280.400 590.700 297.630 ;
        RECT 679.880 296.060 680.200 299.050 ;
        RECT 858.310 297.870 858.640 298.480 ;
        RECT 679.880 294.490 680.190 296.060 ;
        RECT 679.880 282.370 680.200 294.490 ;
        RECT 858.430 293.300 858.580 297.870 ;
        RECT 863.730 293.990 864.090 294.500 ;
        RECT 819.510 292.460 819.810 293.080 ;
        RECT 858.380 292.690 858.710 293.300 ;
        RECT 819.560 288.660 819.700 292.460 ;
        RECT 841.360 290.790 841.830 291.440 ;
        RECT 819.450 288.080 819.800 288.660 ;
        RECT 819.600 283.730 819.780 288.080 ;
        RECT 858.440 288.060 858.590 292.690 ;
        RECT 856.130 286.870 856.730 287.540 ;
        RECT 858.400 287.340 858.860 288.060 ;
        RECT 819.540 283.610 819.840 283.730 ;
        RECT 828.170 283.610 828.570 283.710 ;
        RECT 800.090 283.030 800.500 283.610 ;
        RECT 819.540 283.450 828.570 283.610 ;
        RECT 819.540 283.110 819.840 283.450 ;
        RECT 679.810 281.720 680.350 282.370 ;
        RECT 710.170 281.840 710.670 282.650 ;
        RECT 589.990 279.090 591.010 280.400 ;
        RECT 589.990 262.740 590.700 279.090 ;
        RECT 710.380 277.400 710.570 281.840 ;
        RECT 756.400 279.900 756.960 280.610 ;
        RECT 756.470 279.770 756.710 279.900 ;
        RECT 710.380 277.130 710.900 277.400 ;
        RECT 682.540 276.500 682.920 276.740 ;
        RECT 699.770 276.520 700.150 276.760 ;
        RECT 710.400 276.590 710.900 277.130 ;
        RECT 717.340 276.620 717.720 276.860 ;
        RECT 734.510 276.650 734.890 276.890 ;
        RECT 752.320 276.710 752.700 276.950 ;
        RECT 682.380 276.050 682.920 276.500 ;
        RECT 699.610 276.070 700.150 276.520 ;
        RECT 717.180 276.170 717.720 276.620 ;
        RECT 734.350 276.200 734.890 276.650 ;
        RECT 752.160 276.260 752.700 276.710 ;
        RECT 682.380 271.070 682.680 276.050 ;
        RECT 699.610 271.090 699.910 276.070 ;
        RECT 717.180 271.190 717.480 276.170 ;
        RECT 734.350 271.220 734.650 276.200 ;
        RECT 752.160 271.280 752.460 276.260 ;
        RECT 756.470 274.520 756.690 279.770 ;
        RECT 761.500 276.710 761.980 276.950 ;
        RECT 778.600 276.710 779.440 277.140 ;
        RECT 761.500 276.400 779.440 276.710 ;
        RECT 761.500 276.230 761.980 276.400 ;
        RECT 778.600 275.220 779.440 276.400 ;
        RECT 800.180 275.980 800.370 283.030 ;
        RECT 828.170 283.000 828.570 283.450 ;
        RECT 841.830 283.230 842.300 283.590 ;
        RECT 841.680 282.940 842.300 283.230 ;
        RECT 841.680 282.400 841.980 282.940 ;
        RECT 842.970 282.490 843.600 283.230 ;
        RECT 858.510 282.650 858.650 287.340 ;
        RECT 863.830 285.530 863.980 293.990 ;
        RECT 863.760 285.230 864.120 285.530 ;
        RECT 863.750 285.020 864.120 285.230 ;
        RECT 843.090 276.030 843.330 282.490 ;
        RECT 858.400 281.930 858.860 282.650 ;
        RECT 858.550 276.110 858.740 281.930 ;
        RECT 800.130 275.400 800.540 275.980 ;
        RECT 841.550 274.930 842.180 275.670 ;
        RECT 842.980 275.400 843.620 276.030 ;
        RECT 858.460 275.390 858.920 276.110 ;
        RECT 756.350 273.600 756.840 274.520 ;
        RECT 682.250 270.750 682.680 271.070 ;
        RECT 699.480 270.770 699.910 271.090 ;
        RECT 717.050 270.870 717.480 271.190 ;
        RECT 734.220 270.900 734.650 271.220 ;
        RECT 752.030 270.960 752.460 271.280 ;
        RECT 682.250 270.380 682.630 270.750 ;
        RECT 699.480 270.400 699.860 270.770 ;
        RECT 717.050 270.500 717.430 270.870 ;
        RECT 734.220 270.530 734.600 270.900 ;
        RECT 752.030 270.590 752.410 270.960 ;
        RECT 756.510 268.690 756.680 273.600 ;
        RECT 841.610 270.510 841.800 274.930 ;
        RECT 841.420 269.840 841.810 270.510 ;
        RECT 858.710 269.400 858.910 275.390 ;
        RECT 863.750 272.430 863.920 285.020 ;
        RECT 863.550 271.540 864.300 272.430 ;
        RECT 858.620 268.850 859.080 269.400 ;
        RECT 756.460 268.010 756.820 268.690 ;
        RECT 858.580 268.680 859.080 268.850 ;
        RECT 589.910 261.430 590.910 262.740 ;
        RECT 710.150 260.310 710.650 261.120 ;
        RECT 710.360 255.870 710.550 260.310 ;
        RECT 858.580 260.110 858.800 268.680 ;
        RECT 858.440 259.390 858.900 260.110 ;
        RECT 710.360 255.600 710.880 255.870 ;
        RECT 682.520 254.970 682.900 255.210 ;
        RECT 699.750 254.990 700.130 255.230 ;
        RECT 710.380 255.060 710.880 255.600 ;
        RECT 717.320 255.090 717.700 255.330 ;
        RECT 734.490 255.120 734.870 255.360 ;
        RECT 752.300 255.180 752.680 255.420 ;
        RECT 682.360 254.520 682.900 254.970 ;
        RECT 699.590 254.540 700.130 254.990 ;
        RECT 717.160 254.640 717.700 255.090 ;
        RECT 734.330 254.670 734.870 255.120 ;
        RECT 752.140 254.730 752.680 255.180 ;
        RECT 682.360 249.540 682.660 254.520 ;
        RECT 697.050 252.830 697.510 253.430 ;
        RECT 682.230 249.220 682.660 249.540 ;
        RECT 682.230 248.850 682.610 249.220 ;
        RECT 697.300 247.200 697.480 252.830 ;
        RECT 699.590 249.560 699.890 254.540 ;
        RECT 717.160 249.660 717.460 254.640 ;
        RECT 734.330 249.690 734.630 254.670 ;
        RECT 752.140 249.750 752.440 254.730 ;
        RECT 858.640 254.330 858.820 259.390 ;
        RECT 863.730 257.320 863.920 271.540 ;
        RECT 863.600 256.400 864.210 257.320 ;
        RECT 858.530 253.610 858.990 254.330 ;
        RECT 699.460 249.240 699.890 249.560 ;
        RECT 717.030 249.340 717.460 249.660 ;
        RECT 734.200 249.370 734.630 249.690 ;
        RECT 752.010 249.430 752.440 249.750 ;
        RECT 699.460 248.870 699.840 249.240 ;
        RECT 717.030 248.970 717.410 249.340 ;
        RECT 734.200 249.000 734.580 249.370 ;
        RECT 752.010 249.060 752.390 249.430 ;
        RECT 697.240 246.660 697.650 247.200 ;
        RECT -46.120 236.610 -32.630 239.330 ;
        RECT -46.010 224.500 -32.520 227.220 ;
        RECT -46.010 136.890 -32.520 139.610 ;
        RECT -45.890 17.450 -32.400 20.170 ;
      LAYER via2 ;
        RECT -34.505 378.570 29.375 410.850 ;
        RECT 1087.120 380.240 1130.600 409.720 ;
        RECT -44.415 358.070 -34.535 359.550 ;
        RECT 680.200 319.915 680.480 320.195 ;
        RECT 680.245 314.665 680.525 314.945 ;
        RECT 841.455 290.975 841.735 291.255 ;
        RECT 856.290 287.065 856.570 287.345 ;
        RECT 841.925 283.125 842.205 283.405 ;
        RECT -46.115 236.830 -32.635 239.110 ;
        RECT -46.005 224.720 -32.525 227.000 ;
        RECT -46.005 137.110 -32.525 139.390 ;
        RECT -45.885 17.670 -32.405 19.950 ;
      LAYER met3 ;
        RECT -34.750 378.445 29.620 410.975 ;
        RECT 1086.920 380.125 1130.800 409.835 ;
        RECT -44.640 357.965 -34.310 359.655 ;
        RECT 680.100 319.855 680.580 320.255 ;
        RECT 680.220 315.055 680.540 319.855 ;
        RECT 680.050 314.555 680.720 315.055 ;
        RECT 841.310 291.160 841.880 291.415 ;
        RECT 841.310 291.150 841.940 291.160 ;
        RECT 841.310 290.815 841.990 291.150 ;
        RECT 841.660 287.020 841.990 290.815 ;
        RECT 856.080 287.020 856.780 287.515 ;
        RECT 841.660 286.895 856.780 287.020 ;
        RECT 841.660 286.720 856.390 286.895 ;
        RECT 841.660 283.565 841.990 286.720 ;
        RECT 841.660 283.260 842.350 283.565 ;
        RECT 841.780 282.965 842.350 283.260 ;
        RECT -46.170 236.635 -32.580 239.305 ;
        RECT -46.060 224.525 -32.470 227.195 ;
        RECT -46.060 136.915 -32.470 139.585 ;
        RECT -45.940 17.475 -32.350 20.145 ;
        RECT 1072.580 -61.270 1105.690 -61.180 ;
        RECT 934.600 -61.450 1105.690 -61.270 ;
        RECT -34.820 -62.090 1105.690 -61.450 ;
        RECT -52.790 -62.460 1105.690 -62.090 ;
        RECT -52.790 -104.330 1129.420 -62.460 ;
        RECT -34.820 -104.700 1129.420 -104.330 ;
        RECT -34.820 -105.480 1105.690 -104.700 ;
        RECT -34.820 -106.250 944.550 -105.480 ;
        RECT 1072.580 -105.980 1105.690 -105.480 ;
      LAYER via3 ;
        RECT -34.525 378.550 29.395 410.870 ;
        RECT 1087.100 380.220 1130.620 409.740 ;
        RECT -44.435 358.050 -34.515 359.570 ;
        RECT -45.935 236.810 -32.815 239.130 ;
        RECT -45.825 224.700 -32.705 227.020 ;
        RECT -45.825 137.090 -32.705 139.410 ;
        RECT -45.705 17.650 -32.585 19.970 ;
        RECT -52.620 -104.170 -5.500 -62.250 ;
        RECT 1082.130 -104.540 1129.250 -62.620 ;
      LAYER met4 ;
        RECT 11.030 426.930 20.610 490.310 ;
        RECT 10.840 410.955 20.640 426.930 ;
        RECT -34.705 408.930 29.575 410.955 ;
        RECT 1088.880 409.815 1128.580 409.970 ;
        RECT -53.610 408.590 -53.310 408.620 ;
        RECT -47.450 408.590 29.575 408.930 ;
        RECT -53.610 378.465 29.575 408.590 ;
        RECT 1086.965 380.145 1130.755 409.815 ;
        RECT -53.610 374.400 -23.520 378.465 ;
        RECT -53.610 9.460 -23.530 374.400 ;
        RECT -53.630 9.220 -23.530 9.460 ;
        RECT -53.630 9.150 -23.540 9.220 ;
        RECT -53.610 -6.700 -23.540 9.150 ;
        RECT -53.610 -62.085 -23.530 -6.700 ;
        RECT 1104.390 -13.410 1128.260 380.145 ;
        RECT -53.610 -71.230 -5.375 -62.085 ;
        RECT 1104.100 -62.230 1128.540 -13.410 ;
        RECT 1086.510 -62.455 1128.540 -62.230 ;
        RECT -53.880 -104.335 -5.375 -71.230 ;
        RECT -53.880 -105.480 -10.040 -104.335 ;
        RECT 1082.005 -104.705 1129.375 -62.455 ;
    END
  END vdda2
  PIN re
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 28.980000 ;
    PORT
      LAYER li1 ;
        RECT 664.450 352.675 666.305 352.845 ;
        RECT 661.125 352.115 661.455 352.505 ;
        RECT 664.450 352.145 664.620 352.675 ;
        RECT 669.675 352.470 670.215 353.340 ;
        RECT 682.500 352.635 684.355 352.805 ;
        RECT 665.820 352.145 666.180 352.150 ;
        RECT 661.125 351.945 662.130 352.115 ;
        RECT 661.960 351.285 662.130 351.945 ;
        RECT 664.450 351.975 667.070 352.145 ;
        RECT 664.450 351.285 664.620 351.975 ;
        RECT 665.820 351.970 666.180 351.975 ;
        RECT 666.900 351.480 667.070 351.975 ;
        RECT 669.675 351.480 669.845 352.470 ;
        RECT 679.175 352.075 679.505 352.465 ;
        RECT 682.500 352.105 682.670 352.635 ;
        RECT 687.725 352.430 688.265 353.300 ;
        RECT 700.090 352.655 701.945 352.825 ;
        RECT 679.175 351.905 680.180 352.075 ;
        RECT 666.900 351.310 669.845 351.480 ;
        RECT 661.960 351.115 664.620 351.285 ;
        RECT 680.010 351.245 680.180 351.905 ;
        RECT 682.500 351.935 685.120 352.105 ;
        RECT 682.500 351.245 682.670 351.935 ;
        RECT 684.060 351.900 684.340 351.935 ;
        RECT 684.950 351.440 685.120 351.935 ;
        RECT 687.725 351.440 687.895 352.430 ;
        RECT 696.765 352.095 697.095 352.485 ;
        RECT 700.090 352.125 700.260 352.655 ;
        RECT 705.315 352.450 705.855 353.320 ;
        RECT 717.940 352.655 719.795 352.825 ;
        RECT 696.765 351.925 697.770 352.095 ;
        RECT 684.950 351.270 687.895 351.440 ;
        RECT 680.010 351.075 682.670 351.245 ;
        RECT 697.600 351.265 697.770 351.925 ;
        RECT 700.090 351.955 702.710 352.125 ;
        RECT 700.090 351.265 700.260 351.955 ;
        RECT 701.730 351.900 702.070 351.955 ;
        RECT 702.540 351.460 702.710 351.955 ;
        RECT 705.315 351.460 705.485 352.450 ;
        RECT 714.615 352.095 714.945 352.485 ;
        RECT 717.940 352.125 718.110 352.655 ;
        RECT 723.165 352.450 723.705 353.320 ;
        RECT 736.200 352.655 738.055 352.825 ;
        RECT 714.615 351.925 715.620 352.095 ;
        RECT 702.540 351.290 705.485 351.460 ;
        RECT 697.600 351.095 700.260 351.265 ;
        RECT 715.450 351.265 715.620 351.925 ;
        RECT 717.940 351.955 720.560 352.125 ;
        RECT 717.940 351.265 718.110 351.955 ;
        RECT 719.720 351.880 720.040 351.955 ;
        RECT 720.390 351.460 720.560 351.955 ;
        RECT 723.165 351.460 723.335 352.450 ;
        RECT 732.875 352.095 733.205 352.485 ;
        RECT 736.200 352.125 736.370 352.655 ;
        RECT 741.425 352.450 741.965 353.320 ;
        RECT 753.970 352.625 755.825 352.795 ;
        RECT 732.875 351.925 733.880 352.095 ;
        RECT 720.390 351.290 723.335 351.460 ;
        RECT 715.450 351.095 718.110 351.265 ;
        RECT 733.710 351.265 733.880 351.925 ;
        RECT 736.200 351.955 738.820 352.125 ;
        RECT 736.200 351.265 736.370 351.955 ;
        RECT 737.840 351.840 738.150 351.955 ;
        RECT 738.650 351.460 738.820 351.955 ;
        RECT 741.425 351.460 741.595 352.450 ;
        RECT 750.645 352.065 750.975 352.455 ;
        RECT 753.970 352.095 754.140 352.625 ;
        RECT 759.195 352.420 759.735 353.290 ;
        RECT 772.010 352.545 773.865 352.715 ;
        RECT 750.645 351.895 751.650 352.065 ;
        RECT 738.650 351.290 741.595 351.460 ;
        RECT 733.710 351.095 736.370 351.265 ;
        RECT 751.480 351.235 751.650 351.895 ;
        RECT 753.970 351.925 756.590 352.095 ;
        RECT 753.970 351.235 754.140 351.925 ;
        RECT 755.670 351.810 755.940 351.925 ;
        RECT 756.420 351.430 756.590 351.925 ;
        RECT 759.195 351.430 759.365 352.420 ;
        RECT 768.685 351.985 769.015 352.375 ;
        RECT 772.010 352.015 772.180 352.545 ;
        RECT 777.235 352.340 777.775 353.210 ;
        RECT 790.170 352.585 792.025 352.755 ;
        RECT 768.685 351.815 769.690 351.985 ;
        RECT 756.420 351.260 759.365 351.430 ;
        RECT 751.480 351.065 754.140 351.235 ;
        RECT 769.520 351.155 769.690 351.815 ;
        RECT 772.010 351.845 774.630 352.015 ;
        RECT 772.010 351.155 772.180 351.845 ;
        RECT 773.670 351.700 773.990 351.845 ;
        RECT 774.460 351.350 774.630 351.845 ;
        RECT 777.235 351.350 777.405 352.340 ;
        RECT 786.845 352.025 787.175 352.415 ;
        RECT 790.170 352.055 790.340 352.585 ;
        RECT 795.395 352.380 795.935 353.250 ;
        RECT 808.550 352.595 810.405 352.765 ;
        RECT 786.845 351.855 787.850 352.025 ;
        RECT 774.460 351.180 777.405 351.350 ;
        RECT 787.680 351.195 787.850 351.855 ;
        RECT 790.170 351.885 792.790 352.055 ;
        RECT 790.170 351.195 790.340 351.885 ;
        RECT 791.820 351.800 792.170 351.885 ;
        RECT 792.620 351.390 792.790 351.885 ;
        RECT 795.395 351.390 795.565 352.380 ;
        RECT 805.225 352.035 805.555 352.425 ;
        RECT 808.550 352.065 808.720 352.595 ;
        RECT 813.775 352.390 814.315 353.260 ;
        RECT 805.225 351.865 806.230 352.035 ;
        RECT 792.620 351.220 795.565 351.390 ;
        RECT 769.520 350.985 772.180 351.155 ;
        RECT 787.680 351.025 790.340 351.195 ;
        RECT 806.060 351.205 806.230 351.865 ;
        RECT 808.550 351.895 811.170 352.065 ;
        RECT 808.550 351.205 808.720 351.895 ;
        RECT 810.150 351.800 810.500 351.895 ;
        RECT 811.000 351.400 811.170 351.895 ;
        RECT 813.775 351.400 813.945 352.390 ;
        RECT 811.000 351.230 813.945 351.400 ;
        RECT 806.060 351.035 808.720 351.205 ;
        RECT 800.750 344.505 802.605 344.675 ;
        RECT 797.425 343.945 797.755 344.335 ;
        RECT 800.750 343.975 800.920 344.505 ;
        RECT 805.975 344.300 806.515 345.170 ;
        RECT 820.110 344.415 821.965 344.585 ;
        RECT 797.425 343.775 798.430 343.945 ;
        RECT 798.260 343.115 798.430 343.775 ;
        RECT 800.750 343.805 803.370 343.975 ;
        RECT 800.750 343.115 800.920 343.805 ;
        RECT 802.410 343.600 802.810 343.805 ;
        RECT 803.200 343.310 803.370 343.805 ;
        RECT 805.975 343.310 806.145 344.300 ;
        RECT 816.785 343.855 817.115 344.245 ;
        RECT 820.110 343.885 820.280 344.415 ;
        RECT 825.335 344.210 825.875 345.080 ;
        RECT 816.785 343.685 817.790 343.855 ;
        RECT 803.200 343.140 806.145 343.310 ;
        RECT 798.260 342.945 800.920 343.115 ;
        RECT 817.620 343.025 817.790 343.685 ;
        RECT 820.110 343.715 822.730 343.885 ;
        RECT 820.110 343.025 820.280 343.715 ;
        RECT 821.750 343.540 822.130 343.715 ;
        RECT 822.560 343.220 822.730 343.715 ;
        RECT 825.335 343.220 825.505 344.210 ;
        RECT 822.560 343.050 825.505 343.220 ;
        RECT 817.620 342.855 820.280 343.025 ;
        RECT 799.175 305.650 799.715 306.520 ;
        RECT 803.085 305.855 804.940 306.025 ;
        RECT 799.545 304.660 799.715 305.650 ;
        RECT 804.770 305.325 804.940 305.855 ;
        RECT 802.320 305.155 804.940 305.325 ;
        RECT 807.935 305.295 808.265 305.685 ;
        RECT 816.935 305.650 817.475 306.520 ;
        RECT 820.845 305.855 822.700 306.025 ;
        RECT 802.320 304.660 802.490 305.155 ;
        RECT 802.820 305.050 803.140 305.155 ;
        RECT 799.545 304.490 802.490 304.660 ;
        RECT 804.770 304.465 804.940 305.155 ;
        RECT 807.260 305.125 808.265 305.295 ;
        RECT 807.260 304.465 807.430 305.125 ;
        RECT 817.305 304.660 817.475 305.650 ;
        RECT 822.530 305.325 822.700 305.855 ;
        RECT 820.080 305.155 822.700 305.325 ;
        RECT 825.695 305.295 826.025 305.685 ;
        RECT 820.080 304.660 820.250 305.155 ;
        RECT 820.660 305.050 820.980 305.155 ;
        RECT 817.305 304.490 820.250 304.660 ;
        RECT 804.770 304.295 807.430 304.465 ;
        RECT 822.530 304.465 822.700 305.155 ;
        RECT 825.020 305.125 826.025 305.295 ;
        RECT 825.020 304.465 825.190 305.125 ;
        RECT 822.530 304.295 825.190 304.465 ;
        RECT 682.755 296.590 683.295 297.460 ;
        RECT 686.665 296.795 688.520 296.965 ;
        RECT 683.125 295.600 683.295 296.590 ;
        RECT 688.350 296.265 688.520 296.795 ;
        RECT 685.900 296.095 688.520 296.265 ;
        RECT 691.515 296.235 691.845 296.625 ;
        RECT 700.245 296.550 700.785 297.420 ;
        RECT 704.155 296.755 706.010 296.925 ;
        RECT 685.900 295.600 686.070 296.095 ;
        RECT 683.125 295.430 686.070 295.600 ;
        RECT 688.350 295.405 688.520 296.095 ;
        RECT 690.840 296.065 691.845 296.235 ;
        RECT 690.840 295.405 691.010 296.065 ;
        RECT 688.350 295.235 691.010 295.405 ;
        RECT 700.615 295.560 700.785 296.550 ;
        RECT 705.840 296.225 706.010 296.755 ;
        RECT 717.855 296.610 718.395 297.480 ;
        RECT 721.765 296.815 723.620 296.985 ;
        RECT 703.390 296.055 706.010 296.225 ;
        RECT 709.005 296.195 709.335 296.585 ;
        RECT 703.390 295.560 703.560 296.055 ;
        RECT 700.615 295.390 703.560 295.560 ;
        RECT 705.840 295.365 706.010 296.055 ;
        RECT 708.330 296.025 709.335 296.195 ;
        RECT 708.330 295.365 708.500 296.025 ;
        RECT 718.225 295.620 718.395 296.610 ;
        RECT 723.450 296.285 723.620 296.815 ;
        RECT 721.000 296.115 723.620 296.285 ;
        RECT 726.615 296.255 726.945 296.645 ;
        RECT 735.555 296.560 736.095 297.430 ;
        RECT 739.465 296.765 741.320 296.935 ;
        RECT 721.000 295.620 721.170 296.115 ;
        RECT 718.225 295.450 721.170 295.620 ;
        RECT 705.840 295.195 708.500 295.365 ;
        RECT 723.450 295.425 723.620 296.115 ;
        RECT 725.940 296.085 726.945 296.255 ;
        RECT 725.940 295.425 726.110 296.085 ;
        RECT 723.450 295.255 726.110 295.425 ;
        RECT 735.925 295.570 736.095 296.560 ;
        RECT 741.150 296.235 741.320 296.765 ;
        RECT 738.700 296.065 741.320 296.235 ;
        RECT 744.315 296.205 744.645 296.595 ;
        RECT 753.295 296.550 753.835 297.420 ;
        RECT 757.205 296.755 759.060 296.925 ;
        RECT 738.700 296.020 738.870 296.065 ;
        RECT 738.690 295.770 738.870 296.020 ;
        RECT 738.700 295.570 738.870 295.770 ;
        RECT 735.925 295.400 738.870 295.570 ;
        RECT 741.150 295.375 741.320 296.065 ;
        RECT 743.640 296.035 744.645 296.205 ;
        RECT 743.640 295.375 743.810 296.035 ;
        RECT 753.665 295.560 753.835 296.550 ;
        RECT 758.890 296.225 759.060 296.755 ;
        RECT 756.440 296.055 759.060 296.225 ;
        RECT 762.055 296.195 762.385 296.585 ;
        RECT 756.440 295.790 756.650 296.055 ;
        RECT 756.440 295.560 756.610 295.790 ;
        RECT 753.665 295.390 756.610 295.560 ;
        RECT 741.150 295.205 743.810 295.375 ;
        RECT 758.890 295.365 759.060 296.055 ;
        RECT 761.380 296.025 762.385 296.195 ;
        RECT 761.380 295.365 761.550 296.025 ;
        RECT 758.890 295.195 761.550 295.365 ;
        RECT 783.655 273.030 784.195 273.900 ;
        RECT 787.565 273.235 789.420 273.405 ;
        RECT 784.025 272.040 784.195 273.030 ;
        RECT 789.250 272.705 789.420 273.235 ;
        RECT 786.800 272.535 789.420 272.705 ;
        RECT 792.415 272.675 792.745 273.065 ;
        RECT 802.545 273.020 803.085 273.890 ;
        RECT 806.455 273.225 808.310 273.395 ;
        RECT 786.800 272.040 786.970 272.535 ;
        RECT 787.380 272.360 787.860 272.535 ;
        RECT 784.025 271.870 786.970 272.040 ;
        RECT 789.250 271.845 789.420 272.535 ;
        RECT 791.740 272.505 792.745 272.675 ;
        RECT 791.740 271.845 791.910 272.505 ;
        RECT 802.915 272.030 803.085 273.020 ;
        RECT 808.140 272.695 808.310 273.225 ;
        RECT 805.690 272.525 808.310 272.695 ;
        RECT 811.305 272.665 811.635 273.055 ;
        RECT 821.395 272.990 821.935 273.860 ;
        RECT 825.305 273.195 827.160 273.365 ;
        RECT 805.690 272.030 805.860 272.525 ;
        RECT 806.280 272.390 806.730 272.525 ;
        RECT 802.915 271.860 805.860 272.030 ;
        RECT 789.250 271.675 791.910 271.845 ;
        RECT 808.140 271.835 808.310 272.525 ;
        RECT 810.630 272.495 811.635 272.665 ;
        RECT 810.630 271.835 810.800 272.495 ;
        RECT 808.140 271.665 810.800 271.835 ;
        RECT 821.765 272.000 821.935 272.990 ;
        RECT 826.990 272.665 827.160 273.195 ;
        RECT 824.540 272.495 827.160 272.665 ;
        RECT 830.155 272.635 830.485 273.025 ;
        RECT 824.540 272.000 824.710 272.495 ;
        RECT 825.140 272.320 825.610 272.495 ;
        RECT 821.765 271.830 824.710 272.000 ;
        RECT 826.990 271.805 827.160 272.495 ;
        RECT 829.480 272.465 830.485 272.635 ;
        RECT 829.480 271.805 829.650 272.465 ;
        RECT 826.990 271.635 829.650 271.805 ;
        RECT 772.440 269.950 774.010 270.680 ;
        RECT 781.480 269.950 782.250 270.270 ;
        RECT 772.440 269.520 782.250 269.950 ;
        RECT 772.440 268.880 774.010 269.520 ;
        RECT 781.480 269.480 782.250 269.520 ;
        RECT 783.665 265.470 784.205 266.340 ;
        RECT 787.575 265.675 789.430 265.845 ;
        RECT 784.035 264.480 784.205 265.470 ;
        RECT 789.260 265.145 789.430 265.675 ;
        RECT 802.195 265.530 802.735 266.400 ;
        RECT 806.105 265.735 807.960 265.905 ;
        RECT 786.810 264.975 789.430 265.145 ;
        RECT 792.425 265.115 792.755 265.505 ;
        RECT 786.810 264.480 786.980 264.975 ;
        RECT 787.400 264.800 787.890 264.975 ;
        RECT 784.035 264.310 786.980 264.480 ;
        RECT 789.260 264.285 789.430 264.975 ;
        RECT 791.750 264.945 792.755 265.115 ;
        RECT 791.750 264.285 791.920 264.945 ;
        RECT 802.565 264.540 802.735 265.530 ;
        RECT 807.790 265.205 807.960 265.735 ;
        RECT 805.340 265.035 807.960 265.205 ;
        RECT 810.955 265.175 811.285 265.565 ;
        RECT 805.340 264.540 805.510 265.035 ;
        RECT 805.920 264.880 806.400 265.035 ;
        RECT 802.565 264.370 805.510 264.540 ;
        RECT 789.260 264.115 791.920 264.285 ;
        RECT 807.790 264.345 807.960 265.035 ;
        RECT 810.280 265.005 811.285 265.175 ;
        RECT 810.280 264.345 810.450 265.005 ;
        RECT 807.790 264.175 810.450 264.345 ;
      LAYER mcon ;
        RECT 665.915 351.975 666.085 352.145 ;
        RECT 684.115 351.905 684.285 352.075 ;
        RECT 701.815 351.925 701.985 352.095 ;
        RECT 719.795 351.905 719.965 352.075 ;
        RECT 737.910 351.895 738.080 352.065 ;
        RECT 755.720 351.865 755.890 352.035 ;
        RECT 773.745 351.745 773.915 351.915 ;
        RECT 791.910 351.825 792.080 351.995 ;
        RECT 810.240 351.830 810.410 352.000 ;
        RECT 802.525 343.675 802.695 343.845 ;
        RECT 821.855 343.605 822.025 343.775 ;
        RECT 802.895 305.100 803.065 305.270 ;
        RECT 820.735 305.100 820.905 305.270 ;
        RECT 685.900 295.855 686.070 296.025 ;
        RECT 703.390 295.835 703.560 296.005 ;
        RECT 721.000 295.865 721.170 296.035 ;
        RECT 738.695 295.810 738.865 295.980 ;
        RECT 756.465 295.865 756.635 296.035 ;
        RECT 787.535 272.440 787.705 272.610 ;
        RECT 806.420 272.445 806.590 272.615 ;
        RECT 825.290 272.390 825.460 272.560 ;
        RECT 772.600 268.975 773.850 270.585 ;
        RECT 781.600 269.610 782.130 270.140 ;
        RECT 787.560 264.880 787.730 265.050 ;
        RECT 806.075 264.935 806.245 265.105 ;
      LAYER met1 ;
        RECT 665.690 351.950 666.350 352.230 ;
        RECT 684.000 352.090 684.400 352.110 ;
        RECT 665.760 351.940 666.240 351.950 ;
        RECT 683.980 351.830 684.440 352.090 ;
        RECT 701.620 351.850 702.190 352.150 ;
        RECT 719.580 351.820 720.190 352.140 ;
        RECT 737.780 352.130 738.210 352.150 ;
        RECT 737.720 351.770 738.250 352.130 ;
        RECT 755.620 351.730 756.030 352.150 ;
        RECT 773.560 351.640 774.120 352.020 ;
        RECT 791.690 351.750 792.310 352.050 ;
        RECT 810.050 351.780 810.610 352.060 ;
        RECT 810.090 351.770 810.560 351.780 ;
        RECT 802.350 343.570 802.870 343.950 ;
        RECT 821.690 343.510 822.190 343.870 ;
        RECT 767.200 305.160 769.770 305.670 ;
        RECT 802.760 305.230 803.200 305.350 ;
        RECT 812.730 305.230 813.360 305.320 ;
        RECT 820.600 305.230 821.040 305.350 ;
        RECT 767.200 304.620 775.880 305.160 ;
        RECT 802.760 305.060 821.040 305.230 ;
        RECT 802.760 305.020 803.200 305.060 ;
        RECT 812.730 304.910 813.360 305.060 ;
        RECT 820.600 305.020 821.040 305.060 ;
        RECT 767.200 304.210 776.360 304.620 ;
        RECT 767.200 303.760 769.770 304.210 ;
        RECT 775.270 302.520 776.360 304.210 ;
        RECT 720.970 296.130 721.200 296.140 ;
        RECT 685.870 296.090 686.100 296.130 ;
        RECT 703.360 296.090 703.590 296.120 ;
        RECT 685.810 295.750 686.220 296.090 ;
        RECT 703.290 295.720 703.670 296.090 ;
        RECT 720.900 295.780 721.260 296.130 ;
        RECT 738.660 296.050 738.900 296.080 ;
        RECT 720.970 295.760 721.200 295.780 ;
        RECT 738.610 295.710 738.970 296.050 ;
        RECT 756.370 295.760 756.740 296.170 ;
        RECT 756.420 295.730 756.680 295.760 ;
        RECT 763.730 293.110 764.830 293.740 ;
        RECT 767.190 293.110 769.200 293.740 ;
        RECT 763.730 292.590 769.200 293.110 ;
        RECT 763.730 292.350 764.830 292.590 ;
        RECT 767.190 292.270 769.200 292.590 ;
        RECT 756.110 286.930 757.150 287.950 ;
        RECT 756.440 282.080 756.780 286.930 ;
        RECT 756.440 281.990 773.300 282.080 ;
        RECT 756.440 281.650 773.580 281.990 ;
        RECT 772.920 270.740 773.580 281.650 ;
        RECT 787.320 272.330 787.920 272.720 ;
        RECT 806.220 272.360 806.790 272.700 ;
        RECT 825.080 272.290 825.670 272.660 ;
        RECT 772.410 268.820 774.040 270.740 ;
        RECT 781.450 270.270 782.280 270.330 ;
        RECT 781.430 269.480 782.300 270.270 ;
        RECT 781.450 269.420 782.280 269.480 ;
        RECT 787.340 264.770 787.950 265.160 ;
        RECT 805.860 264.850 806.460 265.190 ;
      LAYER via ;
        RECT 665.890 351.960 666.150 352.220 ;
        RECT 684.080 351.830 684.340 352.090 ;
        RECT 701.775 351.870 702.035 352.130 ;
        RECT 719.755 351.850 720.015 352.110 ;
        RECT 737.855 351.820 738.115 352.080 ;
        RECT 755.695 351.810 755.955 352.070 ;
        RECT 773.710 351.700 773.970 351.960 ;
        RECT 791.870 351.770 792.130 352.030 ;
        RECT 810.200 351.790 810.460 352.050 ;
        RECT 802.480 343.630 802.740 343.890 ;
        RECT 821.810 343.560 822.070 343.820 ;
        RECT 767.395 303.785 769.575 305.645 ;
        RECT 812.915 304.985 813.175 305.245 ;
        RECT 775.365 302.640 776.265 304.500 ;
        RECT 685.885 295.790 686.145 296.050 ;
        RECT 703.350 295.775 703.610 296.035 ;
        RECT 720.950 295.825 721.210 296.085 ;
        RECT 738.660 295.750 738.920 296.010 ;
        RECT 756.425 295.835 756.685 296.095 ;
        RECT 763.830 292.435 764.730 293.655 ;
        RECT 767.265 292.395 769.125 293.615 ;
        RECT 756.180 286.990 757.080 287.890 ;
        RECT 787.490 272.395 787.750 272.655 ;
        RECT 806.375 272.400 806.635 272.660 ;
        RECT 825.245 272.345 825.505 272.605 ;
        RECT 781.575 269.585 782.155 270.165 ;
        RECT 787.515 264.835 787.775 265.095 ;
        RECT 806.030 264.890 806.290 265.150 ;
      LAYER met2 ;
        RECT 755.480 355.540 756.030 356.260 ;
        RECT 665.740 351.900 666.300 352.280 ;
        RECT 755.700 352.200 755.850 355.540 ;
        RECT 665.890 350.320 666.090 351.900 ;
        RECT 684.030 351.780 684.390 352.140 ;
        RECT 701.670 351.800 702.140 352.200 ;
        RECT 684.090 350.320 684.290 351.780 ;
        RECT 665.870 350.270 684.350 350.320 ;
        RECT 701.780 350.270 701.930 351.800 ;
        RECT 719.630 351.770 720.140 352.190 ;
        RECT 719.810 350.270 719.960 351.770 ;
        RECT 737.770 351.720 738.200 352.180 ;
        RECT 737.860 350.270 738.010 351.720 ;
        RECT 755.670 351.680 755.980 352.200 ;
        RECT 755.720 350.270 755.880 351.680 ;
        RECT 773.610 351.590 774.070 352.070 ;
        RECT 791.740 351.700 792.260 352.100 ;
        RECT 810.100 351.730 810.560 352.110 ;
        RECT 767.970 350.270 768.620 350.280 ;
        RECT 773.740 350.270 773.910 351.590 ;
        RECT 791.890 350.270 792.040 351.700 ;
        RECT 810.240 350.270 810.390 351.730 ;
        RECT 665.870 350.120 810.400 350.270 ;
        RECT 665.870 350.090 684.350 350.120 ;
        RECT 701.780 349.870 701.930 350.120 ;
        RECT 719.810 349.880 719.960 350.120 ;
        RECT 767.970 305.720 768.620 350.120 ;
        RECT 773.740 350.060 773.910 350.120 ;
        RECT 791.890 350.110 792.040 350.120 ;
        RECT 802.590 348.410 802.760 350.120 ;
        RECT 802.590 348.330 822.030 348.410 ;
        RECT 802.590 348.140 822.070 348.330 ;
        RECT 802.590 343.970 802.760 348.140 ;
        RECT 802.410 343.550 802.810 343.970 ;
        RECT 821.860 343.890 822.070 348.140 ;
        RECT 821.750 343.490 822.130 343.890 ;
        RECT 767.250 303.710 769.720 305.720 ;
        RECT 685.860 295.700 686.170 296.140 ;
        RECT 685.910 293.170 686.110 295.700 ;
        RECT 703.340 295.670 703.620 296.140 ;
        RECT 720.950 295.730 721.210 296.180 ;
        RECT 703.410 293.920 703.550 295.670 ;
        RECT 703.410 293.170 703.580 293.920 ;
        RECT 720.960 293.740 721.140 295.730 ;
        RECT 738.660 295.660 738.920 296.100 ;
        RECT 756.420 295.710 756.690 296.220 ;
        RECT 738.740 294.300 738.880 295.660 ;
        RECT 738.740 294.180 738.890 294.300 ;
        RECT 720.970 293.170 721.140 293.740 ;
        RECT 738.750 293.170 738.890 294.180 ;
        RECT 756.470 294.130 756.620 295.710 ;
        RECT 756.470 293.940 756.630 294.130 ;
        RECT 756.440 293.230 756.630 293.940 ;
        RECT 767.970 293.790 768.620 303.710 ;
        RECT 775.010 302.310 776.510 305.250 ;
        RECT 812.780 304.860 813.310 305.370 ;
        RECT 763.780 293.230 764.780 293.790 ;
        RECT 756.430 293.170 764.780 293.230 ;
        RECT 685.910 292.940 764.780 293.170 ;
        RECT 703.410 292.930 703.580 292.940 ;
        RECT 720.970 292.920 721.140 292.940 ;
        RECT 738.750 292.920 738.890 292.940 ;
        RECT 756.430 292.710 764.780 292.940 ;
        RECT 756.440 288.000 756.630 292.710 ;
        RECT 763.780 292.300 764.780 292.710 ;
        RECT 767.240 292.220 769.150 293.790 ;
        RECT 767.970 291.990 768.620 292.220 ;
        RECT 756.160 286.880 757.100 288.000 ;
        RECT 787.380 272.310 787.860 272.740 ;
        RECT 806.280 272.340 806.730 272.720 ;
        RECT 781.480 269.990 782.250 270.320 ;
        RECT 787.540 269.990 787.710 272.310 ;
        RECT 806.450 269.990 806.620 272.340 ;
        RECT 825.140 272.270 825.610 272.680 ;
        RECT 825.270 269.990 825.440 272.270 ;
        RECT 781.480 269.690 825.480 269.990 ;
        RECT 781.480 269.430 782.250 269.690 ;
        RECT 787.490 269.670 825.480 269.690 ;
        RECT 787.540 269.660 787.710 269.670 ;
        RECT 787.400 264.750 787.890 265.180 ;
        RECT 805.920 264.830 806.400 265.210 ;
        RECT 787.450 262.060 787.630 264.750 ;
        RECT 805.970 262.820 806.150 264.830 ;
        RECT 805.970 262.660 806.170 262.820 ;
        RECT 805.980 262.090 806.170 262.660 ;
        RECT 823.690 262.090 823.990 269.670 ;
        RECT 805.980 262.060 824.010 262.090 ;
        RECT 787.450 261.790 824.010 262.060 ;
        RECT 805.980 261.780 824.010 261.790 ;
        RECT 823.690 261.740 823.990 261.780 ;
      LAYER via2 ;
        RECT 755.615 355.760 755.895 356.040 ;
        RECT 775.020 302.440 776.500 305.120 ;
        RECT 812.905 304.975 813.185 305.255 ;
      LAYER met3 ;
        RECT 755.240 355.500 756.280 356.500 ;
        RECT 774.960 303.000 776.560 305.225 ;
        RECT 812.730 304.885 813.360 305.345 ;
        RECT 813.000 303.000 813.350 304.885 ;
        RECT 774.960 302.335 813.450 303.000 ;
        RECT 775.610 302.210 813.450 302.335 ;
      LAYER via3 ;
        RECT 755.400 355.640 756.120 356.360 ;
      LAYER met4 ;
        RECT 754.630 475.830 757.050 490.240 ;
        RECT 754.670 376.270 756.870 475.830 ;
        RECT 754.630 358.110 756.870 376.270 ;
        RECT 754.630 357.400 756.990 358.110 ;
        RECT 754.670 355.970 756.990 357.400 ;
        RECT 754.670 355.850 756.870 355.970 ;
        RECT 755.285 355.495 756.235 355.850 ;
    END
  END re
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.220000 ;
    PORT
      LAYER li1 ;
        RECT 840.420 356.750 841.490 358.080 ;
        RECT 839.525 352.660 840.235 352.665 ;
        RECT 840.670 352.660 841.120 356.750 ;
        RECT 839.525 352.280 841.200 352.660 ;
        RECT 840.030 352.240 841.200 352.280 ;
        RECT 808.320 344.730 808.650 344.830 ;
        RECT 808.300 344.370 808.650 344.730 ;
        RECT 808.320 343.855 808.650 344.370 ;
        RECT 827.680 343.765 828.010 344.740 ;
        RECT 840.640 344.190 841.050 352.240 ;
        RECT 840.330 343.530 841.180 344.190 ;
        RECT 781.520 272.585 781.850 273.560 ;
        RECT 800.410 272.575 800.740 273.550 ;
        RECT 819.260 272.545 819.590 273.520 ;
        RECT 781.530 265.025 781.860 266.000 ;
        RECT 800.060 265.085 800.390 266.060 ;
      LAYER mcon ;
        RECT 840.510 356.790 841.400 358.040 ;
        RECT 808.375 344.465 808.545 344.635 ;
        RECT 827.750 343.880 827.920 344.050 ;
        RECT 840.490 343.595 841.020 344.125 ;
        RECT 781.590 273.035 781.760 273.205 ;
        RECT 800.490 273.235 800.660 273.405 ;
        RECT 800.490 272.875 800.660 273.045 ;
        RECT 819.330 273.185 819.500 273.355 ;
        RECT 819.330 272.825 819.500 272.995 ;
        RECT 781.620 265.635 781.790 265.805 ;
        RECT 781.620 265.275 781.790 265.445 ;
        RECT 800.150 265.725 800.320 265.895 ;
        RECT 800.150 265.365 800.320 265.535 ;
      LAYER met1 ;
        RECT 840.390 358.080 841.520 358.140 ;
        RECT 840.370 356.750 841.540 358.080 ;
        RECT 840.390 356.690 841.520 356.750 ;
        RECT 808.270 344.730 808.650 344.790 ;
        RECT 808.250 344.370 808.670 344.730 ;
        RECT 808.270 344.310 808.650 344.370 ;
        RECT 827.660 344.020 828.010 344.190 ;
        RECT 840.270 344.040 841.240 344.220 ;
        RECT 833.600 344.020 841.240 344.040 ;
        RECT 827.660 343.740 841.240 344.020 ;
        RECT 827.790 343.700 841.240 343.740 ;
        RECT 827.790 343.680 835.030 343.700 ;
        RECT 808.160 341.780 808.830 341.840 ;
        RECT 830.520 341.780 831.010 343.680 ;
        RECT 840.270 343.500 841.240 343.700 ;
        RECT 808.160 341.230 831.010 341.780 ;
        RECT 808.160 341.110 808.830 341.230 ;
        RECT 840.620 333.860 841.060 343.500 ;
        RECT 838.460 331.210 843.260 333.860 ;
        RECT 800.410 273.430 800.740 273.490 ;
        RECT 781.490 272.830 781.860 273.410 ;
        RECT 800.390 272.850 800.760 273.430 ;
        RECT 819.250 273.380 819.580 273.440 ;
        RECT 800.410 272.790 800.740 272.850 ;
        RECT 819.230 272.800 819.600 273.380 ;
        RECT 819.250 272.740 819.580 272.800 ;
        RECT 800.070 265.920 800.400 265.980 ;
        RECT 781.540 265.830 781.870 265.890 ;
        RECT 781.520 265.250 781.890 265.830 ;
        RECT 800.050 265.340 800.420 265.920 ;
        RECT 800.070 265.280 800.400 265.340 ;
        RECT 781.540 265.190 781.870 265.250 ;
      LAYER via ;
        RECT 840.505 356.805 841.405 358.025 ;
        RECT 808.330 344.420 808.590 344.680 ;
        RECT 808.365 341.505 808.625 341.765 ;
        RECT 808.365 341.185 808.625 341.445 ;
        RECT 838.650 331.285 843.070 333.785 ;
        RECT 781.545 273.150 781.805 273.410 ;
        RECT 781.545 272.830 781.805 273.090 ;
        RECT 800.445 273.170 800.705 273.430 ;
        RECT 800.445 272.850 800.705 273.110 ;
        RECT 819.285 273.120 819.545 273.380 ;
        RECT 819.285 272.800 819.545 273.060 ;
        RECT 781.575 265.570 781.835 265.830 ;
        RECT 781.575 265.250 781.835 265.510 ;
        RECT 800.105 265.660 800.365 265.920 ;
        RECT 800.105 265.340 800.365 265.600 ;
      LAYER met2 ;
        RECT 840.420 356.700 841.490 358.130 ;
        RECT 808.300 344.650 808.620 344.780 ;
        RECT 808.300 344.320 808.690 344.650 ;
        RECT 808.470 341.890 808.690 344.320 ;
        RECT 808.210 341.060 808.780 341.890 ;
        RECT 838.510 332.870 843.210 333.910 ;
        RECT 773.370 332.800 843.210 332.870 ;
        RECT 773.300 332.120 843.210 332.800 ;
        RECT 773.300 283.870 774.140 332.120 ;
        RECT 838.510 331.160 843.210 332.120 ;
        RECT 773.300 283.670 780.220 283.870 ;
        RECT 773.300 283.570 780.240 283.670 ;
        RECT 779.800 273.180 780.240 283.570 ;
        RECT 779.780 273.160 780.240 273.180 ;
        RECT 781.540 273.160 781.810 273.460 ;
        RECT 779.780 273.120 781.810 273.160 ;
        RECT 800.440 273.120 800.710 273.480 ;
        RECT 819.280 273.120 819.550 273.430 ;
        RECT 779.780 272.960 819.550 273.120 ;
        RECT 779.780 272.880 780.240 272.960 ;
        RECT 781.540 272.920 819.550 272.960 ;
        RECT 779.780 265.620 780.090 272.880 ;
        RECT 781.540 272.780 781.810 272.920 ;
        RECT 800.440 272.800 800.710 272.920 ;
        RECT 819.280 272.750 819.550 272.920 ;
        RECT 781.570 265.640 781.840 265.880 ;
        RECT 800.100 265.640 800.370 265.970 ;
        RECT 781.550 265.620 800.430 265.640 ;
        RECT 779.780 265.440 800.430 265.620 ;
        RECT 779.780 265.420 781.840 265.440 ;
        RECT 781.570 265.200 781.840 265.420 ;
        RECT 800.100 265.290 800.370 265.440 ;
      LAYER via2 ;
        RECT 840.615 356.875 841.295 357.955 ;
      LAYER met3 ;
        RECT 840.210 356.670 841.730 358.310 ;
      LAYER via3 ;
        RECT 840.410 356.730 841.530 358.250 ;
      LAYER met4 ;
        RECT 839.970 475.630 843.590 489.430 ;
        RECT 840.020 462.560 843.460 475.630 ;
        RECT 839.990 461.880 843.460 462.560 ;
        RECT 839.990 376.780 843.390 461.880 ;
        RECT 839.870 357.840 843.500 376.780 ;
        RECT 840.010 356.530 841.840 357.840 ;
    END
  END clk
  PIN y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.090000 ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 695.730 323.960 695.985 325.955 ;
        RECT 701.350 323.990 702.440 324.200 ;
        RECT 696.790 323.960 702.440 323.990 ;
        RECT 695.710 323.690 702.440 323.960 ;
        RECT 695.730 322.695 695.985 323.690 ;
        RECT 696.790 323.670 702.440 323.690 ;
        RECT 697.390 323.580 702.440 323.670 ;
        RECT 701.350 323.200 702.440 323.580 ;
        RECT 736.275 295.750 736.605 297.045 ;
        RECT 716.645 274.465 717.835 274.840 ;
        RECT 714.845 268.185 715.255 268.855 ;
      LAYER mcon ;
        RECT 701.450 323.255 702.340 324.145 ;
        RECT 736.355 295.840 736.525 296.010 ;
        RECT 716.685 274.630 716.855 274.800 ;
        RECT 714.945 268.460 715.115 268.630 ;
      LAYER met1 ;
        RECT 700.760 322.740 702.800 324.640 ;
        RECT 701.300 308.110 702.160 322.740 ;
        RECT 736.140 308.110 737.230 308.190 ;
        RECT 701.300 307.350 737.230 308.110 ;
        RECT 736.140 306.680 737.230 307.350 ;
        RECT 736.230 295.750 736.660 296.140 ;
        RECT 736.280 295.730 736.600 295.750 ;
        RECT 735.900 294.040 737.160 294.660 ;
        RECT 711.600 289.120 712.820 289.450 ;
        RECT 736.190 289.120 736.820 294.040 ;
        RECT 711.600 288.480 736.970 289.120 ;
        RECT 711.600 288.200 712.820 288.480 ;
        RECT 736.190 288.450 736.820 288.480 ;
        RECT 711.640 274.790 712.550 274.960 ;
        RECT 711.640 274.780 713.640 274.790 ;
        RECT 711.640 274.770 714.060 274.780 ;
        RECT 714.590 274.770 715.150 275.010 ;
        RECT 716.640 274.770 716.900 274.900 ;
        RECT 711.640 274.600 716.900 274.770 ;
        RECT 711.640 274.580 714.060 274.600 ;
        RECT 711.640 274.340 712.550 274.580 ;
        RECT 714.590 274.510 715.150 274.600 ;
        RECT 716.640 274.530 716.900 274.600 ;
        RECT 714.780 268.340 715.290 268.780 ;
        RECT 714.850 268.320 715.210 268.340 ;
      LAYER via ;
        RECT 700.850 322.760 702.710 324.620 ;
        RECT 736.235 306.825 737.135 308.045 ;
        RECT 736.315 295.815 736.575 296.075 ;
        RECT 736.080 294.060 736.980 294.640 ;
        RECT 711.760 288.215 712.660 289.435 ;
        RECT 711.805 274.360 712.385 274.940 ;
        RECT 714.740 274.630 715.000 274.890 ;
        RECT 714.905 268.430 715.165 268.690 ;
      LAYER met2 ;
        RECT 700.810 322.690 702.750 324.690 ;
        RECT 736.190 306.630 737.180 308.240 ;
        RECT 736.330 296.190 736.620 306.630 ;
        RECT 736.280 295.980 736.620 296.190 ;
        RECT 736.280 295.700 736.610 295.980 ;
        RECT 736.350 294.710 736.490 295.700 ;
        RECT 735.950 293.990 737.110 294.710 ;
        RECT 711.650 288.150 712.770 289.500 ;
        RECT 711.980 275.010 712.440 288.150 ;
        RECT 711.690 274.290 712.500 275.010 ;
        RECT 714.640 274.460 715.100 275.060 ;
        RECT 714.890 268.830 715.070 274.460 ;
        RECT 714.830 268.290 715.240 268.830 ;
      LAYER via2 ;
        RECT 700.840 322.750 702.720 324.630 ;
      LAYER met3 ;
        RECT 700.760 322.715 702.800 324.665 ;
      LAYER via3 ;
        RECT 700.820 322.930 702.740 324.450 ;
      LAYER met4 ;
        RECT 646.030 346.940 649.120 490.400 ;
        RECT 646.030 344.400 703.190 346.940 ;
        RECT 700.640 323.190 702.920 344.400 ;
        RECT 700.805 322.735 702.755 323.190 ;
    END
  END y1
  PIN y0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.090000 ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 690.450 330.170 690.725 332.205 ;
        RECT 691.820 330.170 693.070 330.390 ;
        RECT 690.440 329.870 693.070 330.170 ;
        RECT 690.450 328.945 690.725 329.870 ;
        RECT 691.350 329.850 693.070 329.870 ;
        RECT 691.820 329.480 693.070 329.850 ;
        RECT 754.015 295.740 754.345 297.035 ;
        RECT 733.815 274.495 735.005 274.870 ;
        RECT 732.015 268.215 732.425 268.885 ;
      LAYER mcon ;
        RECT 691.820 329.490 693.070 330.380 ;
        RECT 754.100 295.835 754.270 296.005 ;
        RECT 733.855 274.660 734.025 274.830 ;
        RECT 732.115 268.490 732.285 268.660 ;
      LAYER met1 ;
        RECT 694.980 330.520 697.630 331.080 ;
        RECT 753.470 330.520 755.510 331.070 ;
        RECT 692.460 330.420 755.510 330.520 ;
        RECT 691.760 329.650 755.510 330.420 ;
        RECT 691.760 329.450 693.130 329.650 ;
        RECT 694.980 329.000 697.630 329.650 ;
        RECT 753.470 328.810 755.510 329.650 ;
        RECT 753.950 295.770 754.420 296.090 ;
        RECT 753.990 295.760 754.380 295.770 ;
        RECT 753.750 293.900 754.660 294.520 ;
        RECT 753.880 291.870 754.410 293.900 ;
        RECT 729.880 290.670 731.510 291.600 ;
        RECT 753.350 290.630 755.110 291.870 ;
        RECT 730.120 274.820 730.720 275.110 ;
        RECT 730.120 274.800 730.910 274.820 ;
        RECT 731.760 274.800 732.320 275.040 ;
        RECT 733.810 274.800 734.070 274.930 ;
        RECT 730.120 274.630 734.070 274.800 ;
        RECT 730.120 274.600 731.270 274.630 ;
        RECT 730.120 274.590 730.910 274.600 ;
        RECT 730.120 274.400 730.720 274.590 ;
        RECT 731.760 274.540 732.320 274.630 ;
        RECT 733.810 274.560 734.070 274.630 ;
        RECT 731.950 268.370 732.460 268.810 ;
        RECT 732.020 268.350 732.380 268.370 ;
      LAYER via ;
        RECT 695.055 329.110 697.555 330.970 ;
        RECT 753.560 328.850 755.420 331.030 ;
        RECT 754.055 295.800 754.315 296.060 ;
        RECT 753.915 293.920 754.495 294.500 ;
        RECT 730.085 290.685 731.305 291.585 ;
        RECT 753.460 290.640 755.000 291.860 ;
        RECT 730.290 274.785 730.550 275.045 ;
        RECT 730.290 274.465 730.550 274.725 ;
        RECT 731.910 274.660 732.170 274.920 ;
        RECT 732.075 268.460 732.335 268.720 ;
      LAYER met2 ;
        RECT 695.030 328.950 697.580 331.130 ;
        RECT 753.520 328.760 755.460 331.120 ;
        RECT 753.920 319.560 754.470 328.760 ;
        RECT 754.010 296.140 754.390 319.560 ;
        RECT 754.000 295.820 754.390 296.140 ;
        RECT 754.000 295.720 754.370 295.820 ;
        RECT 754.110 294.570 754.280 295.720 ;
        RECT 753.800 293.850 754.610 294.570 ;
        RECT 729.930 291.450 731.460 291.650 ;
        RECT 729.930 291.430 747.350 291.450 ;
        RECT 753.400 291.430 755.060 291.920 ;
        RECT 729.930 290.920 755.060 291.430 ;
        RECT 729.930 290.620 731.460 290.920 ;
        RECT 730.300 275.160 730.870 290.620 ;
        RECT 753.400 290.580 755.060 290.920 ;
        RECT 730.170 274.730 730.870 275.160 ;
        RECT 730.170 274.350 730.670 274.730 ;
        RECT 731.810 274.490 732.270 275.090 ;
        RECT 732.060 268.860 732.240 274.490 ;
        RECT 732.000 268.320 732.410 268.860 ;
      LAYER via2 ;
        RECT 695.165 329.100 697.445 330.980 ;
      LAYER met3 ;
        RECT 694.980 328.975 697.630 331.105 ;
      LAYER via3 ;
        RECT 695.145 329.080 697.465 331.000 ;
      LAYER met4 ;
        RECT 641.390 339.960 644.290 490.570 ;
        RECT 641.390 337.610 697.340 339.960 ;
        RECT 694.980 331.085 697.340 337.610 ;
        RECT 694.980 329.900 697.585 331.085 ;
        RECT 695.025 328.995 697.585 329.900 ;
    END
  END y0
  PIN y2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.095000 ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 694.280 323.375 694.610 323.925 ;
        RECT 686.310 318.250 686.585 320.095 ;
        RECT 686.980 318.250 687.240 318.800 ;
        RECT 687.470 318.250 687.930 318.370 ;
        RECT 686.310 317.870 687.930 318.250 ;
        RECT 686.310 316.835 686.585 317.870 ;
        RECT 686.980 317.730 687.240 317.870 ;
        RECT 687.470 317.830 687.930 317.870 ;
        RECT 689.755 317.785 690.085 319.580 ;
        RECT 718.575 295.800 718.905 297.095 ;
        RECT 699.075 274.365 700.265 274.740 ;
        RECT 697.275 268.085 697.685 268.755 ;
      LAYER mcon ;
        RECT 694.385 323.485 694.555 323.655 ;
        RECT 687.615 318.195 687.785 318.365 ;
        RECT 687.615 317.835 687.785 318.005 ;
        RECT 689.830 318.110 690.000 318.280 ;
        RECT 718.650 295.875 718.820 296.045 ;
        RECT 699.115 274.530 699.285 274.700 ;
        RECT 697.375 268.360 697.545 268.530 ;
      LAYER met1 ;
        RECT 694.280 323.400 694.670 323.770 ;
        RECT 694.320 323.370 694.620 323.400 ;
        RECT 687.440 318.420 687.960 318.430 ;
        RECT 687.400 318.280 688.010 318.420 ;
        RECT 689.760 318.280 690.070 318.410 ;
        RECT 687.400 317.980 690.070 318.280 ;
        RECT 687.400 317.940 689.880 317.980 ;
        RECT 687.400 317.770 688.010 317.940 ;
        RECT 687.040 305.650 688.270 305.790 ;
        RECT 717.410 305.650 719.140 306.270 ;
        RECT 687.040 304.980 719.140 305.650 ;
        RECT 687.040 304.740 688.270 304.980 ;
        RECT 717.410 304.670 719.140 304.980 ;
        RECT 718.520 295.810 718.990 296.110 ;
        RECT 718.230 294.120 719.280 294.660 ;
        RECT 718.540 292.600 718.940 294.120 ;
        RECT 718.210 291.010 719.490 292.600 ;
        RECT 694.130 274.670 694.650 274.980 ;
        RECT 697.020 274.670 697.580 274.910 ;
        RECT 699.070 274.670 699.330 274.800 ;
        RECT 694.130 274.500 699.330 274.670 ;
        RECT 694.130 274.490 696.450 274.500 ;
        RECT 694.130 274.460 694.650 274.490 ;
        RECT 695.940 274.470 696.450 274.490 ;
        RECT 697.020 274.410 697.580 274.500 ;
        RECT 699.070 274.430 699.330 274.500 ;
        RECT 697.210 268.240 697.720 268.680 ;
        RECT 697.280 268.220 697.640 268.240 ;
      LAYER via ;
        RECT 694.345 323.455 694.605 323.715 ;
        RECT 687.575 318.125 687.835 318.385 ;
        RECT 687.575 317.805 687.835 318.065 ;
        RECT 687.205 304.815 688.105 305.715 ;
        RECT 717.505 304.700 719.045 306.240 ;
        RECT 718.625 295.830 718.885 296.090 ;
        RECT 718.305 294.260 718.565 294.520 ;
        RECT 718.625 294.260 718.885 294.520 ;
        RECT 718.945 294.260 719.205 294.520 ;
        RECT 718.400 291.035 719.300 292.575 ;
        RECT 694.260 274.590 694.520 274.850 ;
        RECT 697.170 274.530 697.430 274.790 ;
        RECT 697.335 268.330 697.595 268.590 ;
      LAYER met2 ;
        RECT 694.330 323.350 694.620 323.820 ;
        RECT 687.400 321.100 688.050 321.440 ;
        RECT 694.430 321.100 694.580 323.350 ;
        RECT 687.400 320.930 694.590 321.100 ;
        RECT 687.400 320.680 688.050 320.930 ;
        RECT 687.590 318.660 687.820 320.680 ;
        RECT 687.520 318.470 687.890 318.660 ;
        RECT 687.450 317.720 687.960 318.470 ;
        RECT 687.520 305.840 687.890 317.720 ;
        RECT 687.090 304.690 688.220 305.840 ;
        RECT 717.460 304.620 719.090 306.320 ;
        RECT 718.490 296.160 718.760 304.620 ;
        RECT 718.490 295.940 718.940 296.160 ;
        RECT 718.570 295.760 718.940 295.940 ;
        RECT 718.610 294.710 718.810 295.760 ;
        RECT 718.280 294.070 719.230 294.710 ;
        RECT 718.260 292.280 719.440 292.650 ;
        RECT 694.040 291.820 719.440 292.280 ;
        RECT 694.050 275.030 694.370 291.820 ;
        RECT 718.260 290.960 719.440 291.820 ;
        RECT 694.050 274.800 694.600 275.030 ;
        RECT 694.180 274.410 694.600 274.800 ;
        RECT 697.070 274.360 697.530 274.960 ;
        RECT 697.320 268.730 697.500 274.360 ;
        RECT 697.260 268.190 697.670 268.730 ;
      LAYER via2 ;
        RECT 687.585 320.920 687.865 321.200 ;
      LAYER met3 ;
        RECT 687.300 320.970 688.250 321.740 ;
        RECT 687.350 320.705 688.100 320.970 ;
      LAYER via3 ;
        RECT 687.415 321.275 687.735 321.595 ;
        RECT 687.815 321.275 688.135 321.595 ;
        RECT 687.415 320.875 687.735 321.195 ;
      LAYER met4 ;
        RECT 635.190 335.710 638.510 490.240 ;
        RECT 635.190 334.040 689.210 335.710 ;
        RECT 687.520 322.380 689.160 334.040 ;
        RECT 687.070 322.080 689.160 322.380 ;
        RECT 687.070 321.810 689.150 322.080 ;
        RECT 687.070 320.910 688.460 321.810 ;
        RECT 687.395 320.725 688.055 320.910 ;
    END
  END y2
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.670000 ;
    PORT
      LAYER li1 ;
        RECT 716.625 252.935 717.815 253.310 ;
        RECT 714.825 246.655 715.235 247.325 ;
      LAYER mcon ;
        RECT 716.665 253.100 716.835 253.270 ;
        RECT 714.925 246.930 715.095 247.100 ;
      LAYER met1 ;
        RECT 712.950 253.250 713.790 253.640 ;
        RECT 712.950 253.240 714.040 253.250 ;
        RECT 714.570 253.240 715.130 253.480 ;
        RECT 716.620 253.240 716.880 253.370 ;
        RECT 712.950 253.070 716.880 253.240 ;
        RECT 712.950 253.050 714.040 253.070 ;
        RECT 712.950 252.970 713.790 253.050 ;
        RECT 714.570 252.980 715.130 253.070 ;
        RECT 716.620 253.000 716.880 253.070 ;
        RECT 714.760 246.810 715.270 247.250 ;
        RECT 714.830 246.790 715.190 246.810 ;
      LAYER via ;
        RECT 713.080 253.015 713.660 253.595 ;
        RECT 714.720 253.100 714.980 253.360 ;
        RECT 714.885 246.900 715.145 247.160 ;
      LAYER met2 ;
        RECT 713.000 252.920 713.740 253.690 ;
        RECT 714.620 252.930 715.080 253.530 ;
        RECT 714.870 247.300 715.050 252.930 ;
        RECT 714.810 246.760 715.220 247.300 ;
      LAYER via2 ;
        RECT 713.030 253.165 713.310 253.445 ;
        RECT 713.430 253.165 713.710 253.445 ;
      LAYER met3 ;
        RECT 625.150 318.250 627.960 319.770 ;
        RECT 625.860 300.910 627.430 318.250 ;
        RECT 625.290 299.290 628.150 300.910 ;
        RECT 712.870 252.820 713.860 253.750 ;
      LAYER via3 ;
        RECT 625.395 318.250 627.715 319.770 ;
        RECT 625.360 299.340 628.080 300.860 ;
        RECT 713.005 252.925 713.725 253.645 ;
      LAYER met4 ;
        RECT 625.630 319.775 628.240 490.000 ;
        RECT 625.195 318.920 628.240 319.775 ;
        RECT 625.195 318.245 627.915 318.920 ;
        RECT 625.335 299.285 628.105 300.915 ;
        RECT 625.760 242.100 627.560 299.285 ;
        RECT 712.440 252.270 714.390 254.470 ;
        RECT 713.210 245.270 713.580 252.270 ;
        RECT 625.760 241.960 672.740 242.100 ;
        RECT 713.100 241.960 713.650 245.270 ;
        RECT 625.760 240.940 713.650 241.960 ;
        RECT 625.760 240.870 672.740 240.940 ;
        RECT 713.100 240.870 713.650 240.940 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.670000 ;
    PORT
      LAYER li1 ;
        RECT 733.795 252.965 734.985 253.340 ;
        RECT 731.995 246.685 732.405 247.355 ;
      LAYER mcon ;
        RECT 733.835 253.130 734.005 253.300 ;
        RECT 732.095 246.960 732.265 247.130 ;
      LAYER met1 ;
        RECT 729.970 253.280 730.880 253.720 ;
        RECT 729.970 253.270 730.900 253.280 ;
        RECT 731.740 253.270 732.300 253.510 ;
        RECT 733.790 253.270 734.050 253.400 ;
        RECT 729.970 253.100 734.050 253.270 ;
        RECT 729.970 253.070 731.250 253.100 ;
        RECT 729.970 252.630 730.880 253.070 ;
        RECT 731.740 253.010 732.300 253.100 ;
        RECT 733.790 253.030 734.050 253.100 ;
        RECT 731.930 246.840 732.440 247.280 ;
        RECT 732.000 246.820 732.360 246.840 ;
      LAYER via ;
        RECT 730.135 252.725 730.715 253.625 ;
        RECT 731.890 253.130 732.150 253.390 ;
        RECT 732.055 246.930 732.315 247.190 ;
      LAYER met2 ;
        RECT 730.020 252.580 730.830 253.770 ;
        RECT 731.790 252.960 732.250 253.560 ;
        RECT 732.040 247.330 732.220 252.960 ;
        RECT 731.980 246.790 732.390 247.330 ;
      LAYER via2 ;
        RECT 730.085 252.635 730.765 253.715 ;
      LAYER met3 ;
        RECT 617.070 318.180 620.360 320.140 ;
        RECT 617.570 301.290 619.720 318.180 ;
        RECT 617.100 298.840 620.820 301.290 ;
        RECT 729.830 252.480 730.920 253.880 ;
      LAYER via3 ;
        RECT 617.155 318.200 620.275 320.120 ;
        RECT 617.200 298.905 620.720 301.225 ;
        RECT 730.015 252.620 730.735 253.740 ;
      LAYER met4 ;
        RECT 617.270 320.145 620.260 489.770 ;
        RECT 617.115 318.175 620.315 320.145 ;
        RECT 617.145 298.835 620.775 301.295 ;
        RECT 617.640 238.140 620.090 298.835 ;
        RECT 729.520 252.190 731.090 254.520 ;
        RECT 729.530 241.420 730.980 252.190 ;
        RECT 729.480 238.140 731.080 241.420 ;
        RECT 617.640 238.030 731.080 238.140 ;
        RECT 617.640 236.460 731.070 238.030 ;
        RECT 617.770 236.430 731.070 236.460 ;
        RECT 617.770 236.360 731.020 236.430 ;
    END
  END a1
  OBS
      LAYER pwell ;
        RECT 639.390 322.990 640.730 324.250 ;
        RECT 643.440 323.040 644.780 324.300 ;
        RECT 869.740 323.700 872.870 330.840 ;
        RECT 645.910 308.850 646.820 310.420 ;
        RECT 639.240 304.820 640.580 306.080 ;
        RECT 643.290 304.870 644.630 306.130 ;
        RECT 639.190 285.640 640.530 286.900 ;
        RECT 643.240 285.690 644.580 286.950 ;
        RECT 645.720 271.190 646.630 272.760 ;
        RECT 639.110 267.170 640.450 268.430 ;
        RECT 643.160 267.220 644.500 268.480 ;
        RECT 638.960 249.440 640.300 250.700 ;
        RECT 643.010 249.490 644.350 250.750 ;
        RECT 9.600 190.020 36.600 217.160 ;
        RECT 74.700 190.100 101.700 217.240 ;
        RECT 107.150 190.020 134.150 217.160 ;
        RECT 139.760 190.100 166.760 217.240 ;
        RECT 204.760 190.130 231.760 217.270 ;
        RECT 237.700 190.240 264.700 217.380 ;
        RECT 9.600 160.940 36.600 188.080 ;
        RECT 74.700 161.020 101.700 188.160 ;
        RECT 107.150 160.940 134.150 188.080 ;
        RECT 139.760 161.020 166.760 188.160 ;
        RECT 204.760 161.050 231.760 188.190 ;
        RECT 237.700 161.160 264.700 188.300 ;
        RECT 9.600 131.770 36.600 158.910 ;
        RECT 74.700 131.850 101.700 158.990 ;
        RECT 107.150 131.770 134.150 158.910 ;
        RECT 139.760 131.850 166.760 158.990 ;
        RECT 204.760 131.880 231.760 159.020 ;
        RECT 237.700 131.990 264.700 159.130 ;
        RECT 9.600 102.590 36.600 129.730 ;
        RECT 74.700 102.670 101.700 129.810 ;
        RECT 107.150 102.590 134.150 129.730 ;
        RECT 139.760 102.670 166.760 129.810 ;
        RECT 204.760 102.700 231.760 129.840 ;
        RECT 237.700 102.810 264.700 129.950 ;
        RECT 342.680 102.590 369.680 129.730 ;
        RECT 442.320 102.420 469.320 129.560 ;
        RECT 9.600 73.270 36.600 100.410 ;
        RECT 74.700 73.350 101.700 100.490 ;
        RECT 107.150 73.270 134.150 100.410 ;
        RECT 139.760 73.350 166.760 100.490 ;
        RECT 204.760 73.380 231.760 100.520 ;
        RECT 237.700 73.490 264.700 100.630 ;
        RECT 342.720 73.470 369.720 100.610 ;
        RECT 408.500 73.330 435.500 100.470 ;
        RECT 442.350 73.230 469.350 100.370 ;
        RECT 9.650 43.990 36.650 71.130 ;
        RECT 74.750 44.070 101.750 71.210 ;
        RECT 107.200 43.990 134.200 71.130 ;
        RECT 139.810 44.070 166.810 71.210 ;
        RECT 204.810 44.100 231.810 71.240 ;
        RECT 342.740 44.110 369.740 71.250 ;
        RECT 408.520 43.970 435.520 71.110 ;
        RECT 442.350 43.940 469.350 71.080 ;
        RECT 9.740 14.450 36.740 41.590 ;
        RECT 107.290 14.450 134.290 41.590 ;
        RECT 139.900 14.530 166.900 41.670 ;
        RECT 172.450 14.560 199.450 41.700 ;
        RECT 204.900 14.560 231.900 41.700 ;
        RECT 342.760 14.820 369.760 41.960 ;
        RECT 408.540 14.680 435.540 41.820 ;
        RECT 442.350 14.650 469.350 41.790 ;
      LAYER li1 ;
        RECT 379.300 369.530 379.470 370.180 ;
        RECT 379.160 368.850 379.550 369.530 ;
        RECT 385.880 369.480 386.050 370.180 ;
        RECT 385.750 369.380 386.140 369.480 ;
        RECT 385.630 369.310 386.140 369.380 ;
        RECT 385.630 368.860 386.160 369.310 ;
        RECT 385.060 368.850 386.160 368.860 ;
        RECT 379.160 368.470 386.160 368.850 ;
        RECT 379.160 368.460 385.140 368.470 ;
        RECT 379.220 368.450 385.140 368.460 ;
        RECT 385.760 368.430 386.160 368.470 ;
        RECT 379.160 365.450 379.330 365.610 ;
        RECT 379.110 351.450 379.390 365.450 ;
        RECT 385.740 365.220 385.910 365.610 ;
        RECT 379.060 351.230 379.390 351.450 ;
        RECT 385.680 351.440 385.960 365.220 ;
        RECT 654.065 353.035 654.450 354.615 ;
        RECT 652.900 352.630 653.420 352.730 ;
        RECT 654.065 352.630 654.395 353.035 ;
        RECT 652.900 352.320 654.395 352.630 ;
        RECT 654.575 352.750 655.285 352.795 ;
        RECT 657.675 352.750 658.010 354.585 ;
        RECT 659.315 352.855 659.565 353.855 ;
        RECT 660.820 353.555 661.070 354.025 ;
        RECT 663.230 353.695 663.480 354.605 ;
        RECT 665.300 354.485 666.330 354.655 ;
        RECT 665.300 354.125 665.470 354.485 ;
        RECT 654.575 352.490 658.010 352.750 ;
        RECT 658.190 352.525 659.565 352.855 ;
        RECT 654.575 352.410 655.285 352.490 ;
        RECT 652.900 352.150 653.420 352.320 ;
        RECT 379.060 350.240 379.360 351.230 ;
        RECT 385.680 351.000 386.000 351.440 ;
        RECT 654.065 351.355 654.395 352.320 ;
        RECT 385.700 350.260 386.000 351.000 ;
        RECT 656.220 350.290 656.610 352.490 ;
        RECT 657.675 351.515 658.010 352.490 ;
        RECT 659.355 352.345 659.565 352.525 ;
        RECT 660.065 353.385 661.070 353.555 ;
        RECT 662.605 353.525 663.480 353.695 ;
        RECT 663.660 353.955 665.470 354.125 ;
        RECT 660.065 352.855 660.235 353.385 ;
        RECT 662.605 353.205 662.775 353.525 ;
        RECT 660.415 353.035 662.775 353.205 ;
        RECT 660.065 352.685 662.105 352.855 ;
        RECT 659.355 351.845 659.685 352.345 ;
        RECT 660.065 351.845 660.290 352.685 ;
        RECT 661.775 352.295 662.105 352.685 ;
        RECT 659.960 351.345 660.290 351.845 ;
        RECT 662.310 351.635 662.480 353.035 ;
        RECT 662.955 352.785 663.285 353.285 ;
        RECT 663.660 352.605 663.830 353.955 ;
        RECT 662.660 352.435 663.830 352.605 ;
        RECT 664.010 353.195 664.340 353.775 ;
        RECT 665.650 353.545 665.980 354.305 ;
        RECT 666.160 353.895 666.330 354.485 ;
        RECT 667.640 354.485 669.380 354.655 ;
        RECT 667.640 353.895 667.810 354.485 ;
        RECT 668.000 354.050 668.330 354.305 ;
        RECT 666.160 353.850 667.810 353.895 ;
        RECT 666.160 353.725 667.930 353.850 ;
        RECT 665.650 353.375 667.420 353.545 ;
        RECT 667.600 353.530 667.930 353.725 ;
        RECT 667.250 353.350 667.420 353.375 ;
        RECT 668.110 353.350 668.280 354.050 ;
        RECT 664.010 353.025 667.070 353.195 ;
        RECT 662.660 351.935 662.945 352.435 ;
        RECT 664.010 352.175 664.270 353.025 ;
        RECT 666.740 352.675 667.070 353.025 ;
        RECT 667.250 353.180 668.280 353.350 ;
        RECT 668.460 353.520 668.680 353.850 ;
        RECT 668.860 353.690 669.030 354.305 ;
        RECT 669.210 354.040 669.380 354.485 ;
        RECT 670.070 354.485 671.510 354.655 ;
        RECT 670.070 354.040 670.240 354.485 ;
        RECT 669.210 353.870 670.240 354.040 ;
        RECT 670.420 353.690 670.670 354.305 ;
        RECT 668.860 353.520 670.670 353.690 ;
        RECT 667.250 352.495 667.420 353.180 ;
        RECT 668.460 353.000 668.630 353.520 ;
        RECT 668.860 353.340 669.030 353.520 ;
        RECT 664.800 352.325 667.420 352.495 ;
        RECT 663.150 351.635 663.480 352.175 ;
        RECT 662.310 351.465 663.480 351.635 ;
        RECT 663.940 351.465 664.270 352.175 ;
        RECT 667.250 352.095 667.420 352.325 ;
        RECT 667.605 352.770 668.630 353.000 ;
        RECT 668.810 353.170 669.030 353.340 ;
        RECT 667.605 352.275 667.935 352.770 ;
        RECT 668.810 352.175 668.980 353.170 ;
        RECT 670.910 353.000 671.160 354.305 ;
        RECT 667.250 351.925 668.260 352.095 ;
        RECT 667.930 351.675 668.260 351.925 ;
        RECT 668.710 351.675 668.980 352.175 ;
        RECT 669.165 351.660 669.495 352.955 ;
        RECT 670.635 352.770 671.160 353.000 ;
        RECT 670.890 351.845 671.160 352.770 ;
        RECT 671.340 353.375 671.510 354.485 ;
        RECT 672.470 353.375 672.800 354.305 ;
        RECT 671.340 353.205 672.800 353.375 ;
        RECT 671.340 352.705 671.670 353.205 ;
        RECT 672.020 352.025 672.350 353.000 ;
        RECT 670.890 351.345 671.220 351.845 ;
        RECT 672.530 351.345 672.800 353.205 ;
        RECT 675.725 351.475 676.060 354.545 ;
        RECT 677.365 352.815 677.615 353.815 ;
        RECT 678.870 353.515 679.120 353.985 ;
        RECT 681.280 353.655 681.530 354.565 ;
        RECT 683.350 354.445 684.380 354.615 ;
        RECT 683.350 354.085 683.520 354.445 ;
        RECT 676.240 352.485 677.615 352.815 ;
        RECT 677.405 352.305 677.615 352.485 ;
        RECT 678.115 353.345 679.120 353.515 ;
        RECT 680.655 353.485 681.530 353.655 ;
        RECT 681.710 353.915 683.520 354.085 ;
        RECT 678.115 352.815 678.285 353.345 ;
        RECT 680.655 353.165 680.825 353.485 ;
        RECT 678.465 352.995 680.825 353.165 ;
        RECT 678.115 352.645 680.155 352.815 ;
        RECT 677.405 351.805 677.735 352.305 ;
        RECT 678.115 351.805 678.340 352.645 ;
        RECT 679.825 352.255 680.155 352.645 ;
        RECT 678.010 351.305 678.340 351.805 ;
        RECT 680.360 351.595 680.530 352.995 ;
        RECT 681.005 352.745 681.335 353.245 ;
        RECT 681.710 352.565 681.880 353.915 ;
        RECT 680.710 352.395 681.880 352.565 ;
        RECT 682.060 353.155 682.390 353.735 ;
        RECT 683.700 353.505 684.030 354.265 ;
        RECT 684.210 353.855 684.380 354.445 ;
        RECT 685.690 354.445 687.430 354.615 ;
        RECT 685.690 353.855 685.860 354.445 ;
        RECT 686.050 354.010 686.380 354.265 ;
        RECT 684.210 353.810 685.860 353.855 ;
        RECT 684.210 353.685 685.980 353.810 ;
        RECT 683.700 353.335 685.470 353.505 ;
        RECT 685.650 353.490 685.980 353.685 ;
        RECT 685.300 353.310 685.470 353.335 ;
        RECT 686.160 353.310 686.330 354.010 ;
        RECT 682.060 352.985 685.120 353.155 ;
        RECT 680.710 351.895 680.995 352.395 ;
        RECT 682.060 352.135 682.320 352.985 ;
        RECT 684.790 352.635 685.120 352.985 ;
        RECT 685.300 353.140 686.330 353.310 ;
        RECT 686.510 353.480 686.730 353.810 ;
        RECT 686.910 353.650 687.080 354.265 ;
        RECT 687.260 354.000 687.430 354.445 ;
        RECT 688.120 354.445 689.560 354.615 ;
        RECT 688.120 354.000 688.290 354.445 ;
        RECT 687.260 353.830 688.290 354.000 ;
        RECT 688.470 353.650 688.720 354.265 ;
        RECT 686.910 353.480 688.720 353.650 ;
        RECT 685.300 352.455 685.470 353.140 ;
        RECT 686.510 352.960 686.680 353.480 ;
        RECT 686.910 353.300 687.080 353.480 ;
        RECT 682.850 352.285 685.470 352.455 ;
        RECT 681.200 351.595 681.530 352.135 ;
        RECT 680.360 351.425 681.530 351.595 ;
        RECT 681.990 351.425 682.320 352.135 ;
        RECT 685.300 352.055 685.470 352.285 ;
        RECT 685.655 352.730 686.680 352.960 ;
        RECT 686.860 353.130 687.080 353.300 ;
        RECT 685.655 352.235 685.985 352.730 ;
        RECT 686.860 352.135 687.030 353.130 ;
        RECT 688.960 352.960 689.210 354.265 ;
        RECT 685.300 351.885 686.310 352.055 ;
        RECT 685.980 351.635 686.310 351.885 ;
        RECT 686.760 351.635 687.030 352.135 ;
        RECT 687.215 351.620 687.545 352.915 ;
        RECT 688.685 352.730 689.210 352.960 ;
        RECT 688.940 351.805 689.210 352.730 ;
        RECT 689.390 353.335 689.560 354.445 ;
        RECT 690.520 353.335 690.850 354.265 ;
        RECT 689.390 353.165 690.850 353.335 ;
        RECT 689.390 352.665 689.720 353.165 ;
        RECT 690.070 351.985 690.400 352.960 ;
        RECT 688.940 351.305 689.270 351.805 ;
        RECT 690.580 351.305 690.850 353.165 ;
        RECT 693.315 351.495 693.650 354.565 ;
        RECT 694.955 352.835 695.205 353.835 ;
        RECT 696.460 353.535 696.710 354.005 ;
        RECT 698.870 353.675 699.120 354.585 ;
        RECT 700.940 354.465 701.970 354.635 ;
        RECT 700.940 354.105 701.110 354.465 ;
        RECT 693.830 352.505 695.205 352.835 ;
        RECT 694.995 352.325 695.205 352.505 ;
        RECT 695.705 353.365 696.710 353.535 ;
        RECT 698.245 353.505 699.120 353.675 ;
        RECT 699.300 353.935 701.110 354.105 ;
        RECT 695.705 352.835 695.875 353.365 ;
        RECT 698.245 353.185 698.415 353.505 ;
        RECT 696.055 353.015 698.415 353.185 ;
        RECT 695.705 352.665 697.745 352.835 ;
        RECT 694.995 351.825 695.325 352.325 ;
        RECT 695.705 351.825 695.930 352.665 ;
        RECT 697.415 352.275 697.745 352.665 ;
        RECT 695.600 351.325 695.930 351.825 ;
        RECT 697.950 351.615 698.120 353.015 ;
        RECT 698.595 352.765 698.925 353.265 ;
        RECT 699.300 352.585 699.470 353.935 ;
        RECT 698.300 352.415 699.470 352.585 ;
        RECT 699.650 353.175 699.980 353.755 ;
        RECT 701.290 353.525 701.620 354.285 ;
        RECT 701.800 353.875 701.970 354.465 ;
        RECT 703.280 354.465 705.020 354.635 ;
        RECT 703.280 353.875 703.450 354.465 ;
        RECT 703.640 354.030 703.970 354.285 ;
        RECT 701.800 353.830 703.450 353.875 ;
        RECT 701.800 353.705 703.570 353.830 ;
        RECT 701.290 353.355 703.060 353.525 ;
        RECT 703.240 353.510 703.570 353.705 ;
        RECT 702.890 353.330 703.060 353.355 ;
        RECT 703.750 353.330 703.920 354.030 ;
        RECT 699.650 353.005 702.710 353.175 ;
        RECT 698.300 351.915 698.585 352.415 ;
        RECT 699.650 352.155 699.910 353.005 ;
        RECT 702.380 352.655 702.710 353.005 ;
        RECT 702.890 353.160 703.920 353.330 ;
        RECT 704.100 353.500 704.320 353.830 ;
        RECT 704.500 353.670 704.670 354.285 ;
        RECT 704.850 354.020 705.020 354.465 ;
        RECT 705.710 354.465 707.150 354.635 ;
        RECT 705.710 354.020 705.880 354.465 ;
        RECT 704.850 353.850 705.880 354.020 ;
        RECT 706.060 353.670 706.310 354.285 ;
        RECT 704.500 353.500 706.310 353.670 ;
        RECT 702.890 352.475 703.060 353.160 ;
        RECT 704.100 352.980 704.270 353.500 ;
        RECT 704.500 353.320 704.670 353.500 ;
        RECT 700.440 352.305 703.060 352.475 ;
        RECT 698.790 351.615 699.120 352.155 ;
        RECT 697.950 351.445 699.120 351.615 ;
        RECT 699.580 351.445 699.910 352.155 ;
        RECT 702.890 352.075 703.060 352.305 ;
        RECT 703.245 352.750 704.270 352.980 ;
        RECT 704.450 353.150 704.670 353.320 ;
        RECT 703.245 352.255 703.575 352.750 ;
        RECT 704.450 352.155 704.620 353.150 ;
        RECT 706.550 352.980 706.800 354.285 ;
        RECT 702.890 351.905 703.900 352.075 ;
        RECT 703.570 351.655 703.900 351.905 ;
        RECT 704.350 351.655 704.620 352.155 ;
        RECT 704.805 351.640 705.135 352.935 ;
        RECT 706.275 352.750 706.800 352.980 ;
        RECT 706.530 351.825 706.800 352.750 ;
        RECT 706.980 353.355 707.150 354.465 ;
        RECT 708.110 353.355 708.440 354.285 ;
        RECT 706.980 353.185 708.440 353.355 ;
        RECT 706.980 352.685 707.310 353.185 ;
        RECT 707.660 352.005 707.990 352.980 ;
        RECT 706.530 351.325 706.860 351.825 ;
        RECT 708.170 351.325 708.440 353.185 ;
        RECT 711.165 351.495 711.500 354.565 ;
        RECT 712.805 352.835 713.055 353.835 ;
        RECT 714.310 353.535 714.560 354.005 ;
        RECT 716.720 353.675 716.970 354.585 ;
        RECT 718.790 354.465 719.820 354.635 ;
        RECT 718.790 354.105 718.960 354.465 ;
        RECT 711.680 352.505 713.055 352.835 ;
        RECT 712.845 352.325 713.055 352.505 ;
        RECT 713.555 353.365 714.560 353.535 ;
        RECT 716.095 353.505 716.970 353.675 ;
        RECT 717.150 353.935 718.960 354.105 ;
        RECT 713.555 352.835 713.725 353.365 ;
        RECT 716.095 353.185 716.265 353.505 ;
        RECT 713.905 353.015 716.265 353.185 ;
        RECT 713.555 352.665 715.595 352.835 ;
        RECT 712.845 351.825 713.175 352.325 ;
        RECT 713.555 351.825 713.780 352.665 ;
        RECT 715.265 352.275 715.595 352.665 ;
        RECT 713.450 351.325 713.780 351.825 ;
        RECT 715.800 351.615 715.970 353.015 ;
        RECT 716.445 352.765 716.775 353.265 ;
        RECT 717.150 352.585 717.320 353.935 ;
        RECT 716.150 352.415 717.320 352.585 ;
        RECT 717.500 353.175 717.830 353.755 ;
        RECT 719.140 353.525 719.470 354.285 ;
        RECT 719.650 353.875 719.820 354.465 ;
        RECT 721.130 354.465 722.870 354.635 ;
        RECT 721.130 353.875 721.300 354.465 ;
        RECT 721.490 354.030 721.820 354.285 ;
        RECT 719.650 353.830 721.300 353.875 ;
        RECT 719.650 353.705 721.420 353.830 ;
        RECT 719.140 353.355 720.910 353.525 ;
        RECT 721.090 353.510 721.420 353.705 ;
        RECT 720.740 353.330 720.910 353.355 ;
        RECT 721.600 353.330 721.770 354.030 ;
        RECT 717.500 353.005 720.560 353.175 ;
        RECT 716.150 351.915 716.435 352.415 ;
        RECT 717.500 352.155 717.760 353.005 ;
        RECT 720.230 352.655 720.560 353.005 ;
        RECT 720.740 353.160 721.770 353.330 ;
        RECT 721.950 353.500 722.170 353.830 ;
        RECT 722.350 353.670 722.520 354.285 ;
        RECT 722.700 354.020 722.870 354.465 ;
        RECT 723.560 354.465 725.000 354.635 ;
        RECT 723.560 354.020 723.730 354.465 ;
        RECT 722.700 353.850 723.730 354.020 ;
        RECT 723.910 353.670 724.160 354.285 ;
        RECT 722.350 353.500 724.160 353.670 ;
        RECT 720.740 352.475 720.910 353.160 ;
        RECT 721.950 352.980 722.120 353.500 ;
        RECT 722.350 353.320 722.520 353.500 ;
        RECT 718.290 352.305 720.910 352.475 ;
        RECT 716.640 351.615 716.970 352.155 ;
        RECT 715.800 351.445 716.970 351.615 ;
        RECT 717.430 351.445 717.760 352.155 ;
        RECT 720.740 352.075 720.910 352.305 ;
        RECT 721.095 352.750 722.120 352.980 ;
        RECT 722.300 353.150 722.520 353.320 ;
        RECT 721.095 352.255 721.425 352.750 ;
        RECT 722.300 352.155 722.470 353.150 ;
        RECT 724.400 352.980 724.650 354.285 ;
        RECT 720.740 351.905 721.750 352.075 ;
        RECT 721.420 351.655 721.750 351.905 ;
        RECT 722.200 351.655 722.470 352.155 ;
        RECT 722.655 351.640 722.985 352.935 ;
        RECT 724.125 352.750 724.650 352.980 ;
        RECT 724.380 351.825 724.650 352.750 ;
        RECT 724.830 353.355 725.000 354.465 ;
        RECT 725.960 353.355 726.290 354.285 ;
        RECT 724.830 353.185 726.290 353.355 ;
        RECT 724.830 352.685 725.160 353.185 ;
        RECT 725.510 352.005 725.840 352.980 ;
        RECT 724.380 351.325 724.710 351.825 ;
        RECT 726.020 351.325 726.290 353.185 ;
        RECT 729.425 351.495 729.760 354.565 ;
        RECT 731.065 352.835 731.315 353.835 ;
        RECT 732.570 353.535 732.820 354.005 ;
        RECT 734.980 353.675 735.230 354.585 ;
        RECT 737.050 354.465 738.080 354.635 ;
        RECT 737.050 354.105 737.220 354.465 ;
        RECT 729.940 352.505 731.315 352.835 ;
        RECT 731.105 352.325 731.315 352.505 ;
        RECT 731.815 353.365 732.820 353.535 ;
        RECT 734.355 353.505 735.230 353.675 ;
        RECT 735.410 353.935 737.220 354.105 ;
        RECT 731.815 352.835 731.985 353.365 ;
        RECT 734.355 353.185 734.525 353.505 ;
        RECT 732.165 353.015 734.525 353.185 ;
        RECT 731.815 352.665 733.855 352.835 ;
        RECT 731.105 351.825 731.435 352.325 ;
        RECT 731.815 351.825 732.040 352.665 ;
        RECT 733.525 352.275 733.855 352.665 ;
        RECT 731.710 351.325 732.040 351.825 ;
        RECT 734.060 351.615 734.230 353.015 ;
        RECT 734.705 352.765 735.035 353.265 ;
        RECT 735.410 352.585 735.580 353.935 ;
        RECT 734.410 352.415 735.580 352.585 ;
        RECT 735.760 353.175 736.090 353.755 ;
        RECT 737.400 353.525 737.730 354.285 ;
        RECT 737.910 353.875 738.080 354.465 ;
        RECT 739.390 354.465 741.130 354.635 ;
        RECT 739.390 353.875 739.560 354.465 ;
        RECT 739.750 354.030 740.080 354.285 ;
        RECT 737.910 353.830 739.560 353.875 ;
        RECT 737.910 353.705 739.680 353.830 ;
        RECT 737.400 353.355 739.170 353.525 ;
        RECT 739.350 353.510 739.680 353.705 ;
        RECT 739.000 353.330 739.170 353.355 ;
        RECT 739.860 353.330 740.030 354.030 ;
        RECT 735.760 353.005 738.820 353.175 ;
        RECT 734.410 351.915 734.695 352.415 ;
        RECT 735.760 352.155 736.020 353.005 ;
        RECT 738.490 352.655 738.820 353.005 ;
        RECT 739.000 353.160 740.030 353.330 ;
        RECT 740.210 353.500 740.430 353.830 ;
        RECT 740.610 353.670 740.780 354.285 ;
        RECT 740.960 354.020 741.130 354.465 ;
        RECT 741.820 354.465 743.260 354.635 ;
        RECT 741.820 354.020 741.990 354.465 ;
        RECT 740.960 353.850 741.990 354.020 ;
        RECT 742.170 353.670 742.420 354.285 ;
        RECT 740.610 353.500 742.420 353.670 ;
        RECT 739.000 352.475 739.170 353.160 ;
        RECT 740.210 352.980 740.380 353.500 ;
        RECT 740.610 353.320 740.780 353.500 ;
        RECT 736.550 352.305 739.170 352.475 ;
        RECT 734.900 351.615 735.230 352.155 ;
        RECT 734.060 351.445 735.230 351.615 ;
        RECT 735.690 351.445 736.020 352.155 ;
        RECT 739.000 352.075 739.170 352.305 ;
        RECT 739.355 352.750 740.380 352.980 ;
        RECT 740.560 353.150 740.780 353.320 ;
        RECT 739.355 352.255 739.685 352.750 ;
        RECT 740.560 352.155 740.730 353.150 ;
        RECT 742.660 352.980 742.910 354.285 ;
        RECT 739.000 351.905 740.010 352.075 ;
        RECT 739.680 351.655 740.010 351.905 ;
        RECT 740.460 351.655 740.730 352.155 ;
        RECT 740.915 351.640 741.245 352.935 ;
        RECT 742.385 352.750 742.910 352.980 ;
        RECT 742.640 351.825 742.910 352.750 ;
        RECT 743.090 353.355 743.260 354.465 ;
        RECT 744.220 353.355 744.550 354.285 ;
        RECT 743.090 353.185 744.550 353.355 ;
        RECT 743.090 352.685 743.420 353.185 ;
        RECT 743.770 352.005 744.100 352.980 ;
        RECT 742.640 351.325 742.970 351.825 ;
        RECT 744.280 351.325 744.550 353.185 ;
        RECT 747.195 351.465 747.530 354.535 ;
        RECT 748.835 352.805 749.085 353.805 ;
        RECT 750.340 353.505 750.590 353.975 ;
        RECT 752.750 353.645 753.000 354.555 ;
        RECT 754.820 354.435 755.850 354.605 ;
        RECT 754.820 354.075 754.990 354.435 ;
        RECT 747.710 352.475 749.085 352.805 ;
        RECT 748.875 352.295 749.085 352.475 ;
        RECT 749.585 353.335 750.590 353.505 ;
        RECT 752.125 353.475 753.000 353.645 ;
        RECT 753.180 353.905 754.990 354.075 ;
        RECT 749.585 352.805 749.755 353.335 ;
        RECT 752.125 353.155 752.295 353.475 ;
        RECT 749.935 352.985 752.295 353.155 ;
        RECT 749.585 352.635 751.625 352.805 ;
        RECT 748.875 351.795 749.205 352.295 ;
        RECT 749.585 351.795 749.810 352.635 ;
        RECT 751.295 352.245 751.625 352.635 ;
        RECT 749.480 351.295 749.810 351.795 ;
        RECT 751.830 351.585 752.000 352.985 ;
        RECT 752.475 352.735 752.805 353.235 ;
        RECT 753.180 352.555 753.350 353.905 ;
        RECT 752.180 352.385 753.350 352.555 ;
        RECT 753.530 353.145 753.860 353.725 ;
        RECT 755.170 353.495 755.500 354.255 ;
        RECT 755.680 353.845 755.850 354.435 ;
        RECT 757.160 354.435 758.900 354.605 ;
        RECT 757.160 353.845 757.330 354.435 ;
        RECT 757.520 354.000 757.850 354.255 ;
        RECT 755.680 353.800 757.330 353.845 ;
        RECT 755.680 353.675 757.450 353.800 ;
        RECT 755.170 353.325 756.940 353.495 ;
        RECT 757.120 353.480 757.450 353.675 ;
        RECT 756.770 353.300 756.940 353.325 ;
        RECT 757.630 353.300 757.800 354.000 ;
        RECT 753.530 352.975 756.590 353.145 ;
        RECT 752.180 351.885 752.465 352.385 ;
        RECT 753.530 352.125 753.790 352.975 ;
        RECT 756.260 352.625 756.590 352.975 ;
        RECT 756.770 353.130 757.800 353.300 ;
        RECT 757.980 353.470 758.200 353.800 ;
        RECT 758.380 353.640 758.550 354.255 ;
        RECT 758.730 353.990 758.900 354.435 ;
        RECT 759.590 354.435 761.030 354.605 ;
        RECT 759.590 353.990 759.760 354.435 ;
        RECT 758.730 353.820 759.760 353.990 ;
        RECT 759.940 353.640 760.190 354.255 ;
        RECT 758.380 353.470 760.190 353.640 ;
        RECT 756.770 352.445 756.940 353.130 ;
        RECT 757.980 352.950 758.150 353.470 ;
        RECT 758.380 353.290 758.550 353.470 ;
        RECT 754.320 352.275 756.940 352.445 ;
        RECT 752.670 351.585 753.000 352.125 ;
        RECT 751.830 351.415 753.000 351.585 ;
        RECT 753.460 351.415 753.790 352.125 ;
        RECT 756.770 352.045 756.940 352.275 ;
        RECT 757.125 352.720 758.150 352.950 ;
        RECT 758.330 353.120 758.550 353.290 ;
        RECT 757.125 352.225 757.455 352.720 ;
        RECT 758.330 352.125 758.500 353.120 ;
        RECT 760.430 352.950 760.680 354.255 ;
        RECT 756.770 351.875 757.780 352.045 ;
        RECT 757.450 351.625 757.780 351.875 ;
        RECT 758.230 351.625 758.500 352.125 ;
        RECT 758.685 351.840 759.015 352.905 ;
        RECT 760.155 352.720 760.680 352.950 ;
        RECT 758.685 351.610 759.020 351.840 ;
        RECT 760.410 351.795 760.680 352.720 ;
        RECT 760.860 353.325 761.030 354.435 ;
        RECT 761.990 353.325 762.320 354.255 ;
        RECT 760.860 353.155 762.320 353.325 ;
        RECT 760.860 352.655 761.190 353.155 ;
        RECT 761.540 351.975 761.870 352.950 ;
        RECT 760.410 351.295 760.740 351.795 ;
        RECT 762.050 351.295 762.320 353.155 ;
        RECT 765.235 351.385 765.570 354.455 ;
        RECT 766.875 352.725 767.125 353.725 ;
        RECT 768.380 353.425 768.630 353.895 ;
        RECT 770.790 353.565 771.040 354.475 ;
        RECT 772.860 354.355 773.890 354.525 ;
        RECT 772.860 353.995 773.030 354.355 ;
        RECT 765.750 352.395 767.125 352.725 ;
        RECT 766.915 352.215 767.125 352.395 ;
        RECT 767.625 353.255 768.630 353.425 ;
        RECT 770.165 353.395 771.040 353.565 ;
        RECT 771.220 353.825 773.030 353.995 ;
        RECT 767.625 352.725 767.795 353.255 ;
        RECT 770.165 353.075 770.335 353.395 ;
        RECT 767.975 352.905 770.335 353.075 ;
        RECT 767.625 352.555 769.665 352.725 ;
        RECT 766.915 351.715 767.245 352.215 ;
        RECT 767.625 351.715 767.850 352.555 ;
        RECT 769.335 352.165 769.665 352.555 ;
        RECT 767.520 351.215 767.850 351.715 ;
        RECT 769.870 351.505 770.040 352.905 ;
        RECT 770.515 352.655 770.845 353.155 ;
        RECT 771.220 352.475 771.390 353.825 ;
        RECT 770.220 352.305 771.390 352.475 ;
        RECT 771.570 353.065 771.900 353.645 ;
        RECT 773.210 353.415 773.540 354.175 ;
        RECT 773.720 353.765 773.890 354.355 ;
        RECT 775.200 354.355 776.940 354.525 ;
        RECT 775.200 353.765 775.370 354.355 ;
        RECT 775.560 353.920 775.890 354.175 ;
        RECT 773.720 353.720 775.370 353.765 ;
        RECT 773.720 353.595 775.490 353.720 ;
        RECT 773.210 353.245 774.980 353.415 ;
        RECT 775.160 353.400 775.490 353.595 ;
        RECT 774.810 353.220 774.980 353.245 ;
        RECT 775.670 353.220 775.840 353.920 ;
        RECT 771.570 352.895 774.630 353.065 ;
        RECT 770.220 351.805 770.505 352.305 ;
        RECT 771.570 352.045 771.830 352.895 ;
        RECT 774.300 352.545 774.630 352.895 ;
        RECT 774.810 353.050 775.840 353.220 ;
        RECT 776.020 353.390 776.240 353.720 ;
        RECT 776.420 353.560 776.590 354.175 ;
        RECT 776.770 353.910 776.940 354.355 ;
        RECT 777.630 354.355 779.070 354.525 ;
        RECT 777.630 353.910 777.800 354.355 ;
        RECT 776.770 353.740 777.800 353.910 ;
        RECT 777.980 353.560 778.230 354.175 ;
        RECT 776.420 353.390 778.230 353.560 ;
        RECT 774.810 352.365 774.980 353.050 ;
        RECT 776.020 352.870 776.190 353.390 ;
        RECT 776.420 353.210 776.590 353.390 ;
        RECT 772.360 352.195 774.980 352.365 ;
        RECT 770.710 351.505 771.040 352.045 ;
        RECT 769.870 351.335 771.040 351.505 ;
        RECT 771.500 351.335 771.830 352.045 ;
        RECT 774.810 351.965 774.980 352.195 ;
        RECT 775.165 352.640 776.190 352.870 ;
        RECT 776.370 353.040 776.590 353.210 ;
        RECT 775.165 352.145 775.495 352.640 ;
        RECT 776.370 352.045 776.540 353.040 ;
        RECT 778.470 352.870 778.720 354.175 ;
        RECT 774.810 351.795 775.820 351.965 ;
        RECT 775.490 351.545 775.820 351.795 ;
        RECT 776.270 351.545 776.540 352.045 ;
        RECT 776.725 351.530 777.055 352.825 ;
        RECT 778.195 352.640 778.720 352.870 ;
        RECT 778.450 351.715 778.720 352.640 ;
        RECT 778.900 353.245 779.070 354.355 ;
        RECT 780.030 353.245 780.360 354.175 ;
        RECT 778.900 353.075 780.360 353.245 ;
        RECT 778.900 352.575 779.230 353.075 ;
        RECT 779.580 351.895 779.910 352.870 ;
        RECT 778.450 351.215 778.780 351.715 ;
        RECT 780.090 351.215 780.360 353.075 ;
        RECT 783.395 351.425 783.730 354.495 ;
        RECT 785.035 352.765 785.285 353.765 ;
        RECT 786.540 353.465 786.790 353.935 ;
        RECT 788.950 353.605 789.200 354.515 ;
        RECT 791.020 354.395 792.050 354.565 ;
        RECT 791.020 354.035 791.190 354.395 ;
        RECT 783.910 352.435 785.285 352.765 ;
        RECT 785.075 352.255 785.285 352.435 ;
        RECT 785.785 353.295 786.790 353.465 ;
        RECT 788.325 353.435 789.200 353.605 ;
        RECT 789.380 353.865 791.190 354.035 ;
        RECT 785.785 352.765 785.955 353.295 ;
        RECT 788.325 353.115 788.495 353.435 ;
        RECT 786.135 352.945 788.495 353.115 ;
        RECT 785.785 352.595 787.825 352.765 ;
        RECT 785.075 351.755 785.405 352.255 ;
        RECT 785.785 351.755 786.010 352.595 ;
        RECT 787.495 352.205 787.825 352.595 ;
        RECT 785.680 351.255 786.010 351.755 ;
        RECT 788.030 351.545 788.200 352.945 ;
        RECT 788.675 352.695 789.005 353.195 ;
        RECT 789.380 352.515 789.550 353.865 ;
        RECT 788.380 352.345 789.550 352.515 ;
        RECT 789.730 353.105 790.060 353.685 ;
        RECT 791.370 353.455 791.700 354.215 ;
        RECT 791.880 353.805 792.050 354.395 ;
        RECT 793.360 354.395 795.100 354.565 ;
        RECT 793.360 353.805 793.530 354.395 ;
        RECT 793.720 353.960 794.050 354.215 ;
        RECT 791.880 353.760 793.530 353.805 ;
        RECT 791.880 353.635 793.650 353.760 ;
        RECT 791.370 353.285 793.140 353.455 ;
        RECT 793.320 353.440 793.650 353.635 ;
        RECT 792.970 353.260 793.140 353.285 ;
        RECT 793.830 353.260 794.000 353.960 ;
        RECT 789.730 352.935 792.790 353.105 ;
        RECT 788.380 351.845 788.665 352.345 ;
        RECT 789.730 352.085 789.990 352.935 ;
        RECT 792.460 352.585 792.790 352.935 ;
        RECT 792.970 353.090 794.000 353.260 ;
        RECT 794.180 353.430 794.400 353.760 ;
        RECT 794.580 353.600 794.750 354.215 ;
        RECT 794.930 353.950 795.100 354.395 ;
        RECT 795.790 354.395 797.230 354.565 ;
        RECT 795.790 353.950 795.960 354.395 ;
        RECT 794.930 353.780 795.960 353.950 ;
        RECT 796.140 353.600 796.390 354.215 ;
        RECT 794.580 353.430 796.390 353.600 ;
        RECT 792.970 352.405 793.140 353.090 ;
        RECT 794.180 352.910 794.350 353.430 ;
        RECT 794.580 353.250 794.750 353.430 ;
        RECT 790.520 352.235 793.140 352.405 ;
        RECT 788.870 351.545 789.200 352.085 ;
        RECT 788.030 351.375 789.200 351.545 ;
        RECT 789.660 351.375 789.990 352.085 ;
        RECT 792.970 352.005 793.140 352.235 ;
        RECT 793.325 352.680 794.350 352.910 ;
        RECT 794.530 353.080 794.750 353.250 ;
        RECT 793.325 352.185 793.655 352.680 ;
        RECT 794.530 352.085 794.700 353.080 ;
        RECT 796.630 352.910 796.880 354.215 ;
        RECT 792.970 351.835 793.980 352.005 ;
        RECT 793.650 351.585 793.980 351.835 ;
        RECT 794.430 351.585 794.700 352.085 ;
        RECT 794.885 351.570 795.215 352.865 ;
        RECT 796.355 352.680 796.880 352.910 ;
        RECT 796.610 351.755 796.880 352.680 ;
        RECT 797.060 353.285 797.230 354.395 ;
        RECT 798.190 353.285 798.520 354.215 ;
        RECT 797.060 353.115 798.520 353.285 ;
        RECT 797.060 352.615 797.390 353.115 ;
        RECT 797.740 352.860 798.070 352.910 ;
        RECT 797.730 352.490 798.070 352.860 ;
        RECT 797.740 351.935 798.070 352.490 ;
        RECT 796.610 351.255 796.940 351.755 ;
        RECT 798.250 351.255 798.520 353.115 ;
        RECT 801.775 351.435 802.110 354.505 ;
        RECT 803.415 352.775 803.665 353.775 ;
        RECT 804.920 353.475 805.170 353.945 ;
        RECT 807.330 353.615 807.580 354.525 ;
        RECT 809.400 354.405 810.430 354.575 ;
        RECT 809.400 354.045 809.570 354.405 ;
        RECT 802.290 352.445 803.665 352.775 ;
        RECT 803.455 352.265 803.665 352.445 ;
        RECT 804.165 353.305 805.170 353.475 ;
        RECT 806.705 353.445 807.580 353.615 ;
        RECT 807.760 353.875 809.570 354.045 ;
        RECT 804.165 352.775 804.335 353.305 ;
        RECT 806.705 353.125 806.875 353.445 ;
        RECT 804.515 352.955 806.875 353.125 ;
        RECT 804.165 352.605 806.205 352.775 ;
        RECT 803.455 351.765 803.785 352.265 ;
        RECT 804.165 351.765 804.390 352.605 ;
        RECT 805.875 352.215 806.205 352.605 ;
        RECT 804.060 351.265 804.390 351.765 ;
        RECT 806.410 351.555 806.580 352.955 ;
        RECT 807.055 352.705 807.385 353.205 ;
        RECT 807.760 352.525 807.930 353.875 ;
        RECT 806.760 352.355 807.930 352.525 ;
        RECT 808.110 353.115 808.440 353.695 ;
        RECT 809.750 353.465 810.080 354.225 ;
        RECT 810.260 353.815 810.430 354.405 ;
        RECT 811.740 354.405 813.480 354.575 ;
        RECT 811.740 353.815 811.910 354.405 ;
        RECT 812.100 353.970 812.430 354.225 ;
        RECT 810.260 353.770 811.910 353.815 ;
        RECT 810.260 353.645 812.030 353.770 ;
        RECT 809.750 353.295 811.520 353.465 ;
        RECT 811.700 353.450 812.030 353.645 ;
        RECT 811.350 353.270 811.520 353.295 ;
        RECT 812.210 353.270 812.380 353.970 ;
        RECT 808.110 352.945 811.170 353.115 ;
        RECT 806.760 351.855 807.045 352.355 ;
        RECT 808.110 352.095 808.370 352.945 ;
        RECT 810.840 352.595 811.170 352.945 ;
        RECT 811.350 353.100 812.380 353.270 ;
        RECT 812.560 353.440 812.780 353.770 ;
        RECT 812.960 353.610 813.130 354.225 ;
        RECT 813.310 353.960 813.480 354.405 ;
        RECT 814.170 354.405 815.610 354.575 ;
        RECT 814.170 353.960 814.340 354.405 ;
        RECT 813.310 353.790 814.340 353.960 ;
        RECT 814.520 353.610 814.770 354.225 ;
        RECT 812.960 353.440 814.770 353.610 ;
        RECT 811.350 352.415 811.520 353.100 ;
        RECT 812.560 352.920 812.730 353.440 ;
        RECT 812.960 353.260 813.130 353.440 ;
        RECT 808.900 352.245 811.520 352.415 ;
        RECT 807.250 351.555 807.580 352.095 ;
        RECT 806.410 351.385 807.580 351.555 ;
        RECT 808.040 351.385 808.370 352.095 ;
        RECT 811.350 352.015 811.520 352.245 ;
        RECT 811.705 352.690 812.730 352.920 ;
        RECT 812.910 353.090 813.130 353.260 ;
        RECT 811.705 352.195 812.035 352.690 ;
        RECT 812.910 352.095 813.080 353.090 ;
        RECT 815.010 352.920 815.260 354.225 ;
        RECT 811.350 351.845 812.360 352.015 ;
        RECT 812.030 351.595 812.360 351.845 ;
        RECT 812.810 351.595 813.080 352.095 ;
        RECT 813.265 351.580 813.595 352.875 ;
        RECT 814.735 352.690 815.260 352.920 ;
        RECT 814.990 351.765 815.260 352.690 ;
        RECT 815.440 353.295 815.610 354.405 ;
        RECT 816.570 353.295 816.900 354.225 ;
        RECT 815.440 353.125 816.900 353.295 ;
        RECT 815.440 352.625 815.770 353.125 ;
        RECT 816.120 351.945 816.450 352.920 ;
        RECT 814.990 351.265 815.320 351.765 ;
        RECT 816.630 351.265 816.900 353.125 ;
        RECT 818.540 351.610 819.530 352.340 ;
        RECT 385.700 350.240 386.490 350.260 ;
        RECT 379.060 349.930 386.490 350.240 ;
        RECT 379.060 349.900 379.360 349.930 ;
        RECT 385.610 349.910 386.000 349.930 ;
        RECT 385.700 349.890 386.000 349.910 ;
        RECT 656.060 349.530 656.690 350.290 ;
        RECT 818.740 347.710 819.530 351.610 ;
        RECT 820.575 351.415 820.910 354.485 ;
        RECT 822.215 352.755 822.465 353.755 ;
        RECT 823.720 353.455 823.970 353.925 ;
        RECT 826.130 353.595 826.380 354.505 ;
        RECT 828.200 354.385 829.230 354.555 ;
        RECT 828.200 354.025 828.370 354.385 ;
        RECT 821.090 352.425 822.465 352.755 ;
        RECT 822.255 352.245 822.465 352.425 ;
        RECT 822.965 353.285 823.970 353.455 ;
        RECT 825.505 353.425 826.380 353.595 ;
        RECT 826.560 353.855 828.370 354.025 ;
        RECT 822.965 352.755 823.135 353.285 ;
        RECT 825.505 353.105 825.675 353.425 ;
        RECT 823.315 352.935 825.675 353.105 ;
        RECT 822.965 352.585 825.005 352.755 ;
        RECT 822.255 351.745 822.585 352.245 ;
        RECT 822.965 351.745 823.190 352.585 ;
        RECT 824.025 352.015 824.355 352.405 ;
        RECT 824.675 352.195 825.005 352.585 ;
        RECT 824.025 351.845 825.030 352.015 ;
        RECT 822.860 351.245 823.190 351.745 ;
        RECT 824.860 351.185 825.030 351.845 ;
        RECT 825.210 351.535 825.380 352.935 ;
        RECT 825.855 352.685 826.185 353.185 ;
        RECT 826.560 352.505 826.730 353.855 ;
        RECT 825.560 352.335 826.730 352.505 ;
        RECT 826.910 353.095 827.240 353.675 ;
        RECT 828.550 353.445 828.880 354.205 ;
        RECT 829.060 353.795 829.230 354.385 ;
        RECT 830.540 354.385 832.280 354.555 ;
        RECT 830.540 353.795 830.710 354.385 ;
        RECT 830.900 353.950 831.230 354.205 ;
        RECT 829.060 353.750 830.710 353.795 ;
        RECT 829.060 353.625 830.830 353.750 ;
        RECT 828.550 353.275 830.320 353.445 ;
        RECT 830.500 353.430 830.830 353.625 ;
        RECT 830.150 353.250 830.320 353.275 ;
        RECT 831.010 353.250 831.180 353.950 ;
        RECT 826.910 352.925 829.970 353.095 ;
        RECT 825.560 351.835 825.845 352.335 ;
        RECT 826.910 352.075 827.170 352.925 ;
        RECT 826.050 351.535 826.380 352.075 ;
        RECT 825.210 351.365 826.380 351.535 ;
        RECT 826.840 351.365 827.170 352.075 ;
        RECT 827.350 352.575 829.205 352.745 ;
        RECT 829.640 352.575 829.970 352.925 ;
        RECT 830.150 353.080 831.180 353.250 ;
        RECT 831.360 353.420 831.580 353.750 ;
        RECT 831.760 353.590 831.930 354.205 ;
        RECT 832.110 353.940 832.280 354.385 ;
        RECT 832.970 354.385 834.410 354.555 ;
        RECT 832.970 353.940 833.140 354.385 ;
        RECT 832.110 353.770 833.140 353.940 ;
        RECT 833.320 353.590 833.570 354.205 ;
        RECT 831.760 353.420 833.570 353.590 ;
        RECT 827.350 352.045 827.520 352.575 ;
        RECT 830.150 352.395 830.320 353.080 ;
        RECT 831.360 352.900 831.530 353.420 ;
        RECT 831.760 353.240 831.930 353.420 ;
        RECT 827.700 352.225 830.320 352.395 ;
        RECT 827.350 351.875 829.970 352.045 ;
        RECT 827.350 351.185 827.520 351.875 ;
        RECT 828.970 351.730 829.320 351.875 ;
        RECT 829.800 351.380 829.970 351.875 ;
        RECT 830.150 351.995 830.320 352.225 ;
        RECT 830.505 352.670 831.530 352.900 ;
        RECT 831.710 353.070 831.930 353.240 ;
        RECT 830.505 352.175 830.835 352.670 ;
        RECT 831.710 352.075 831.880 353.070 ;
        RECT 830.150 351.825 831.160 351.995 ;
        RECT 830.830 351.575 831.160 351.825 ;
        RECT 831.610 351.575 831.880 352.075 ;
        RECT 832.575 352.370 833.115 353.240 ;
        RECT 833.810 352.900 834.060 354.205 ;
        RECT 833.535 352.670 834.060 352.900 ;
        RECT 832.575 351.380 832.745 352.370 ;
        RECT 829.800 351.210 832.745 351.380 ;
        RECT 833.790 351.745 834.060 352.670 ;
        RECT 834.240 353.275 834.410 354.385 ;
        RECT 835.370 353.275 835.700 354.205 ;
        RECT 834.240 353.105 835.700 353.275 ;
        RECT 834.240 352.605 834.570 353.105 ;
        RECT 834.920 351.925 835.250 352.900 ;
        RECT 833.790 351.245 834.120 351.745 ;
        RECT 835.430 351.245 835.700 353.105 ;
        RECT 839.015 352.905 839.400 354.485 ;
        RECT 839.015 352.640 839.345 352.905 ;
        RECT 838.040 352.260 839.345 352.640 ;
        RECT 836.110 351.290 836.770 351.870 ;
        RECT 824.860 351.015 827.520 351.185 ;
        RECT 832.110 349.180 834.130 349.470 ;
        RECT 836.190 349.180 836.580 351.290 ;
        RECT 839.015 351.225 839.345 352.260 ;
        RECT 832.110 348.600 836.630 349.180 ;
        RECT 832.110 348.360 834.210 348.600 ;
        RECT 832.110 348.030 834.130 348.360 ;
        RECT 837.430 347.710 838.740 348.300 ;
        RECT 818.700 347.270 838.740 347.710 ;
        RECT 818.700 347.110 837.950 347.270 ;
        RECT 379.140 346.570 379.310 346.730 ;
        RECT 379.090 332.570 379.370 346.570 ;
        RECT 385.720 346.340 385.890 346.730 ;
        RECT 379.040 332.350 379.370 332.570 ;
        RECT 385.660 332.560 385.940 346.340 ;
        RECT 780.120 344.370 781.000 344.730 ;
        RECT 783.935 344.380 784.210 346.345 ;
        RECT 785.820 344.665 785.990 345.265 ;
        RECT 790.485 344.795 790.870 346.375 ;
        RECT 783.200 344.370 784.210 344.380 ;
        RECT 780.120 344.070 784.210 344.370 ;
        RECT 784.415 344.495 786.475 344.665 ;
        RECT 784.415 344.315 784.745 344.495 ;
        RECT 780.120 344.050 783.740 344.070 ;
        RECT 780.120 343.390 781.000 344.050 ;
        RECT 783.935 343.085 784.210 344.070 ;
        RECT 785.735 343.400 786.125 344.315 ;
        RECT 786.305 343.585 786.475 344.495 ;
        RECT 786.655 344.300 787.065 344.435 ;
        RECT 790.485 344.300 790.815 344.795 ;
        RECT 786.655 344.080 790.815 344.300 ;
        RECT 790.995 344.460 791.705 344.555 ;
        RECT 793.975 344.460 794.310 346.415 ;
        RECT 795.615 344.685 795.865 345.685 ;
        RECT 797.120 345.385 797.370 345.855 ;
        RECT 799.530 345.525 799.780 346.435 ;
        RECT 801.600 346.315 802.630 346.485 ;
        RECT 801.600 345.955 801.770 346.315 ;
        RECT 790.995 344.230 794.310 344.460 ;
        RECT 794.490 344.355 795.865 344.685 ;
        RECT 790.995 344.170 791.705 344.230 ;
        RECT 786.655 343.765 787.065 344.080 ;
        RECT 786.305 343.415 787.060 343.585 ;
        RECT 786.810 343.085 787.060 343.415 ;
        RECT 790.485 343.115 790.815 344.080 ;
        RECT 793.975 343.345 794.310 344.230 ;
        RECT 795.655 344.175 795.865 344.355 ;
        RECT 796.365 345.215 797.370 345.385 ;
        RECT 798.905 345.355 799.780 345.525 ;
        RECT 799.960 345.785 801.770 345.955 ;
        RECT 796.365 344.685 796.535 345.215 ;
        RECT 798.905 345.035 799.075 345.355 ;
        RECT 796.715 344.865 799.075 345.035 ;
        RECT 796.365 344.515 798.405 344.685 ;
        RECT 795.655 343.675 795.985 344.175 ;
        RECT 796.365 343.675 796.590 344.515 ;
        RECT 798.075 344.125 798.405 344.515 ;
        RECT 796.260 343.175 796.590 343.675 ;
        RECT 798.610 343.465 798.780 344.865 ;
        RECT 799.255 344.615 799.585 345.115 ;
        RECT 799.960 344.435 800.130 345.785 ;
        RECT 798.960 344.265 800.130 344.435 ;
        RECT 800.310 345.025 800.640 345.605 ;
        RECT 801.950 345.375 802.280 346.135 ;
        RECT 802.460 345.725 802.630 346.315 ;
        RECT 803.940 346.315 805.680 346.485 ;
        RECT 803.940 345.725 804.110 346.315 ;
        RECT 804.300 345.880 804.630 346.135 ;
        RECT 802.460 345.680 804.110 345.725 ;
        RECT 802.460 345.555 804.230 345.680 ;
        RECT 801.950 345.205 803.720 345.375 ;
        RECT 803.900 345.360 804.230 345.555 ;
        RECT 803.550 345.180 803.720 345.205 ;
        RECT 804.410 345.180 804.580 345.880 ;
        RECT 800.310 344.855 803.370 345.025 ;
        RECT 798.960 343.765 799.245 344.265 ;
        RECT 800.310 344.005 800.570 344.855 ;
        RECT 803.040 344.505 803.370 344.855 ;
        RECT 803.550 345.010 804.580 345.180 ;
        RECT 804.760 345.350 804.980 345.680 ;
        RECT 805.160 345.520 805.330 346.135 ;
        RECT 805.510 345.870 805.680 346.315 ;
        RECT 806.370 346.315 807.810 346.485 ;
        RECT 806.370 345.870 806.540 346.315 ;
        RECT 805.510 345.700 806.540 345.870 ;
        RECT 806.720 345.520 806.970 346.135 ;
        RECT 805.160 345.350 806.970 345.520 ;
        RECT 803.550 344.325 803.720 345.010 ;
        RECT 804.760 344.830 804.930 345.350 ;
        RECT 805.160 345.170 805.330 345.350 ;
        RECT 801.100 344.155 803.720 344.325 ;
        RECT 799.450 343.465 799.780 344.005 ;
        RECT 798.610 343.295 799.780 343.465 ;
        RECT 800.240 343.295 800.570 344.005 ;
        RECT 803.550 343.925 803.720 344.155 ;
        RECT 803.905 344.600 804.930 344.830 ;
        RECT 805.110 345.000 805.330 345.170 ;
        RECT 803.905 344.105 804.235 344.600 ;
        RECT 805.110 344.005 805.280 345.000 ;
        RECT 807.210 344.830 807.460 346.135 ;
        RECT 803.550 343.755 804.560 343.925 ;
        RECT 804.230 343.505 804.560 343.755 ;
        RECT 805.010 343.505 805.280 344.005 ;
        RECT 805.465 343.490 805.795 344.785 ;
        RECT 806.935 344.600 807.460 344.830 ;
        RECT 807.190 343.675 807.460 344.600 ;
        RECT 807.640 345.205 807.810 346.315 ;
        RECT 808.770 345.205 809.100 346.135 ;
        RECT 813.335 345.530 813.670 346.325 ;
        RECT 813.320 345.230 813.680 345.530 ;
        RECT 807.640 345.035 809.100 345.205 ;
        RECT 807.640 344.535 807.970 345.035 ;
        RECT 807.190 343.175 807.520 343.675 ;
        RECT 808.830 343.175 809.100 345.035 ;
        RECT 813.335 343.255 813.670 345.230 ;
        RECT 814.975 344.595 815.225 345.595 ;
        RECT 816.480 345.295 816.730 345.765 ;
        RECT 818.890 345.435 819.140 346.345 ;
        RECT 820.960 346.225 821.990 346.395 ;
        RECT 820.960 345.865 821.130 346.225 ;
        RECT 813.850 344.265 815.225 344.595 ;
        RECT 815.015 344.085 815.225 344.265 ;
        RECT 815.725 345.125 816.730 345.295 ;
        RECT 818.265 345.265 819.140 345.435 ;
        RECT 819.320 345.695 821.130 345.865 ;
        RECT 815.725 344.595 815.895 345.125 ;
        RECT 818.265 344.945 818.435 345.265 ;
        RECT 816.075 344.775 818.435 344.945 ;
        RECT 815.725 344.425 817.765 344.595 ;
        RECT 815.015 343.585 815.345 344.085 ;
        RECT 815.725 343.585 815.950 344.425 ;
        RECT 817.435 344.035 817.765 344.425 ;
        RECT 815.620 343.085 815.950 343.585 ;
        RECT 817.970 343.375 818.140 344.775 ;
        RECT 818.615 344.525 818.945 345.025 ;
        RECT 819.320 344.345 819.490 345.695 ;
        RECT 818.320 344.175 819.490 344.345 ;
        RECT 819.670 344.935 820.000 345.515 ;
        RECT 821.310 345.285 821.640 346.045 ;
        RECT 821.820 345.635 821.990 346.225 ;
        RECT 823.300 346.225 825.040 346.395 ;
        RECT 823.300 345.635 823.470 346.225 ;
        RECT 823.660 345.790 823.990 346.045 ;
        RECT 821.820 345.590 823.470 345.635 ;
        RECT 821.820 345.465 823.590 345.590 ;
        RECT 821.310 345.115 823.080 345.285 ;
        RECT 823.260 345.270 823.590 345.465 ;
        RECT 822.910 345.090 823.080 345.115 ;
        RECT 823.770 345.090 823.940 345.790 ;
        RECT 819.670 344.765 822.730 344.935 ;
        RECT 818.320 343.675 818.605 344.175 ;
        RECT 819.670 343.915 819.930 344.765 ;
        RECT 822.400 344.415 822.730 344.765 ;
        RECT 822.910 344.920 823.940 345.090 ;
        RECT 824.120 345.260 824.340 345.590 ;
        RECT 824.520 345.430 824.690 346.045 ;
        RECT 824.870 345.780 825.040 346.225 ;
        RECT 825.730 346.225 827.170 346.395 ;
        RECT 825.730 345.780 825.900 346.225 ;
        RECT 824.870 345.610 825.900 345.780 ;
        RECT 826.080 345.430 826.330 346.045 ;
        RECT 824.520 345.260 826.330 345.430 ;
        RECT 822.910 344.235 823.080 344.920 ;
        RECT 824.120 344.740 824.290 345.260 ;
        RECT 824.520 345.080 824.690 345.260 ;
        RECT 820.460 344.065 823.080 344.235 ;
        RECT 818.810 343.375 819.140 343.915 ;
        RECT 817.970 343.205 819.140 343.375 ;
        RECT 819.600 343.205 819.930 343.915 ;
        RECT 822.910 343.835 823.080 344.065 ;
        RECT 823.265 344.510 824.290 344.740 ;
        RECT 824.470 344.910 824.690 345.080 ;
        RECT 823.265 344.015 823.595 344.510 ;
        RECT 824.470 343.915 824.640 344.910 ;
        RECT 826.570 344.740 826.820 346.045 ;
        RECT 822.910 343.665 823.920 343.835 ;
        RECT 823.590 343.415 823.920 343.665 ;
        RECT 824.370 343.415 824.640 343.915 ;
        RECT 824.825 343.400 825.155 344.695 ;
        RECT 826.295 344.510 826.820 344.740 ;
        RECT 826.550 343.585 826.820 344.510 ;
        RECT 827.000 345.115 827.170 346.225 ;
        RECT 828.130 345.115 828.460 346.045 ;
        RECT 870.600 345.690 871.940 347.950 ;
        RECT 827.000 344.945 828.460 345.115 ;
        RECT 827.000 344.445 827.330 344.945 ;
        RECT 826.550 343.085 826.880 343.585 ;
        RECT 828.190 343.085 828.460 344.945 ;
        RECT 865.730 341.690 866.540 341.760 ;
        RECT 846.150 341.660 866.540 341.690 ;
        RECT 844.580 341.000 866.540 341.660 ;
        RECT 632.020 333.330 633.420 334.450 ;
        RECT 844.580 332.640 845.130 341.000 ;
        RECT 853.410 338.540 854.490 339.280 ;
        RECT 852.620 337.520 852.790 337.940 ;
        RECT 855.200 337.520 855.370 337.940 ;
        RECT 852.620 336.050 852.790 336.470 ;
        RECT 855.200 336.050 855.370 336.470 ;
        RECT 852.620 334.580 852.790 335.000 ;
        RECT 855.200 334.580 855.370 335.000 ;
        RECT 865.730 334.410 866.540 341.000 ;
        RECT 865.730 333.680 866.550 334.410 ;
        RECT 852.620 333.110 852.790 333.530 ;
        RECT 855.200 333.110 855.370 333.530 ;
        RECT 379.040 331.360 379.340 332.350 ;
        RECT 385.660 332.120 385.980 332.560 ;
        RECT 844.600 332.510 845.130 332.640 ;
        RECT 385.680 331.380 385.980 332.120 ;
        RECT 603.420 332.050 603.590 332.470 ;
        RECT 605.000 332.050 605.170 332.470 ;
        RECT 607.940 332.060 608.110 332.480 ;
        RECT 609.520 332.060 609.690 332.480 ;
        RECT 612.460 332.060 612.630 332.480 ;
        RECT 614.040 332.060 614.210 332.480 ;
        RECT 616.890 332.040 617.060 332.460 ;
        RECT 618.470 332.040 618.640 332.460 ;
        RECT 621.270 332.050 621.440 332.470 ;
        RECT 622.850 332.050 623.020 332.470 ;
        RECT 625.590 332.040 625.760 332.460 ;
        RECT 627.170 332.040 627.340 332.460 ;
        RECT 385.680 331.360 386.470 331.380 ;
        RECT 379.040 331.050 386.470 331.360 ;
        RECT 379.040 331.020 379.340 331.050 ;
        RECT 385.680 331.010 385.980 331.050 ;
        RECT 603.420 330.580 603.590 331.000 ;
        RECT 605.000 330.580 605.170 331.000 ;
        RECT 607.940 330.590 608.110 331.010 ;
        RECT 609.520 330.590 609.690 331.010 ;
        RECT 612.460 330.590 612.630 331.010 ;
        RECT 614.040 330.590 614.210 331.010 ;
        RECT 616.890 330.570 617.060 330.990 ;
        RECT 618.470 330.570 618.640 330.990 ;
        RECT 621.270 330.580 621.440 331.000 ;
        RECT 622.850 330.580 623.020 331.000 ;
        RECT 625.590 330.570 625.760 330.990 ;
        RECT 627.170 330.570 627.340 330.990 ;
        RECT 595.465 328.885 595.850 330.465 ;
        RECT 613.510 329.630 613.980 330.010 ;
        RECT 616.350 329.590 616.780 329.910 ;
        RECT 620.760 329.730 621.170 330.160 ;
        RECT 636.220 329.335 636.605 330.915 ;
        RECT 640.410 329.425 640.795 331.005 ;
        RECT 635.385 329.080 636.095 329.095 ;
        RECT 594.470 328.550 595.150 328.640 ;
        RECT 595.465 328.550 595.795 328.885 ;
        RECT 634.240 328.710 636.095 329.080 ;
        RECT 636.275 329.010 636.605 329.335 ;
        RECT 639.400 329.185 639.770 329.210 ;
        RECT 637.030 329.010 637.870 329.020 ;
        RECT 636.275 328.970 637.870 329.010 ;
        RECT 636.275 328.730 637.880 328.970 ;
        RECT 639.400 328.800 640.285 329.185 ;
        RECT 640.465 329.070 640.795 329.425 ;
        RECT 644.510 329.405 644.895 330.985 ;
        RECT 664.390 330.575 664.560 331.175 ;
        RECT 666.170 331.160 666.445 332.255 ;
        RECT 666.170 330.850 666.480 331.160 ;
        RECT 663.905 330.405 665.965 330.575 ;
        RECT 663.315 329.675 663.725 330.345 ;
        RECT 663.905 329.495 664.075 330.405 ;
        RECT 665.635 330.225 665.965 330.405 ;
        RECT 643.675 329.070 644.385 329.165 ;
        RECT 640.465 328.860 644.385 329.070 ;
        RECT 639.400 328.760 639.770 328.800 ;
        RECT 594.470 328.310 595.795 328.550 ;
        RECT 594.470 328.240 595.150 328.310 ;
        RECT 379.140 327.720 379.310 327.880 ;
        RECT 208.860 320.380 210.530 321.860 ;
        RECT 211.060 319.550 212.490 319.620 ;
        RECT 211.060 319.490 226.740 319.550 ;
        RECT 231.100 319.540 232.530 319.610 ;
        RECT 251.160 319.540 252.590 319.610 ;
        RECT 271.210 319.540 272.640 319.610 ;
        RECT 211.060 319.320 226.770 319.490 ;
        RECT 231.100 319.480 246.780 319.540 ;
        RECT 251.160 319.480 266.840 319.540 ;
        RECT 271.210 319.480 286.890 319.540 ;
        RECT 211.060 319.280 226.740 319.320 ;
        RECT 231.100 319.310 246.810 319.480 ;
        RECT 251.160 319.310 266.870 319.480 ;
        RECT 271.210 319.310 286.920 319.480 ;
        RECT 211.060 319.240 212.490 319.280 ;
        RECT 231.100 319.270 246.780 319.310 ;
        RECT 251.160 319.270 266.840 319.310 ;
        RECT 271.210 319.270 286.890 319.310 ;
        RECT 211.060 313.010 211.470 319.240 ;
        RECT 231.100 319.230 232.530 319.270 ;
        RECT 251.160 319.230 252.590 319.270 ;
        RECT 271.210 319.230 272.640 319.270 ;
        RECT 211.040 312.970 212.640 313.010 ;
        RECT 231.100 313.000 231.510 319.230 ;
        RECT 251.160 313.000 251.570 319.230 ;
        RECT 271.210 313.000 271.620 319.230 ;
        RECT 379.090 313.720 379.370 327.720 ;
        RECT 385.720 327.490 385.890 327.880 ;
        RECT 379.040 313.500 379.370 313.720 ;
        RECT 385.660 313.710 385.940 327.490 ;
        RECT 595.465 327.205 595.795 328.310 ;
        RECT 595.975 328.600 596.685 328.645 ;
        RECT 597.150 328.600 597.780 328.710 ;
        RECT 595.975 328.260 597.780 328.600 ;
        RECT 596.420 328.240 597.780 328.260 ;
        RECT 597.150 327.860 597.780 328.240 ;
        RECT 634.240 328.670 635.800 328.710 ;
        RECT 634.240 328.220 634.520 328.670 ;
        RECT 631.640 326.950 632.470 327.630 ;
        RECT 634.020 327.540 634.730 328.220 ;
        RECT 636.275 327.655 636.605 328.730 ;
        RECT 610.400 325.820 610.570 326.240 ;
        RECT 611.190 325.820 611.360 326.240 ;
        RECT 611.980 325.820 612.150 326.240 ;
        RECT 612.770 325.820 612.940 326.240 ;
        RECT 613.560 325.820 613.730 326.240 ;
        RECT 617.990 325.790 618.160 326.210 ;
        RECT 618.780 325.790 618.950 326.210 ;
        RECT 619.570 325.790 619.740 326.210 ;
        RECT 620.360 325.790 620.530 326.210 ;
        RECT 621.150 325.790 621.320 326.210 ;
        RECT 600.950 325.040 601.120 325.460 ;
        RECT 601.740 325.040 601.910 325.460 ;
        RECT 602.530 325.040 602.700 325.460 ;
        RECT 603.320 325.040 603.490 325.460 ;
        RECT 604.110 325.040 604.280 325.460 ;
        RECT 615.510 325.310 615.990 325.730 ;
        RECT 627.730 325.170 627.900 325.590 ;
        RECT 628.520 325.170 628.690 325.590 ;
        RECT 629.310 325.170 629.480 325.590 ;
        RECT 630.100 325.170 630.270 325.590 ;
        RECT 630.890 325.170 631.060 325.590 ;
        RECT 637.480 324.800 637.880 328.730 ;
        RECT 640.465 327.745 640.795 328.860 ;
        RECT 641.950 328.520 642.180 328.860 ;
        RECT 643.675 328.780 644.385 328.860 ;
        RECT 644.565 328.960 644.895 329.405 ;
        RECT 663.320 329.325 664.075 329.495 ;
        RECT 663.320 328.995 663.570 329.325 ;
        RECT 664.255 329.310 664.645 330.225 ;
        RECT 666.170 328.995 666.445 330.850 ;
        RECT 670.020 330.575 670.190 331.175 ;
        RECT 669.535 330.405 671.595 330.575 ;
        RECT 668.945 330.130 669.355 330.345 ;
        RECT 668.910 329.720 669.355 330.130 ;
        RECT 668.945 329.675 669.355 329.720 ;
        RECT 669.535 329.495 669.705 330.405 ;
        RECT 671.265 330.225 671.595 330.405 ;
        RECT 668.950 329.325 669.705 329.495 ;
        RECT 668.950 328.995 669.200 329.325 ;
        RECT 669.885 329.310 670.275 330.225 ;
        RECT 671.800 329.840 672.075 332.255 ;
        RECT 674.980 330.475 675.230 331.075 ;
        RECT 674.980 330.305 677.355 330.475 ;
        RECT 675.185 329.840 675.515 330.125 ;
        RECT 671.800 329.590 675.515 329.840 ;
        RECT 671.800 328.995 672.075 329.590 ;
        RECT 675.185 329.575 675.515 329.590 ;
        RECT 675.760 329.395 675.930 330.305 ;
        RECT 677.025 330.125 677.355 330.305 ;
        RECT 677.560 330.420 677.815 332.155 ;
        RECT 681.740 330.435 681.990 331.485 ;
        RECT 682.215 330.615 683.175 330.930 ;
        RECT 683.380 330.435 683.630 331.485 ;
        RECT 684.975 330.615 685.325 332.195 ;
        RECT 676.110 329.575 676.440 330.125 ;
        RECT 677.560 330.050 677.830 330.420 ;
        RECT 681.740 330.265 684.850 330.435 ;
        RECT 645.460 328.960 645.770 328.980 ;
        RECT 644.565 328.780 645.770 328.960 ;
        RECT 675.760 328.895 676.090 329.395 ;
        RECT 677.560 328.895 677.815 330.050 ;
        RECT 681.740 329.265 682.035 330.265 ;
        RECT 684.520 330.105 684.850 330.265 ;
        RECT 682.215 329.970 682.545 330.085 ;
        RECT 682.215 329.520 682.550 329.970 ;
        RECT 682.215 329.250 682.545 329.520 ;
        RECT 682.725 329.250 683.865 330.085 ;
        RECT 685.020 329.850 685.325 330.615 ;
        RECT 688.670 330.525 688.840 331.125 ;
        RECT 688.185 330.355 690.245 330.525 ;
        RECT 687.595 329.850 688.005 330.295 ;
        RECT 685.020 329.670 688.005 329.850 ;
        RECT 685.020 328.935 685.325 329.670 ;
        RECT 687.595 329.625 688.005 329.670 ;
        RECT 688.185 329.445 688.355 330.355 ;
        RECT 689.915 330.175 690.245 330.355 ;
        RECT 687.600 329.275 688.355 329.445 ;
        RECT 687.600 328.945 687.850 329.275 ;
        RECT 688.535 329.260 688.925 330.175 ;
        RECT 641.880 328.200 642.260 328.520 ;
        RECT 644.565 327.725 644.895 328.780 ;
        RECT 645.460 328.630 645.770 328.780 ;
        RECT 639.840 324.800 640.290 324.900 ;
        RECT 610.400 324.350 610.570 324.770 ;
        RECT 611.190 324.350 611.360 324.770 ;
        RECT 611.980 324.350 612.150 324.770 ;
        RECT 612.770 324.350 612.940 324.770 ;
        RECT 613.560 324.350 613.730 324.770 ;
        RECT 614.230 324.300 614.400 324.720 ;
        RECT 615.810 324.300 615.980 324.720 ;
        RECT 617.390 324.300 617.560 324.720 ;
        RECT 617.990 324.320 618.160 324.740 ;
        RECT 618.780 324.320 618.950 324.740 ;
        RECT 619.570 324.320 619.740 324.740 ;
        RECT 620.360 324.320 620.530 324.740 ;
        RECT 621.150 324.320 621.320 324.740 ;
        RECT 637.480 324.610 640.290 324.800 ;
        RECT 637.480 324.600 637.880 324.610 ;
        RECT 600.950 323.570 601.120 323.990 ;
        RECT 601.740 323.570 601.910 323.990 ;
        RECT 602.530 323.570 602.700 323.990 ;
        RECT 603.320 323.570 603.490 323.990 ;
        RECT 604.110 323.570 604.280 323.990 ;
        RECT 608.520 323.880 609.190 324.190 ;
        RECT 623.110 323.770 623.800 324.320 ;
        RECT 639.840 324.210 640.290 324.610 ;
        RECT 643.900 324.270 644.320 324.950 ;
        RECT 659.720 324.375 660.105 325.955 ;
        RECT 657.710 324.130 658.240 324.200 ;
        RECT 658.885 324.130 659.595 324.135 ;
        RECT 627.730 323.700 627.900 324.120 ;
        RECT 628.520 323.700 628.690 324.120 ;
        RECT 629.310 323.700 629.480 324.120 ;
        RECT 630.100 323.700 630.270 324.120 ;
        RECT 630.890 323.700 631.060 324.120 ;
        RECT 639.580 323.410 639.750 323.830 ;
        RECT 643.630 323.460 643.800 323.880 ;
        RECT 657.710 323.760 659.595 324.130 ;
        RECT 657.710 323.650 658.240 323.760 ;
        RECT 658.885 323.750 659.595 323.760 ;
        RECT 659.775 324.100 660.105 324.375 ;
        RECT 664.620 324.335 665.005 325.915 ;
        RECT 669.210 324.365 669.595 325.945 ;
        RECT 659.775 323.810 661.160 324.100 ;
        RECT 662.430 324.090 663.090 324.170 ;
        RECT 663.785 324.090 664.495 324.095 ;
        RECT 606.650 322.830 606.820 323.250 ;
        RECT 607.440 322.830 607.610 323.250 ;
        RECT 608.230 322.830 608.400 323.250 ;
        RECT 609.020 322.830 609.190 323.250 ;
        RECT 609.810 322.830 609.980 323.250 ;
        RECT 610.400 322.880 610.570 323.300 ;
        RECT 611.190 322.880 611.360 323.300 ;
        RECT 611.980 322.880 612.150 323.300 ;
        RECT 612.770 322.880 612.940 323.300 ;
        RECT 613.560 322.880 613.730 323.300 ;
        RECT 614.230 322.830 614.400 323.250 ;
        RECT 615.810 322.830 615.980 323.250 ;
        RECT 617.390 322.830 617.560 323.250 ;
        RECT 617.990 322.850 618.160 323.270 ;
        RECT 618.780 322.850 618.950 323.270 ;
        RECT 619.570 322.850 619.740 323.270 ;
        RECT 620.360 322.850 620.530 323.270 ;
        RECT 621.150 322.850 621.320 323.270 ;
        RECT 621.740 322.830 621.910 323.250 ;
        RECT 622.530 322.830 622.700 323.250 ;
        RECT 623.320 322.830 623.490 323.250 ;
        RECT 624.110 322.830 624.280 323.250 ;
        RECT 624.900 322.830 625.070 323.250 ;
        RECT 659.775 322.695 660.105 323.810 ;
        RECT 660.280 323.540 660.910 323.810 ;
        RECT 662.430 323.720 664.495 324.090 ;
        RECT 662.430 323.630 663.090 323.720 ;
        RECT 663.785 323.710 664.495 323.720 ;
        RECT 664.675 324.050 665.005 324.335 ;
        RECT 667.170 324.130 667.850 324.160 ;
        RECT 667.170 324.125 668.600 324.130 ;
        RECT 665.510 324.050 665.990 324.080 ;
        RECT 664.675 323.760 665.990 324.050 ;
        RECT 664.675 322.655 665.005 323.760 ;
        RECT 665.510 323.420 665.990 323.760 ;
        RECT 667.170 323.750 669.085 324.125 ;
        RECT 667.630 323.740 669.085 323.750 ;
        RECT 669.265 324.060 669.595 324.365 ;
        RECT 673.750 324.345 674.135 325.925 ;
        RECT 669.990 324.060 670.570 324.220 ;
        RECT 669.265 323.770 670.570 324.060 ;
        RECT 667.630 323.720 668.600 323.740 ;
        RECT 669.265 322.685 669.595 323.770 ;
        RECT 669.990 323.620 670.570 323.770 ;
        RECT 671.700 324.070 672.170 324.120 ;
        RECT 672.915 324.070 673.625 324.105 ;
        RECT 671.700 323.720 673.625 324.070 ;
        RECT 673.805 324.060 674.135 324.345 ;
        RECT 676.350 324.175 676.600 325.225 ;
        RECT 676.825 324.355 677.785 324.670 ;
        RECT 677.990 324.175 678.240 325.225 ;
        RECT 679.585 324.355 679.935 325.935 ;
        RECT 673.805 323.780 674.920 324.060 ;
        RECT 676.350 324.005 679.460 324.175 ;
        RECT 671.700 323.710 673.180 323.720 ;
        RECT 671.700 323.560 672.170 323.710 ;
        RECT 673.805 323.630 674.135 323.780 ;
        RECT 673.800 323.400 674.135 323.630 ;
        RECT 673.805 322.665 674.135 323.400 ;
        RECT 676.350 323.005 676.645 324.005 ;
        RECT 679.130 323.845 679.460 324.005 ;
        RECT 676.825 322.990 677.155 323.825 ;
        RECT 677.335 322.990 678.475 323.825 ;
        RECT 679.630 322.675 679.935 324.355 ;
        RECT 683.190 324.255 683.360 324.855 ;
        RECT 682.705 324.085 684.765 324.255 ;
        RECT 682.115 323.355 682.525 324.025 ;
        RECT 682.705 323.175 682.875 324.085 ;
        RECT 684.435 323.905 684.765 324.085 ;
        RECT 684.970 323.910 685.245 325.935 ;
        RECT 688.640 324.255 688.810 324.855 ;
        RECT 688.155 324.085 690.215 324.255 ;
        RECT 687.565 323.910 687.975 324.025 ;
        RECT 682.120 323.005 682.875 323.175 ;
        RECT 682.120 322.675 682.370 323.005 ;
        RECT 683.055 322.990 683.445 323.905 ;
        RECT 684.970 323.640 687.975 323.910 ;
        RECT 684.970 322.675 685.245 323.640 ;
        RECT 687.565 323.355 687.975 323.640 ;
        RECT 688.155 323.175 688.325 324.085 ;
        RECT 689.885 323.905 690.215 324.085 ;
        RECT 687.570 323.005 688.325 323.175 ;
        RECT 687.570 322.675 687.820 323.005 ;
        RECT 688.505 322.990 688.895 323.905 ;
        RECT 690.420 323.780 690.695 325.935 ;
        RECT 693.150 324.275 693.400 324.875 ;
        RECT 693.150 324.105 695.525 324.275 ;
        RECT 693.355 323.780 693.685 323.925 ;
        RECT 690.420 323.470 693.685 323.780 ;
        RECT 690.420 322.675 690.695 323.470 ;
        RECT 693.355 323.375 693.685 323.470 ;
        RECT 693.930 323.195 694.100 324.105 ;
        RECT 695.195 323.925 695.525 324.105 ;
        RECT 693.930 322.695 694.260 323.195 ;
        RECT 591.830 320.310 592.180 322.470 ;
        RECT 602.290 321.890 603.070 322.260 ;
        RECT 661.530 318.315 661.780 319.365 ;
        RECT 662.005 318.495 662.965 318.810 ;
        RECT 663.170 318.315 663.420 319.365 ;
        RECT 664.765 318.495 665.115 320.075 ;
        RECT 670.200 319.360 670.475 320.085 ;
        RECT 670.200 319.040 670.480 319.360 ;
        RECT 661.530 318.145 664.640 318.315 ;
        RECT 661.530 317.145 661.825 318.145 ;
        RECT 664.310 317.985 664.640 318.145 ;
        RECT 662.005 317.930 662.335 317.965 ;
        RECT 662.000 317.650 662.335 317.930 ;
        RECT 662.005 317.130 662.335 317.650 ;
        RECT 662.515 317.130 663.655 317.965 ;
        RECT 664.810 316.815 665.115 318.495 ;
        RECT 666.640 318.180 666.950 318.790 ;
        RECT 668.420 318.405 668.590 319.005 ;
        RECT 667.390 318.180 667.670 318.390 ;
        RECT 666.640 318.175 667.670 318.180 ;
        RECT 667.935 318.235 669.995 318.405 ;
        RECT 666.640 317.910 667.755 318.175 ;
        RECT 632.390 315.440 633.540 316.340 ;
        RECT 603.270 313.880 603.440 314.300 ;
        RECT 604.850 313.880 605.020 314.300 ;
        RECT 607.790 313.890 607.960 314.310 ;
        RECT 609.370 313.890 609.540 314.310 ;
        RECT 612.310 313.890 612.480 314.310 ;
        RECT 613.890 313.890 614.060 314.310 ;
        RECT 616.740 313.870 616.910 314.290 ;
        RECT 618.320 313.870 618.490 314.290 ;
        RECT 621.120 313.880 621.290 314.300 ;
        RECT 622.700 313.880 622.870 314.300 ;
        RECT 625.440 313.870 625.610 314.290 ;
        RECT 627.020 313.870 627.190 314.290 ;
        RECT 211.040 312.700 226.780 312.970 ;
        RECT 231.080 312.960 232.680 313.000 ;
        RECT 251.140 312.960 252.740 313.000 ;
        RECT 271.190 312.960 272.790 313.000 ;
        RECT 211.040 312.630 212.640 312.700 ;
        RECT 231.080 312.690 246.820 312.960 ;
        RECT 251.140 312.690 266.880 312.960 ;
        RECT 271.190 312.690 286.930 312.960 ;
        RECT 211.060 306.510 211.470 312.630 ;
        RECT 231.080 312.620 232.680 312.690 ;
        RECT 251.140 312.620 252.740 312.690 ;
        RECT 271.190 312.620 272.790 312.690 ;
        RECT 210.970 306.480 211.470 306.510 ;
        RECT 210.970 306.430 212.540 306.480 ;
        RECT 231.100 306.470 231.510 312.620 ;
        RECT 251.160 306.470 251.570 312.620 ;
        RECT 271.210 306.470 271.620 312.620 ;
        RECT 379.040 312.510 379.340 313.500 ;
        RECT 385.660 313.270 385.980 313.710 ;
        RECT 385.680 312.530 385.980 313.270 ;
        RECT 666.640 313.080 666.950 317.910 ;
        RECT 667.345 317.505 667.755 317.910 ;
        RECT 667.935 317.325 668.105 318.235 ;
        RECT 669.665 318.055 669.995 318.235 ;
        RECT 667.350 317.155 668.105 317.325 ;
        RECT 667.350 316.825 667.600 317.155 ;
        RECT 668.285 317.140 668.675 318.055 ;
        RECT 670.200 316.825 670.475 319.040 ;
        RECT 673.860 318.415 674.030 319.015 ;
        RECT 672.820 318.185 673.100 318.350 ;
        RECT 673.375 318.245 675.435 318.415 ;
        RECT 672.785 317.515 673.195 318.185 ;
        RECT 673.375 317.335 673.545 318.245 ;
        RECT 675.105 318.065 675.435 318.245 ;
        RECT 672.790 317.165 673.545 317.335 ;
        RECT 672.790 316.835 673.040 317.165 ;
        RECT 673.725 317.150 674.115 318.065 ;
        RECT 675.640 317.700 675.915 320.095 ;
        RECT 678.380 318.415 678.630 319.015 ;
        RECT 678.380 318.245 680.755 318.415 ;
        RECT 678.585 317.700 678.915 318.065 ;
        RECT 675.620 317.530 678.915 317.700 ;
        RECT 675.640 316.835 675.915 317.530 ;
        RECT 678.585 317.515 678.915 317.530 ;
        RECT 679.160 317.335 679.330 318.245 ;
        RECT 680.425 318.065 680.755 318.245 ;
        RECT 679.510 317.515 679.840 318.065 ;
        RECT 680.960 317.950 681.215 320.095 ;
        RECT 684.530 318.415 684.700 319.015 ;
        RECT 684.045 318.245 686.105 318.415 ;
        RECT 683.455 317.950 683.865 318.185 ;
        RECT 680.960 317.760 683.865 317.950 ;
        RECT 679.160 316.835 679.490 317.335 ;
        RECT 680.960 316.835 681.215 317.760 ;
        RECT 683.455 317.515 683.865 317.760 ;
        RECT 684.045 317.335 684.215 318.245 ;
        RECT 685.775 318.065 686.105 318.245 ;
        RECT 683.460 317.165 684.215 317.335 ;
        RECT 683.460 316.835 683.710 317.165 ;
        RECT 684.395 317.150 684.785 318.065 ;
        RECT 689.325 317.605 689.575 319.325 ;
        RECT 691.000 318.495 691.435 320.075 ;
        RECT 691.185 318.110 691.435 318.495 ;
        RECT 691.870 318.110 692.160 318.200 ;
        RECT 690.545 317.605 690.875 318.065 ;
        RECT 689.325 317.435 690.875 317.605 ;
        RECT 691.185 317.880 692.160 318.110 ;
        RECT 689.325 316.815 689.575 317.435 ;
        RECT 691.185 316.815 691.435 317.880 ;
        RECT 691.870 317.850 692.160 317.880 ;
        RECT 693.725 317.605 693.975 319.325 ;
        RECT 694.155 317.785 694.485 319.580 ;
        RECT 695.400 318.495 695.835 320.075 ;
        RECT 695.585 318.150 695.835 318.495 ;
        RECT 696.790 318.160 697.000 318.170 ;
        RECT 696.370 318.150 697.000 318.160 ;
        RECT 694.945 317.605 695.275 318.065 ;
        RECT 693.725 317.435 695.275 317.605 ;
        RECT 695.585 317.940 697.000 318.150 ;
        RECT 695.585 317.930 696.520 317.940 ;
        RECT 693.725 316.815 693.975 317.435 ;
        RECT 695.585 316.815 695.835 317.930 ;
        RECT 696.790 315.840 697.000 317.940 ;
        RECT 385.680 312.510 386.470 312.530 ;
        RECT 379.040 312.200 386.470 312.510 ;
        RECT 603.270 312.410 603.440 312.830 ;
        RECT 604.850 312.410 605.020 312.830 ;
        RECT 607.790 312.420 607.960 312.840 ;
        RECT 609.370 312.420 609.540 312.840 ;
        RECT 612.310 312.420 612.480 312.840 ;
        RECT 613.890 312.420 614.060 312.840 ;
        RECT 616.740 312.400 616.910 312.820 ;
        RECT 618.320 312.400 618.490 312.820 ;
        RECT 621.120 312.410 621.290 312.830 ;
        RECT 622.700 312.410 622.870 312.830 ;
        RECT 625.440 312.400 625.610 312.820 ;
        RECT 627.020 312.400 627.190 312.820 ;
        RECT 379.040 312.170 379.340 312.200 ;
        RECT 385.680 312.160 385.980 312.200 ;
        RECT 595.315 310.715 595.700 312.295 ;
        RECT 613.360 311.460 613.830 311.840 ;
        RECT 616.200 311.420 616.630 311.740 ;
        RECT 620.610 311.560 621.020 311.990 ;
        RECT 636.070 311.165 636.455 312.745 ;
        RECT 640.260 311.255 640.645 312.835 ;
        RECT 635.235 310.910 635.945 310.925 ;
        RECT 594.320 310.380 595.000 310.470 ;
        RECT 595.315 310.380 595.645 310.715 ;
        RECT 634.090 310.540 635.945 310.910 ;
        RECT 636.125 310.840 636.455 311.165 ;
        RECT 639.250 311.015 639.620 311.040 ;
        RECT 636.880 310.840 637.720 310.850 ;
        RECT 636.125 310.800 637.720 310.840 ;
        RECT 636.125 310.560 637.730 310.800 ;
        RECT 639.250 310.630 640.135 311.015 ;
        RECT 640.315 310.900 640.645 311.255 ;
        RECT 644.360 311.235 644.745 312.815 ;
        RECT 643.525 310.900 644.235 310.995 ;
        RECT 640.315 310.690 644.235 310.900 ;
        RECT 639.250 310.590 639.620 310.630 ;
        RECT 594.320 310.140 595.645 310.380 ;
        RECT 594.320 310.070 595.000 310.140 ;
        RECT 379.140 308.900 379.310 309.060 ;
        RECT 231.080 306.430 232.580 306.470 ;
        RECT 251.140 306.430 252.640 306.470 ;
        RECT 271.190 306.430 272.690 306.470 ;
        RECT 210.970 306.370 286.270 306.430 ;
        RECT 210.970 306.320 286.900 306.370 ;
        RECT 210.970 306.170 286.920 306.320 ;
        RECT 210.970 306.160 226.770 306.170 ;
        RECT 210.970 306.110 226.750 306.160 ;
        RECT 231.080 306.150 246.810 306.170 ;
        RECT 251.140 306.150 266.870 306.170 ;
        RECT 271.190 306.150 286.920 306.170 ;
        RECT 210.970 306.100 212.450 306.110 ;
        RECT 231.080 306.100 246.790 306.150 ;
        RECT 251.140 306.100 266.850 306.150 ;
        RECT 271.190 306.100 286.900 306.150 ;
        RECT 210.970 306.090 211.470 306.100 ;
        RECT 231.080 306.090 232.490 306.100 ;
        RECT 251.140 306.090 252.550 306.100 ;
        RECT 271.190 306.090 272.600 306.100 ;
        RECT 210.970 298.630 211.380 306.090 ;
        RECT 231.100 306.080 231.510 306.090 ;
        RECT 251.160 306.080 251.570 306.090 ;
        RECT 271.210 306.080 271.620 306.090 ;
        RECT 288.530 301.980 290.200 306.490 ;
        RECT 210.970 298.560 212.450 298.630 ;
        RECT 230.990 298.560 232.420 298.630 ;
        RECT 251.100 298.560 252.530 298.630 ;
        RECT 271.210 298.560 272.640 298.630 ;
        RECT 210.970 298.500 226.700 298.560 ;
        RECT 230.990 298.500 246.670 298.560 ;
        RECT 251.100 298.500 266.780 298.560 ;
        RECT 271.210 298.500 286.890 298.560 ;
        RECT 210.970 298.330 226.730 298.500 ;
        RECT 230.990 298.330 246.700 298.500 ;
        RECT 251.100 298.330 266.810 298.500 ;
        RECT 271.210 298.330 286.920 298.500 ;
        RECT 210.970 298.290 226.700 298.330 ;
        RECT 230.990 298.290 246.670 298.330 ;
        RECT 251.100 298.290 266.780 298.330 ;
        RECT 271.210 298.290 286.890 298.330 ;
        RECT 210.970 298.250 212.450 298.290 ;
        RECT 230.990 298.250 232.420 298.290 ;
        RECT 251.100 298.250 252.530 298.290 ;
        RECT 271.210 298.250 272.640 298.290 ;
        RECT 210.970 297.750 211.430 298.250 ;
        RECT 11.800 296.920 102.640 297.070 ;
        RECT 11.800 296.600 104.200 296.920 ;
        RECT 4.540 296.280 104.200 296.600 ;
        RECT 11.800 296.220 104.200 296.280 ;
        RECT 13.050 289.970 13.390 296.220 ;
        RECT 4.780 289.930 13.390 289.970 ;
        RECT 26.390 289.950 26.730 296.220 ;
        RECT 39.760 289.980 40.100 296.220 ;
        RECT 52.990 289.980 53.330 296.220 ;
        RECT 4.610 289.760 13.390 289.930 ;
        RECT 18.120 289.910 26.730 289.950 ;
        RECT 31.490 289.940 40.100 289.980 ;
        RECT 44.720 289.940 53.330 289.980 ;
        RECT 66.260 289.950 66.600 296.220 ;
        RECT 79.530 289.980 79.870 296.220 ;
        RECT 92.660 290.000 93.000 296.220 ;
        RECT 102.150 296.180 104.200 296.220 ;
        RECT 98.060 290.200 102.070 290.230 ;
        RECT 102.390 290.200 102.800 296.180 ;
        RECT 211.020 292.020 211.430 297.750 ;
        RECT 230.990 292.020 231.400 298.250 ;
        RECT 251.100 292.020 251.510 298.250 ;
        RECT 271.210 292.020 271.620 298.250 ;
        RECT 379.090 294.900 379.370 308.900 ;
        RECT 385.720 308.670 385.890 309.060 ;
        RECT 595.315 309.035 595.645 310.140 ;
        RECT 595.825 310.430 596.535 310.475 ;
        RECT 597.000 310.430 597.630 310.540 ;
        RECT 595.825 310.090 597.630 310.430 ;
        RECT 596.270 310.070 597.630 310.090 ;
        RECT 597.000 309.690 597.630 310.070 ;
        RECT 634.090 310.500 635.650 310.540 ;
        RECT 634.090 310.050 634.370 310.500 ;
        RECT 379.040 294.680 379.370 294.900 ;
        RECT 385.660 294.890 385.940 308.670 ;
        RECT 631.570 308.560 632.520 309.450 ;
        RECT 633.870 309.370 634.580 310.050 ;
        RECT 636.125 309.485 636.455 310.560 ;
        RECT 610.250 307.650 610.420 308.070 ;
        RECT 611.040 307.650 611.210 308.070 ;
        RECT 611.830 307.650 612.000 308.070 ;
        RECT 612.620 307.650 612.790 308.070 ;
        RECT 613.410 307.650 613.580 308.070 ;
        RECT 617.840 307.620 618.010 308.040 ;
        RECT 618.630 307.620 618.800 308.040 ;
        RECT 619.420 307.620 619.590 308.040 ;
        RECT 620.210 307.620 620.380 308.040 ;
        RECT 621.000 307.620 621.170 308.040 ;
        RECT 600.800 306.870 600.970 307.290 ;
        RECT 601.590 306.870 601.760 307.290 ;
        RECT 602.380 306.870 602.550 307.290 ;
        RECT 603.170 306.870 603.340 307.290 ;
        RECT 603.960 306.870 604.130 307.290 ;
        RECT 615.360 307.140 615.840 307.560 ;
        RECT 627.580 307.000 627.750 307.420 ;
        RECT 628.370 307.000 628.540 307.420 ;
        RECT 629.160 307.000 629.330 307.420 ;
        RECT 629.950 307.000 630.120 307.420 ;
        RECT 630.740 307.000 630.910 307.420 ;
        RECT 637.330 306.630 637.730 310.560 ;
        RECT 640.315 309.575 640.645 310.690 ;
        RECT 641.800 310.350 642.030 310.690 ;
        RECT 643.525 310.610 644.235 310.690 ;
        RECT 644.415 310.790 644.745 311.235 ;
        RECT 645.310 310.790 645.620 310.810 ;
        RECT 644.415 310.610 645.620 310.790 ;
        RECT 641.730 310.030 642.110 310.350 ;
        RECT 644.415 309.555 644.745 310.610 ;
        RECT 645.310 310.460 645.620 310.610 ;
        RECT 666.600 310.600 666.960 313.080 ;
        RECT 646.040 308.960 646.680 310.320 ;
        RECT 666.600 309.280 666.980 310.600 ;
        RECT 666.230 307.830 667.540 309.280 ;
        RECT 639.690 306.630 640.140 306.730 ;
        RECT 591.850 304.210 592.200 306.370 ;
        RECT 610.250 306.180 610.420 306.600 ;
        RECT 611.040 306.180 611.210 306.600 ;
        RECT 611.830 306.180 612.000 306.600 ;
        RECT 612.620 306.180 612.790 306.600 ;
        RECT 613.410 306.180 613.580 306.600 ;
        RECT 614.080 306.130 614.250 306.550 ;
        RECT 615.660 306.130 615.830 306.550 ;
        RECT 617.240 306.130 617.410 306.550 ;
        RECT 617.840 306.150 618.010 306.570 ;
        RECT 618.630 306.150 618.800 306.570 ;
        RECT 619.420 306.150 619.590 306.570 ;
        RECT 620.210 306.150 620.380 306.570 ;
        RECT 621.000 306.150 621.170 306.570 ;
        RECT 637.330 306.440 640.140 306.630 ;
        RECT 637.330 306.430 637.730 306.440 ;
        RECT 600.800 305.400 600.970 305.820 ;
        RECT 601.590 305.400 601.760 305.820 ;
        RECT 602.380 305.400 602.550 305.820 ;
        RECT 603.170 305.400 603.340 305.820 ;
        RECT 603.960 305.400 604.130 305.820 ;
        RECT 608.370 305.710 609.040 306.020 ;
        RECT 622.960 305.600 623.650 306.150 ;
        RECT 639.690 306.040 640.140 306.440 ;
        RECT 643.750 306.100 644.170 306.780 ;
        RECT 627.580 305.530 627.750 305.950 ;
        RECT 628.370 305.530 628.540 305.950 ;
        RECT 629.160 305.530 629.330 305.950 ;
        RECT 629.950 305.530 630.120 305.950 ;
        RECT 630.740 305.530 630.910 305.950 ;
        RECT 639.430 305.240 639.600 305.660 ;
        RECT 643.480 305.290 643.650 305.710 ;
        RECT 606.500 304.660 606.670 305.080 ;
        RECT 607.290 304.660 607.460 305.080 ;
        RECT 608.080 304.660 608.250 305.080 ;
        RECT 608.870 304.660 609.040 305.080 ;
        RECT 609.660 304.660 609.830 305.080 ;
        RECT 610.250 304.710 610.420 305.130 ;
        RECT 611.040 304.710 611.210 305.130 ;
        RECT 611.830 304.710 612.000 305.130 ;
        RECT 612.620 304.710 612.790 305.130 ;
        RECT 613.410 304.710 613.580 305.130 ;
        RECT 614.080 304.660 614.250 305.080 ;
        RECT 615.660 304.660 615.830 305.080 ;
        RECT 617.240 304.660 617.410 305.080 ;
        RECT 617.840 304.680 618.010 305.100 ;
        RECT 618.630 304.680 618.800 305.100 ;
        RECT 619.420 304.680 619.590 305.100 ;
        RECT 620.210 304.680 620.380 305.100 ;
        RECT 621.000 304.680 621.170 305.100 ;
        RECT 621.590 304.660 621.760 305.080 ;
        RECT 622.380 304.660 622.550 305.080 ;
        RECT 623.170 304.660 623.340 305.080 ;
        RECT 623.960 304.660 624.130 305.080 ;
        RECT 624.750 304.660 624.920 305.080 ;
        RECT 602.070 303.750 602.850 304.190 ;
        RECT 591.850 301.050 592.200 303.210 ;
        RECT 696.730 302.210 697.100 315.840 ;
        RECT 797.880 307.665 799.320 307.835 ;
        RECT 796.590 306.555 796.920 307.485 ;
        RECT 797.880 306.555 798.050 307.665 ;
        RECT 796.590 306.385 798.050 306.555 ;
        RECT 796.590 304.525 796.860 306.385 ;
        RECT 797.040 305.205 797.370 306.180 ;
        RECT 797.720 305.885 798.050 306.385 ;
        RECT 798.230 306.180 798.480 307.485 ;
        RECT 798.720 306.870 798.970 307.485 ;
        RECT 799.150 307.220 799.320 307.665 ;
        RECT 800.010 307.665 801.750 307.835 ;
        RECT 800.010 307.220 800.180 307.665 ;
        RECT 799.150 307.050 800.180 307.220 ;
        RECT 800.360 306.870 800.530 307.485 ;
        RECT 801.060 307.230 801.390 307.485 ;
        RECT 798.720 306.700 800.530 306.870 ;
        RECT 800.710 306.700 800.930 307.030 ;
        RECT 800.360 306.520 800.530 306.700 ;
        RECT 800.360 306.350 800.580 306.520 ;
        RECT 798.230 305.950 798.755 306.180 ;
        RECT 798.230 305.025 798.500 305.950 ;
        RECT 798.170 304.525 798.500 305.025 ;
        RECT 799.895 304.840 800.225 306.135 ;
        RECT 800.410 305.355 800.580 306.350 ;
        RECT 800.760 306.180 800.930 306.700 ;
        RECT 801.110 306.530 801.280 307.230 ;
        RECT 801.580 307.075 801.750 307.665 ;
        RECT 803.060 307.665 804.090 307.835 ;
        RECT 803.060 307.075 803.230 307.665 ;
        RECT 801.580 307.030 803.230 307.075 ;
        RECT 801.460 306.905 803.230 307.030 ;
        RECT 801.460 306.710 801.790 306.905 ;
        RECT 803.410 306.725 803.740 307.485 ;
        RECT 803.920 307.305 804.090 307.665 ;
        RECT 803.920 307.135 805.730 307.305 ;
        RECT 801.970 306.555 803.740 306.725 ;
        RECT 801.970 306.530 802.140 306.555 ;
        RECT 801.110 306.360 802.140 306.530 ;
        RECT 805.050 306.375 805.380 306.955 ;
        RECT 800.760 305.950 801.785 306.180 ;
        RECT 801.455 305.455 801.785 305.950 ;
        RECT 801.970 305.675 802.140 306.360 ;
        RECT 802.320 306.205 805.380 306.375 ;
        RECT 802.320 305.855 802.650 306.205 ;
        RECT 801.970 305.505 804.590 305.675 ;
        RECT 800.410 304.855 800.680 305.355 ;
        RECT 801.970 305.275 802.140 305.505 ;
        RECT 801.130 305.105 802.140 305.275 ;
        RECT 805.120 305.355 805.380 306.205 ;
        RECT 805.560 305.785 805.730 307.135 ;
        RECT 805.910 306.875 806.160 307.785 ;
        RECT 805.910 306.705 806.785 306.875 ;
        RECT 806.105 305.965 806.435 306.465 ;
        RECT 806.615 306.385 806.785 306.705 ;
        RECT 808.320 306.735 808.570 307.205 ;
        RECT 808.320 306.565 809.325 306.735 ;
        RECT 806.615 306.215 808.975 306.385 ;
        RECT 805.560 305.615 806.730 305.785 ;
        RECT 801.130 304.855 801.460 305.105 ;
        RECT 805.120 304.645 805.450 305.355 ;
        RECT 805.910 304.815 806.240 305.355 ;
        RECT 806.445 305.115 806.730 305.615 ;
        RECT 806.910 304.815 807.080 306.215 ;
        RECT 809.155 306.035 809.325 306.565 ;
        RECT 807.285 305.865 809.325 306.035 ;
        RECT 807.285 305.475 807.615 305.865 ;
        RECT 805.910 304.645 807.080 304.815 ;
        RECT 809.100 305.025 809.325 305.865 ;
        RECT 809.825 306.035 810.075 307.035 ;
        RECT 809.825 305.705 811.200 306.035 ;
        RECT 811.380 305.860 811.715 307.765 ;
        RECT 815.640 307.665 817.080 307.835 ;
        RECT 814.350 306.555 814.680 307.485 ;
        RECT 815.640 306.555 815.810 307.665 ;
        RECT 814.350 306.385 815.810 306.555 ;
        RECT 809.825 305.525 810.035 305.705 ;
        RECT 809.705 305.025 810.035 305.525 ;
        RECT 811.380 305.630 811.720 305.860 ;
        RECT 809.100 304.525 809.430 305.025 ;
        RECT 811.380 304.695 811.715 305.630 ;
        RECT 814.350 304.525 814.620 306.385 ;
        RECT 814.840 306.180 815.130 306.200 ;
        RECT 814.800 305.205 815.130 306.180 ;
        RECT 815.480 305.885 815.810 306.385 ;
        RECT 815.990 306.180 816.240 307.485 ;
        RECT 816.480 306.870 816.730 307.485 ;
        RECT 816.910 307.220 817.080 307.665 ;
        RECT 817.770 307.665 819.510 307.835 ;
        RECT 817.770 307.220 817.940 307.665 ;
        RECT 816.910 307.050 817.940 307.220 ;
        RECT 818.120 306.870 818.290 307.485 ;
        RECT 818.820 307.230 819.150 307.485 ;
        RECT 816.480 306.700 818.290 306.870 ;
        RECT 818.470 306.700 818.690 307.030 ;
        RECT 818.120 306.520 818.290 306.700 ;
        RECT 818.120 306.350 818.340 306.520 ;
        RECT 815.990 305.950 816.515 306.180 ;
        RECT 815.990 305.025 816.260 305.950 ;
        RECT 815.930 304.525 816.260 305.025 ;
        RECT 817.655 304.840 817.985 306.135 ;
        RECT 818.170 305.355 818.340 306.350 ;
        RECT 818.520 306.180 818.690 306.700 ;
        RECT 818.870 306.530 819.040 307.230 ;
        RECT 819.340 307.075 819.510 307.665 ;
        RECT 820.820 307.665 821.850 307.835 ;
        RECT 820.820 307.075 820.990 307.665 ;
        RECT 819.340 307.030 820.990 307.075 ;
        RECT 819.220 306.905 820.990 307.030 ;
        RECT 819.220 306.710 819.550 306.905 ;
        RECT 821.170 306.725 821.500 307.485 ;
        RECT 821.680 307.305 821.850 307.665 ;
        RECT 821.680 307.135 823.490 307.305 ;
        RECT 819.730 306.555 821.500 306.725 ;
        RECT 819.730 306.530 819.900 306.555 ;
        RECT 818.870 306.360 819.900 306.530 ;
        RECT 822.810 306.375 823.140 306.955 ;
        RECT 818.520 305.950 819.545 306.180 ;
        RECT 819.215 305.455 819.545 305.950 ;
        RECT 819.730 305.675 819.900 306.360 ;
        RECT 820.080 306.205 823.140 306.375 ;
        RECT 820.080 305.855 820.410 306.205 ;
        RECT 819.730 305.505 822.350 305.675 ;
        RECT 818.170 304.855 818.440 305.355 ;
        RECT 819.730 305.275 819.900 305.505 ;
        RECT 818.890 305.105 819.900 305.275 ;
        RECT 822.880 305.355 823.140 306.205 ;
        RECT 823.320 305.785 823.490 307.135 ;
        RECT 823.670 306.875 823.920 307.785 ;
        RECT 823.670 306.705 824.545 306.875 ;
        RECT 823.865 305.965 824.195 306.465 ;
        RECT 824.375 306.385 824.545 306.705 ;
        RECT 826.080 306.735 826.330 307.205 ;
        RECT 826.080 306.565 827.085 306.735 ;
        RECT 824.375 306.215 826.735 306.385 ;
        RECT 823.320 305.615 824.490 305.785 ;
        RECT 818.890 304.855 819.220 305.105 ;
        RECT 822.880 304.645 823.210 305.355 ;
        RECT 823.670 304.815 824.000 305.355 ;
        RECT 824.205 305.115 824.490 305.615 ;
        RECT 824.670 304.815 824.840 306.215 ;
        RECT 826.915 306.035 827.085 306.565 ;
        RECT 825.045 305.865 827.085 306.035 ;
        RECT 825.045 305.475 825.375 305.865 ;
        RECT 823.670 304.645 824.840 304.815 ;
        RECT 826.860 305.025 827.085 305.865 ;
        RECT 827.585 306.035 827.835 307.035 ;
        RECT 827.585 305.705 828.960 306.035 ;
        RECT 829.140 305.850 829.475 307.765 ;
        RECT 832.740 306.175 833.125 307.755 ;
        RECT 834.140 306.630 834.430 306.970 ;
        RECT 831.905 305.850 832.615 305.935 ;
        RECT 827.585 305.525 827.795 305.705 ;
        RECT 827.465 305.025 827.795 305.525 ;
        RECT 829.140 305.650 832.615 305.850 ;
        RECT 826.860 304.525 827.190 305.025 ;
        RECT 829.140 304.695 829.475 305.650 ;
        RECT 831.905 305.550 832.615 305.650 ;
        RECT 832.795 304.495 833.125 306.175 ;
        RECT 834.260 305.700 834.430 306.630 ;
        RECT 835.550 306.665 835.800 307.815 ;
        RECT 838.130 307.185 838.300 307.815 ;
        RECT 840.320 307.185 840.570 307.815 ;
        RECT 838.130 307.015 840.570 307.185 ;
        RECT 838.130 306.845 838.300 307.015 ;
        RECT 838.480 306.665 840.140 306.835 ;
        RECT 835.550 306.495 838.650 306.665 ;
        RECT 834.180 305.460 834.530 305.700 ;
        RECT 835.550 305.655 835.800 306.495 ;
        RECT 835.980 305.835 836.930 306.115 ;
        RECT 837.465 305.835 838.655 306.210 ;
        RECT 836.760 305.655 836.930 305.835 ;
        RECT 838.835 305.655 839.135 305.895 ;
        RECT 835.550 305.485 836.580 305.655 ;
        RECT 836.760 305.565 839.135 305.655 ;
        RECT 836.760 305.485 839.005 305.565 ;
        RECT 836.330 304.555 836.580 305.485 ;
        RECT 839.385 305.385 839.790 306.485 ;
        RECT 839.970 306.055 840.140 306.665 ;
        RECT 840.320 306.235 840.570 307.015 ;
        RECT 843.650 306.235 844.035 307.815 ;
        RECT 839.970 305.725 840.300 306.055 ;
        RECT 842.815 305.610 843.525 305.995 ;
        RECT 843.705 305.820 844.035 306.235 ;
        RECT 844.600 305.820 845.200 332.510 ;
        RECT 852.620 331.640 852.790 332.060 ;
        RECT 855.200 331.640 855.370 332.060 ;
        RECT 865.750 331.110 866.550 333.680 ;
        RECT 870.930 332.200 871.690 345.690 ;
        RECT 870.740 331.110 871.790 332.200 ;
        RECT 852.620 330.170 852.790 330.590 ;
        RECT 855.200 330.170 855.370 330.590 ;
        RECT 865.520 330.490 866.770 331.110 ;
        RECT 869.930 330.000 870.100 330.420 ;
        RECT 871.220 330.000 871.390 330.420 ;
        RECT 872.510 330.000 872.680 330.420 ;
        RECT 864.740 329.450 864.910 329.870 ;
        RECT 866.030 329.450 866.200 329.870 ;
        RECT 867.320 329.450 867.490 329.870 ;
        RECT 852.620 328.700 852.790 329.120 ;
        RECT 855.200 328.700 855.370 329.120 ;
        RECT 869.930 328.530 870.100 328.950 ;
        RECT 871.220 328.530 871.390 328.950 ;
        RECT 872.510 328.530 872.680 328.950 ;
        RECT 864.740 327.980 864.910 328.400 ;
        RECT 866.030 327.980 866.200 328.400 ;
        RECT 867.320 327.980 867.490 328.400 ;
        RECT 852.620 327.230 852.790 327.650 ;
        RECT 855.200 327.230 855.370 327.650 ;
        RECT 859.460 327.420 859.630 327.840 ;
        RECT 862.040 327.420 862.210 327.840 ;
        RECT 869.930 327.060 870.100 327.480 ;
        RECT 871.220 327.060 871.390 327.480 ;
        RECT 872.510 327.060 872.680 327.480 ;
        RECT 864.740 326.510 864.910 326.930 ;
        RECT 866.030 326.510 866.200 326.930 ;
        RECT 867.320 326.510 867.490 326.930 ;
        RECT 852.620 325.760 852.790 326.180 ;
        RECT 855.200 325.760 855.370 326.180 ;
        RECT 859.460 325.950 859.630 326.370 ;
        RECT 862.040 325.950 862.210 326.370 ;
        RECT 869.930 325.590 870.100 326.010 ;
        RECT 871.220 325.590 871.390 326.010 ;
        RECT 872.510 325.590 872.680 326.010 ;
        RECT 864.740 325.040 864.910 325.460 ;
        RECT 866.030 325.040 866.200 325.460 ;
        RECT 867.320 325.040 867.490 325.460 ;
        RECT 852.620 324.290 852.790 324.710 ;
        RECT 855.200 324.290 855.370 324.710 ;
        RECT 859.460 324.480 859.630 324.900 ;
        RECT 862.040 324.480 862.210 324.900 ;
        RECT 869.930 324.120 870.100 324.540 ;
        RECT 871.220 324.120 871.390 324.540 ;
        RECT 872.510 324.120 872.680 324.540 ;
        RECT 864.740 323.570 864.910 323.990 ;
        RECT 866.030 323.570 866.200 323.990 ;
        RECT 867.320 323.570 867.490 323.990 ;
        RECT 852.620 322.820 852.790 323.240 ;
        RECT 855.200 322.820 855.370 323.240 ;
        RECT 859.460 323.010 859.630 323.430 ;
        RECT 862.040 323.010 862.210 323.430 ;
        RECT 852.620 321.350 852.790 321.770 ;
        RECT 855.200 321.350 855.370 321.770 ;
        RECT 859.460 321.540 859.630 321.960 ;
        RECT 862.040 321.540 862.210 321.960 ;
        RECT 874.010 321.430 875.020 321.930 ;
        RECT 852.620 319.880 852.790 320.300 ;
        RECT 855.200 319.880 855.370 320.300 ;
        RECT 859.460 320.070 859.630 320.490 ;
        RECT 862.040 320.070 862.210 320.490 ;
        RECT 869.970 320.440 870.140 320.860 ;
        RECT 873.220 320.380 873.390 320.800 ;
        RECT 875.800 320.380 875.970 320.800 ;
        RECT 852.620 318.410 852.790 318.830 ;
        RECT 855.200 318.410 855.370 318.830 ;
        RECT 859.460 318.600 859.630 319.020 ;
        RECT 862.040 318.600 862.210 319.020 ;
        RECT 869.970 318.970 870.140 319.390 ;
        RECT 873.220 318.910 873.390 319.330 ;
        RECT 875.800 318.910 875.970 319.330 ;
        RECT 852.620 316.940 852.790 317.360 ;
        RECT 855.200 316.940 855.370 317.360 ;
        RECT 859.460 317.130 859.630 317.550 ;
        RECT 862.040 317.130 862.210 317.550 ;
        RECT 869.970 317.500 870.140 317.920 ;
        RECT 873.220 317.440 873.390 317.860 ;
        RECT 875.800 317.440 875.970 317.860 ;
        RECT 852.620 315.470 852.790 315.890 ;
        RECT 855.200 315.470 855.370 315.890 ;
        RECT 859.460 315.660 859.630 316.080 ;
        RECT 862.040 315.660 862.210 316.080 ;
        RECT 869.970 316.030 870.140 316.450 ;
        RECT 873.220 315.970 873.390 316.390 ;
        RECT 875.800 315.970 875.970 316.390 ;
        RECT 852.620 314.000 852.790 314.420 ;
        RECT 855.200 314.000 855.370 314.420 ;
        RECT 859.460 314.190 859.630 314.610 ;
        RECT 862.040 314.190 862.210 314.610 ;
        RECT 869.970 314.560 870.140 314.980 ;
        RECT 873.220 314.500 873.390 314.920 ;
        RECT 875.800 314.500 875.970 314.920 ;
        RECT 839.270 304.555 839.790 305.385 ;
        RECT 843.705 305.590 845.200 305.820 ;
        RECT 843.705 304.555 844.035 305.590 ;
        RECT 844.600 305.580 845.200 305.590 ;
        RECT 696.400 300.840 697.500 302.210 ;
        RECT 681.460 298.605 682.900 298.775 ;
        RECT 680.170 297.495 680.500 298.425 ;
        RECT 681.460 297.495 681.630 298.605 ;
        RECT 680.170 297.325 681.630 297.495 ;
        RECT 632.300 296.050 633.790 297.100 ;
        RECT 680.170 295.465 680.440 297.325 ;
        RECT 680.620 296.145 680.950 297.120 ;
        RECT 681.300 296.825 681.630 297.325 ;
        RECT 681.810 297.120 682.060 298.425 ;
        RECT 682.300 297.810 682.550 298.425 ;
        RECT 682.730 298.160 682.900 298.605 ;
        RECT 683.590 298.605 685.330 298.775 ;
        RECT 683.590 298.160 683.760 298.605 ;
        RECT 682.730 297.990 683.760 298.160 ;
        RECT 683.940 297.810 684.110 298.425 ;
        RECT 684.640 298.170 684.970 298.425 ;
        RECT 682.300 297.640 684.110 297.810 ;
        RECT 684.290 297.640 684.510 297.970 ;
        RECT 683.940 297.460 684.110 297.640 ;
        RECT 683.940 297.290 684.160 297.460 ;
        RECT 681.810 296.890 682.335 297.120 ;
        RECT 681.810 295.965 682.080 296.890 ;
        RECT 681.750 295.465 682.080 295.965 ;
        RECT 683.475 295.780 683.805 297.075 ;
        RECT 683.990 296.295 684.160 297.290 ;
        RECT 684.340 297.120 684.510 297.640 ;
        RECT 684.690 297.470 684.860 298.170 ;
        RECT 685.160 298.015 685.330 298.605 ;
        RECT 686.640 298.605 687.670 298.775 ;
        RECT 686.640 298.015 686.810 298.605 ;
        RECT 685.160 297.970 686.810 298.015 ;
        RECT 685.040 297.845 686.810 297.970 ;
        RECT 685.040 297.650 685.370 297.845 ;
        RECT 686.990 297.665 687.320 298.425 ;
        RECT 687.500 298.245 687.670 298.605 ;
        RECT 687.500 298.075 689.310 298.245 ;
        RECT 685.550 297.495 687.320 297.665 ;
        RECT 685.550 297.470 685.720 297.495 ;
        RECT 684.690 297.300 685.720 297.470 ;
        RECT 688.630 297.315 688.960 297.895 ;
        RECT 684.340 296.890 685.365 297.120 ;
        RECT 685.035 296.395 685.365 296.890 ;
        RECT 685.550 296.615 685.720 297.300 ;
        RECT 685.900 297.145 688.960 297.315 ;
        RECT 685.900 296.795 686.230 297.145 ;
        RECT 685.550 296.445 688.170 296.615 ;
        RECT 683.990 295.795 684.260 296.295 ;
        RECT 685.550 296.215 685.720 296.445 ;
        RECT 684.710 296.045 685.720 296.215 ;
        RECT 688.700 296.295 688.960 297.145 ;
        RECT 689.140 296.725 689.310 298.075 ;
        RECT 689.490 297.815 689.740 298.725 ;
        RECT 689.490 297.645 690.365 297.815 ;
        RECT 689.685 296.905 690.015 297.405 ;
        RECT 690.195 297.325 690.365 297.645 ;
        RECT 691.900 297.675 692.150 298.145 ;
        RECT 691.900 297.505 692.905 297.675 ;
        RECT 690.195 297.155 692.555 297.325 ;
        RECT 689.140 296.555 690.310 296.725 ;
        RECT 684.710 295.795 685.040 296.045 ;
        RECT 688.700 295.585 689.030 296.295 ;
        RECT 689.490 295.755 689.820 296.295 ;
        RECT 690.025 296.055 690.310 296.555 ;
        RECT 690.490 295.755 690.660 297.155 ;
        RECT 692.735 296.975 692.905 297.505 ;
        RECT 690.865 296.805 692.905 296.975 ;
        RECT 690.865 296.415 691.195 296.805 ;
        RECT 689.490 295.585 690.660 295.755 ;
        RECT 692.680 295.965 692.905 296.805 ;
        RECT 693.405 296.975 693.655 297.975 ;
        RECT 693.405 296.645 694.780 296.975 ;
        RECT 693.405 296.465 693.615 296.645 ;
        RECT 693.285 295.965 693.615 296.465 ;
        RECT 692.680 295.465 693.010 295.965 ;
        RECT 694.960 295.635 695.295 298.705 ;
        RECT 698.950 298.565 700.390 298.735 ;
        RECT 697.660 297.455 697.990 298.385 ;
        RECT 698.950 297.455 699.120 298.565 ;
        RECT 697.660 297.285 699.120 297.455 ;
        RECT 697.660 295.425 697.930 297.285 ;
        RECT 698.110 296.580 698.440 297.080 ;
        RECT 698.790 296.785 699.120 297.285 ;
        RECT 699.300 297.080 699.550 298.385 ;
        RECT 699.790 297.770 700.040 298.385 ;
        RECT 700.220 298.120 700.390 298.565 ;
        RECT 701.080 298.565 702.820 298.735 ;
        RECT 701.080 298.120 701.250 298.565 ;
        RECT 700.220 297.950 701.250 298.120 ;
        RECT 701.430 297.770 701.600 298.385 ;
        RECT 702.130 298.130 702.460 298.385 ;
        RECT 699.790 297.600 701.600 297.770 ;
        RECT 701.780 297.600 702.000 297.930 ;
        RECT 701.430 297.420 701.600 297.600 ;
        RECT 701.430 297.250 701.650 297.420 ;
        RECT 699.300 296.850 699.825 297.080 ;
        RECT 698.110 296.300 698.480 296.580 ;
        RECT 698.110 296.105 698.440 296.300 ;
        RECT 699.300 295.925 699.570 296.850 ;
        RECT 699.240 295.425 699.570 295.925 ;
        RECT 700.965 295.740 701.295 297.035 ;
        RECT 701.480 296.255 701.650 297.250 ;
        RECT 701.830 297.080 702.000 297.600 ;
        RECT 702.180 297.430 702.350 298.130 ;
        RECT 702.650 297.975 702.820 298.565 ;
        RECT 704.130 298.565 705.160 298.735 ;
        RECT 704.130 297.975 704.300 298.565 ;
        RECT 702.650 297.930 704.300 297.975 ;
        RECT 702.530 297.805 704.300 297.930 ;
        RECT 702.530 297.610 702.860 297.805 ;
        RECT 704.480 297.625 704.810 298.385 ;
        RECT 704.990 298.205 705.160 298.565 ;
        RECT 704.990 298.035 706.800 298.205 ;
        RECT 703.040 297.455 704.810 297.625 ;
        RECT 703.040 297.430 703.210 297.455 ;
        RECT 702.180 297.260 703.210 297.430 ;
        RECT 706.120 297.275 706.450 297.855 ;
        RECT 701.830 296.850 702.855 297.080 ;
        RECT 702.525 296.355 702.855 296.850 ;
        RECT 703.040 296.575 703.210 297.260 ;
        RECT 703.390 297.105 706.450 297.275 ;
        RECT 703.390 296.755 703.720 297.105 ;
        RECT 703.040 296.405 705.660 296.575 ;
        RECT 701.480 295.755 701.750 296.255 ;
        RECT 703.040 296.175 703.210 296.405 ;
        RECT 702.200 296.005 703.210 296.175 ;
        RECT 706.190 296.255 706.450 297.105 ;
        RECT 706.630 296.685 706.800 298.035 ;
        RECT 706.980 297.775 707.230 298.685 ;
        RECT 706.980 297.605 707.855 297.775 ;
        RECT 707.175 296.865 707.505 297.365 ;
        RECT 707.685 297.285 707.855 297.605 ;
        RECT 709.390 297.635 709.640 298.105 ;
        RECT 709.390 297.465 710.395 297.635 ;
        RECT 707.685 297.115 710.045 297.285 ;
        RECT 706.630 296.515 707.800 296.685 ;
        RECT 702.200 295.755 702.530 296.005 ;
        RECT 706.190 295.545 706.520 296.255 ;
        RECT 706.980 295.715 707.310 296.255 ;
        RECT 707.515 296.015 707.800 296.515 ;
        RECT 707.980 295.715 708.150 297.115 ;
        RECT 710.225 296.935 710.395 297.465 ;
        RECT 708.355 296.765 710.395 296.935 ;
        RECT 708.355 296.375 708.685 296.765 ;
        RECT 706.980 295.545 708.150 295.715 ;
        RECT 710.170 295.925 710.395 296.765 ;
        RECT 710.895 296.935 711.145 297.935 ;
        RECT 712.450 297.790 712.785 298.665 ;
        RECT 716.560 298.625 718.000 298.795 ;
        RECT 712.450 297.020 712.800 297.790 ;
        RECT 715.270 297.515 715.600 298.445 ;
        RECT 716.560 297.515 716.730 298.625 ;
        RECT 715.270 297.345 716.730 297.515 ;
        RECT 710.895 296.605 712.270 296.935 ;
        RECT 710.895 296.425 711.105 296.605 ;
        RECT 710.775 295.925 711.105 296.425 ;
        RECT 710.170 295.425 710.500 295.925 ;
        RECT 712.450 295.595 712.785 297.020 ;
        RECT 715.270 295.485 715.540 297.345 ;
        RECT 715.720 296.165 716.050 297.140 ;
        RECT 716.400 296.845 716.730 297.345 ;
        RECT 716.910 297.140 717.160 298.445 ;
        RECT 717.400 297.830 717.650 298.445 ;
        RECT 717.830 298.180 718.000 298.625 ;
        RECT 718.690 298.625 720.430 298.795 ;
        RECT 718.690 298.180 718.860 298.625 ;
        RECT 717.830 298.010 718.860 298.180 ;
        RECT 719.040 297.830 719.210 298.445 ;
        RECT 719.740 298.190 720.070 298.445 ;
        RECT 717.400 297.660 719.210 297.830 ;
        RECT 719.390 297.660 719.610 297.990 ;
        RECT 719.040 297.480 719.210 297.660 ;
        RECT 719.040 297.310 719.260 297.480 ;
        RECT 716.910 296.910 717.435 297.140 ;
        RECT 716.910 295.985 717.180 296.910 ;
        RECT 716.850 295.485 717.180 295.985 ;
        RECT 719.090 296.315 719.260 297.310 ;
        RECT 719.440 297.140 719.610 297.660 ;
        RECT 719.790 297.490 719.960 298.190 ;
        RECT 720.260 298.035 720.430 298.625 ;
        RECT 721.740 298.625 722.770 298.795 ;
        RECT 721.740 298.035 721.910 298.625 ;
        RECT 720.260 297.990 721.910 298.035 ;
        RECT 720.140 297.865 721.910 297.990 ;
        RECT 720.140 297.670 720.470 297.865 ;
        RECT 722.090 297.685 722.420 298.445 ;
        RECT 722.600 298.265 722.770 298.625 ;
        RECT 722.600 298.095 724.410 298.265 ;
        RECT 720.650 297.515 722.420 297.685 ;
        RECT 720.650 297.490 720.820 297.515 ;
        RECT 719.790 297.320 720.820 297.490 ;
        RECT 723.730 297.335 724.060 297.915 ;
        RECT 719.440 296.910 720.465 297.140 ;
        RECT 720.135 296.415 720.465 296.910 ;
        RECT 720.650 296.635 720.820 297.320 ;
        RECT 721.000 297.165 724.060 297.335 ;
        RECT 721.000 296.815 721.330 297.165 ;
        RECT 720.650 296.465 723.270 296.635 ;
        RECT 719.090 295.815 719.360 296.315 ;
        RECT 720.650 296.235 720.820 296.465 ;
        RECT 719.810 296.065 720.820 296.235 ;
        RECT 723.800 296.315 724.060 297.165 ;
        RECT 724.240 296.745 724.410 298.095 ;
        RECT 724.590 297.835 724.840 298.745 ;
        RECT 724.590 297.665 725.465 297.835 ;
        RECT 724.785 296.925 725.115 297.425 ;
        RECT 725.295 297.345 725.465 297.665 ;
        RECT 727.000 297.695 727.250 298.165 ;
        RECT 727.000 297.525 728.005 297.695 ;
        RECT 725.295 297.175 727.655 297.345 ;
        RECT 724.240 296.575 725.410 296.745 ;
        RECT 719.810 295.815 720.140 296.065 ;
        RECT 723.800 295.605 724.130 296.315 ;
        RECT 724.590 295.775 724.920 296.315 ;
        RECT 725.125 296.075 725.410 296.575 ;
        RECT 725.590 295.775 725.760 297.175 ;
        RECT 727.835 296.995 728.005 297.525 ;
        RECT 725.965 296.825 728.005 296.995 ;
        RECT 725.965 296.435 726.295 296.825 ;
        RECT 724.590 295.605 725.760 295.775 ;
        RECT 727.780 295.985 728.005 296.825 ;
        RECT 728.505 296.995 728.755 297.995 ;
        RECT 728.505 296.665 729.880 296.995 ;
        RECT 728.505 296.485 728.715 296.665 ;
        RECT 728.385 295.985 728.715 296.485 ;
        RECT 727.780 295.485 728.110 295.985 ;
        RECT 730.060 295.655 730.395 298.725 ;
        RECT 734.260 298.575 735.700 298.745 ;
        RECT 732.970 297.465 733.300 298.395 ;
        RECT 734.260 297.465 734.430 298.575 ;
        RECT 732.970 297.295 734.430 297.465 ;
        RECT 732.970 295.435 733.240 297.295 ;
        RECT 733.420 296.600 733.750 297.090 ;
        RECT 734.100 296.795 734.430 297.295 ;
        RECT 734.610 297.090 734.860 298.395 ;
        RECT 735.100 297.780 735.350 298.395 ;
        RECT 735.530 298.130 735.700 298.575 ;
        RECT 736.390 298.575 738.130 298.745 ;
        RECT 736.390 298.130 736.560 298.575 ;
        RECT 735.530 297.960 736.560 298.130 ;
        RECT 736.740 297.780 736.910 298.395 ;
        RECT 737.440 298.140 737.770 298.395 ;
        RECT 735.100 297.610 736.910 297.780 ;
        RECT 737.090 297.610 737.310 297.940 ;
        RECT 736.740 297.430 736.910 297.610 ;
        RECT 736.740 297.260 736.960 297.430 ;
        RECT 734.610 296.860 735.135 297.090 ;
        RECT 733.420 296.320 733.770 296.600 ;
        RECT 733.420 296.115 733.750 296.320 ;
        RECT 734.610 295.935 734.880 296.860 ;
        RECT 734.550 295.435 734.880 295.935 ;
        RECT 736.790 296.265 736.960 297.260 ;
        RECT 737.140 297.090 737.310 297.610 ;
        RECT 737.490 297.440 737.660 298.140 ;
        RECT 737.960 297.985 738.130 298.575 ;
        RECT 739.440 298.575 740.470 298.745 ;
        RECT 739.440 297.985 739.610 298.575 ;
        RECT 737.960 297.940 739.610 297.985 ;
        RECT 737.840 297.815 739.610 297.940 ;
        RECT 737.840 297.620 738.170 297.815 ;
        RECT 739.790 297.635 740.120 298.395 ;
        RECT 740.300 298.215 740.470 298.575 ;
        RECT 740.300 298.045 742.110 298.215 ;
        RECT 738.350 297.465 740.120 297.635 ;
        RECT 738.350 297.440 738.520 297.465 ;
        RECT 737.490 297.270 738.520 297.440 ;
        RECT 741.430 297.285 741.760 297.865 ;
        RECT 737.140 296.860 738.165 297.090 ;
        RECT 737.835 296.365 738.165 296.860 ;
        RECT 738.350 296.585 738.520 297.270 ;
        RECT 738.700 297.115 741.760 297.285 ;
        RECT 738.700 296.765 739.030 297.115 ;
        RECT 738.350 296.415 740.970 296.585 ;
        RECT 736.790 295.765 737.060 296.265 ;
        RECT 738.350 296.185 738.520 296.415 ;
        RECT 737.510 296.015 738.520 296.185 ;
        RECT 741.500 296.265 741.760 297.115 ;
        RECT 741.940 296.695 742.110 298.045 ;
        RECT 742.290 297.785 742.540 298.695 ;
        RECT 742.290 297.615 743.165 297.785 ;
        RECT 742.485 296.875 742.815 297.375 ;
        RECT 742.995 297.295 743.165 297.615 ;
        RECT 744.700 297.645 744.950 298.115 ;
        RECT 744.700 297.475 745.705 297.645 ;
        RECT 742.995 297.125 745.355 297.295 ;
        RECT 741.940 296.525 743.110 296.695 ;
        RECT 737.510 295.765 737.840 296.015 ;
        RECT 741.500 295.555 741.830 296.265 ;
        RECT 742.290 295.725 742.620 296.265 ;
        RECT 742.825 296.025 743.110 296.525 ;
        RECT 743.290 295.725 743.460 297.125 ;
        RECT 745.535 296.945 745.705 297.475 ;
        RECT 743.665 296.775 745.705 296.945 ;
        RECT 743.665 296.385 743.995 296.775 ;
        RECT 742.290 295.555 743.460 295.725 ;
        RECT 745.480 295.935 745.705 296.775 ;
        RECT 746.205 296.945 746.455 297.945 ;
        RECT 746.205 296.615 747.580 296.945 ;
        RECT 746.205 296.435 746.415 296.615 ;
        RECT 746.085 295.935 746.415 296.435 ;
        RECT 745.480 295.435 745.810 295.935 ;
        RECT 747.760 295.605 748.095 298.675 ;
        RECT 752.000 298.565 753.440 298.735 ;
        RECT 750.710 297.455 751.040 298.385 ;
        RECT 752.000 297.455 752.170 298.565 ;
        RECT 750.710 297.285 752.170 297.455 ;
        RECT 750.710 295.425 750.980 297.285 ;
        RECT 751.160 296.580 751.490 297.080 ;
        RECT 751.840 296.785 752.170 297.285 ;
        RECT 752.350 297.080 752.600 298.385 ;
        RECT 752.840 297.770 753.090 298.385 ;
        RECT 753.270 298.120 753.440 298.565 ;
        RECT 754.130 298.565 755.870 298.735 ;
        RECT 754.130 298.120 754.300 298.565 ;
        RECT 753.270 297.950 754.300 298.120 ;
        RECT 754.480 297.770 754.650 298.385 ;
        RECT 755.180 298.130 755.510 298.385 ;
        RECT 752.840 297.600 754.650 297.770 ;
        RECT 754.830 297.600 755.050 297.930 ;
        RECT 754.480 297.420 754.650 297.600 ;
        RECT 754.480 297.250 754.700 297.420 ;
        RECT 752.350 296.850 752.875 297.080 ;
        RECT 751.160 296.300 751.500 296.580 ;
        RECT 751.160 296.105 751.490 296.300 ;
        RECT 752.350 295.925 752.620 296.850 ;
        RECT 752.290 295.425 752.620 295.925 ;
        RECT 754.530 296.255 754.700 297.250 ;
        RECT 754.880 297.080 755.050 297.600 ;
        RECT 755.230 297.430 755.400 298.130 ;
        RECT 755.700 297.975 755.870 298.565 ;
        RECT 757.180 298.565 758.210 298.735 ;
        RECT 757.180 297.975 757.350 298.565 ;
        RECT 755.700 297.930 757.350 297.975 ;
        RECT 755.580 297.805 757.350 297.930 ;
        RECT 755.580 297.610 755.910 297.805 ;
        RECT 757.530 297.625 757.860 298.385 ;
        RECT 758.040 298.205 758.210 298.565 ;
        RECT 758.040 298.035 759.850 298.205 ;
        RECT 756.090 297.455 757.860 297.625 ;
        RECT 756.090 297.430 756.260 297.455 ;
        RECT 755.230 297.260 756.260 297.430 ;
        RECT 759.170 297.275 759.500 297.855 ;
        RECT 754.880 296.850 755.905 297.080 ;
        RECT 755.575 296.355 755.905 296.850 ;
        RECT 756.090 296.575 756.260 297.260 ;
        RECT 756.440 297.105 759.500 297.275 ;
        RECT 756.440 296.755 756.770 297.105 ;
        RECT 756.090 296.405 758.710 296.575 ;
        RECT 754.530 295.755 754.800 296.255 ;
        RECT 756.090 296.175 756.260 296.405 ;
        RECT 755.250 296.005 756.260 296.175 ;
        RECT 759.240 296.255 759.500 297.105 ;
        RECT 759.680 296.685 759.850 298.035 ;
        RECT 760.030 297.775 760.280 298.685 ;
        RECT 760.030 297.605 760.905 297.775 ;
        RECT 760.225 296.865 760.555 297.365 ;
        RECT 760.735 297.285 760.905 297.605 ;
        RECT 762.440 297.635 762.690 298.105 ;
        RECT 762.440 297.465 763.445 297.635 ;
        RECT 760.735 297.115 763.095 297.285 ;
        RECT 759.680 296.515 760.850 296.685 ;
        RECT 755.250 295.755 755.580 296.005 ;
        RECT 759.240 295.545 759.570 296.255 ;
        RECT 760.030 295.715 760.360 296.255 ;
        RECT 760.565 296.015 760.850 296.515 ;
        RECT 761.030 295.715 761.200 297.115 ;
        RECT 763.275 296.935 763.445 297.465 ;
        RECT 761.405 296.765 763.445 296.935 ;
        RECT 761.405 296.375 761.735 296.765 ;
        RECT 760.030 295.545 761.200 295.715 ;
        RECT 763.220 295.925 763.445 296.765 ;
        RECT 763.945 296.935 764.195 297.935 ;
        RECT 763.945 296.605 765.320 296.935 ;
        RECT 763.945 296.425 764.155 296.605 ;
        RECT 763.825 295.925 764.155 296.425 ;
        RECT 763.220 295.425 763.550 295.925 ;
        RECT 765.500 295.595 765.835 298.665 ;
        RECT 857.000 296.365 857.170 296.965 ;
        RECT 856.515 296.195 858.575 296.365 ;
        RECT 379.040 293.690 379.340 294.680 ;
        RECT 385.660 294.450 385.980 294.890 ;
        RECT 603.220 294.700 603.390 295.120 ;
        RECT 604.800 294.700 604.970 295.120 ;
        RECT 607.740 294.710 607.910 295.130 ;
        RECT 609.320 294.710 609.490 295.130 ;
        RECT 612.260 294.710 612.430 295.130 ;
        RECT 613.840 294.710 614.010 295.130 ;
        RECT 616.690 294.690 616.860 295.110 ;
        RECT 618.270 294.690 618.440 295.110 ;
        RECT 621.070 294.700 621.240 295.120 ;
        RECT 622.650 294.700 622.820 295.120 ;
        RECT 625.390 294.690 625.560 295.110 ;
        RECT 626.970 294.690 627.140 295.110 ;
        RECT 385.680 293.710 385.980 294.450 ;
        RECT 840.590 294.385 840.760 294.985 ;
        RECT 840.105 294.215 842.165 294.385 ;
        RECT 836.030 293.820 836.420 293.920 ;
        RECT 839.515 293.820 839.925 294.155 ;
        RECT 385.680 293.690 386.470 293.710 ;
        RECT 379.040 293.380 386.470 293.690 ;
        RECT 379.040 293.350 379.340 293.380 ;
        RECT 385.680 293.340 385.980 293.380 ;
        RECT 603.220 293.230 603.390 293.650 ;
        RECT 604.800 293.230 604.970 293.650 ;
        RECT 607.740 293.240 607.910 293.660 ;
        RECT 609.320 293.240 609.490 293.660 ;
        RECT 612.260 293.240 612.430 293.660 ;
        RECT 613.840 293.240 614.010 293.660 ;
        RECT 616.690 293.220 616.860 293.640 ;
        RECT 618.270 293.220 618.440 293.640 ;
        RECT 621.070 293.230 621.240 293.650 ;
        RECT 622.650 293.230 622.820 293.650 ;
        RECT 625.390 293.220 625.560 293.640 ;
        RECT 626.970 293.220 627.140 293.640 ;
        RECT 211.000 291.980 212.600 292.020 ;
        RECT 230.970 291.980 232.570 292.020 ;
        RECT 251.080 291.980 252.680 292.020 ;
        RECT 271.190 291.980 272.790 292.020 ;
        RECT 211.000 291.710 226.740 291.980 ;
        RECT 230.970 291.710 246.710 291.980 ;
        RECT 251.080 291.710 266.820 291.980 ;
        RECT 271.190 291.710 286.930 291.980 ;
        RECT 211.000 291.640 212.600 291.710 ;
        RECT 230.970 291.640 232.570 291.710 ;
        RECT 251.080 291.640 252.680 291.710 ;
        RECT 271.190 291.640 272.790 291.710 ;
        RECT 98.060 290.180 102.800 290.200 ;
        RECT 97.640 290.010 102.800 290.180 ;
        RECT 4.780 289.710 13.390 289.760 ;
        RECT 17.950 289.740 26.730 289.910 ;
        RECT 31.320 289.770 40.100 289.940 ;
        RECT 44.550 289.770 53.330 289.940 ;
        RECT 57.990 289.910 66.600 289.950 ;
        RECT 71.260 289.940 79.870 289.980 ;
        RECT 84.390 289.960 93.000 290.000 ;
        RECT 11.950 289.700 13.390 289.710 ;
        RECT 13.050 283.410 13.390 289.700 ;
        RECT 18.120 289.690 26.730 289.740 ;
        RECT 31.490 289.720 40.100 289.770 ;
        RECT 44.720 289.720 53.330 289.770 ;
        RECT 57.820 289.740 66.600 289.910 ;
        RECT 71.090 289.770 79.870 289.940 ;
        RECT 84.220 289.790 93.000 289.960 ;
        RECT 98.060 289.940 102.800 290.010 ;
        RECT 101.520 289.850 102.800 289.940 ;
        RECT 38.660 289.710 40.100 289.720 ;
        RECT 51.890 289.710 53.330 289.720 ;
        RECT 25.290 289.680 26.730 289.690 ;
        RECT 12.010 283.400 13.390 283.410 ;
        RECT 4.850 283.350 13.390 283.400 ;
        RECT 26.390 283.390 26.730 289.680 ;
        RECT 39.760 283.420 40.100 289.710 ;
        RECT 52.990 283.420 53.330 289.710 ;
        RECT 57.990 289.690 66.600 289.740 ;
        RECT 71.260 289.720 79.870 289.770 ;
        RECT 84.390 289.740 93.000 289.790 ;
        RECT 91.560 289.730 93.000 289.740 ;
        RECT 78.430 289.710 79.870 289.720 ;
        RECT 65.160 289.680 66.600 289.690 ;
        RECT 38.720 283.410 40.100 283.420 ;
        RECT 51.950 283.410 53.330 283.420 ;
        RECT 25.350 283.380 26.730 283.390 ;
        RECT 4.610 283.180 13.390 283.350 ;
        RECT 18.190 283.330 26.730 283.380 ;
        RECT 31.560 283.360 40.100 283.410 ;
        RECT 44.790 283.360 53.330 283.410 ;
        RECT 66.260 283.390 66.600 289.680 ;
        RECT 79.530 283.420 79.870 289.710 ;
        RECT 92.660 283.440 93.000 289.730 ;
        RECT 98.120 283.610 102.130 283.630 ;
        RECT 102.390 283.610 102.800 289.850 ;
        RECT 211.020 285.490 211.430 291.640 ;
        RECT 230.990 285.490 231.400 291.640 ;
        RECT 251.100 285.490 251.510 291.640 ;
        RECT 271.210 285.490 271.620 291.640 ;
        RECT 595.265 291.535 595.650 293.115 ;
        RECT 613.310 292.280 613.780 292.660 ;
        RECT 616.150 292.240 616.580 292.560 ;
        RECT 620.560 292.380 620.970 292.810 ;
        RECT 636.020 291.985 636.405 293.565 ;
        RECT 640.210 292.075 640.595 293.655 ;
        RECT 635.185 291.730 635.895 291.745 ;
        RECT 594.270 291.200 594.950 291.290 ;
        RECT 595.265 291.200 595.595 291.535 ;
        RECT 634.040 291.360 635.895 291.730 ;
        RECT 636.075 291.660 636.405 291.985 ;
        RECT 639.200 291.835 639.570 291.860 ;
        RECT 636.830 291.660 637.670 291.670 ;
        RECT 636.075 291.620 637.670 291.660 ;
        RECT 636.075 291.380 637.680 291.620 ;
        RECT 639.200 291.450 640.085 291.835 ;
        RECT 640.265 291.720 640.595 292.075 ;
        RECT 644.310 292.055 644.695 293.635 ;
        RECT 836.030 293.530 839.925 293.820 ;
        RECT 836.030 293.180 836.420 293.530 ;
        RECT 839.515 293.485 839.925 293.530 ;
        RECT 840.105 293.305 840.275 294.215 ;
        RECT 841.835 294.035 842.165 294.215 ;
        RECT 839.520 293.135 840.275 293.305 ;
        RECT 643.475 291.720 644.185 291.815 ;
        RECT 640.265 291.510 644.185 291.720 ;
        RECT 639.200 291.410 639.570 291.450 ;
        RECT 594.270 290.960 595.595 291.200 ;
        RECT 594.270 290.890 594.950 290.960 ;
        RECT 379.140 290.020 379.310 290.180 ;
        RECT 285.950 285.560 290.460 285.620 ;
        RECT 294.340 285.560 295.920 286.440 ;
        RECT 211.000 285.430 212.500 285.490 ;
        RECT 230.970 285.430 232.470 285.490 ;
        RECT 251.080 285.430 252.580 285.490 ;
        RECT 271.190 285.430 272.690 285.490 ;
        RECT 285.950 285.430 295.920 285.560 ;
        RECT 211.000 285.170 295.920 285.430 ;
        RECT 211.000 285.120 226.710 285.170 ;
        RECT 230.970 285.120 246.680 285.170 ;
        RECT 251.080 285.120 266.790 285.170 ;
        RECT 271.190 285.120 295.920 285.170 ;
        RECT 211.000 285.110 212.410 285.120 ;
        RECT 230.970 285.110 232.380 285.120 ;
        RECT 251.080 285.110 252.490 285.120 ;
        RECT 271.190 285.110 272.600 285.120 ;
        RECT 211.020 285.100 211.430 285.110 ;
        RECT 230.990 285.100 231.400 285.110 ;
        RECT 251.100 285.100 251.510 285.110 ;
        RECT 271.210 285.100 271.620 285.110 ;
        RECT 285.950 284.610 295.920 285.120 ;
        RECT 285.950 284.480 290.460 284.610 ;
        RECT 294.340 284.200 295.920 284.610 ;
        RECT 98.120 283.600 102.890 283.610 ;
        RECT 91.620 283.430 93.000 283.440 ;
        RECT 97.640 283.430 102.890 283.600 ;
        RECT 78.490 283.410 79.870 283.420 ;
        RECT 65.220 283.380 66.600 283.390 ;
        RECT 4.850 283.140 13.390 283.180 ;
        RECT 17.950 283.160 26.730 283.330 ;
        RECT 31.320 283.190 40.100 283.360 ;
        RECT 44.550 283.190 53.330 283.360 ;
        RECT 58.060 283.330 66.600 283.380 ;
        RECT 71.330 283.360 79.870 283.410 ;
        RECT 84.460 283.380 93.000 283.430 ;
        RECT 13.050 276.820 13.390 283.140 ;
        RECT 18.190 283.120 26.730 283.160 ;
        RECT 31.560 283.150 40.100 283.190 ;
        RECT 44.790 283.150 53.330 283.190 ;
        RECT 57.820 283.160 66.600 283.330 ;
        RECT 71.090 283.190 79.870 283.360 ;
        RECT 84.220 283.210 93.000 283.380 ;
        RECT 98.120 283.340 102.890 283.430 ;
        RECT 101.670 283.260 102.890 283.340 ;
        RECT 11.960 276.810 13.390 276.820 ;
        RECT 4.970 276.770 13.390 276.810 ;
        RECT 26.390 276.800 26.730 283.120 ;
        RECT 39.760 276.830 40.100 283.150 ;
        RECT 52.990 276.830 53.330 283.150 ;
        RECT 58.060 283.120 66.600 283.160 ;
        RECT 71.330 283.150 79.870 283.190 ;
        RECT 84.460 283.170 93.000 283.210 ;
        RECT 38.670 276.820 40.100 276.830 ;
        RECT 51.900 276.820 53.330 276.830 ;
        RECT 25.300 276.790 26.730 276.800 ;
        RECT 4.610 276.600 13.390 276.770 ;
        RECT 18.310 276.750 26.730 276.790 ;
        RECT 31.680 276.780 40.100 276.820 ;
        RECT 44.910 276.780 53.330 276.820 ;
        RECT 66.260 276.800 66.600 283.120 ;
        RECT 79.530 276.830 79.870 283.150 ;
        RECT 92.660 276.850 93.000 283.170 ;
        RECT 102.390 278.070 102.800 283.260 ;
        RECT 102.320 277.980 118.870 278.070 ;
        RECT 150.770 277.990 151.070 278.260 ;
        RECT 150.140 277.980 151.070 277.990 ;
        RECT 102.320 277.710 151.070 277.980 ;
        RECT 102.320 277.670 150.230 277.710 ;
        RECT 102.320 277.660 118.870 277.670 ;
        RECT 102.390 277.090 102.800 277.660 ;
        RECT 101.580 277.030 102.800 277.090 ;
        RECT 98.040 277.020 102.800 277.030 ;
        RECT 97.640 276.850 102.800 277.020 ;
        RECT 91.570 276.840 93.000 276.850 ;
        RECT 78.440 276.820 79.870 276.830 ;
        RECT 65.170 276.790 66.600 276.800 ;
        RECT 4.970 276.550 13.390 276.600 ;
        RECT 17.950 276.580 26.730 276.750 ;
        RECT 31.320 276.610 40.100 276.780 ;
        RECT 44.550 276.610 53.330 276.780 ;
        RECT 58.180 276.750 66.600 276.790 ;
        RECT 71.450 276.780 79.870 276.820 ;
        RECT 84.580 276.800 93.000 276.840 ;
        RECT 13.050 273.390 13.390 276.550 ;
        RECT 18.310 276.530 26.730 276.580 ;
        RECT 31.680 276.560 40.100 276.610 ;
        RECT 44.910 276.560 53.330 276.610 ;
        RECT 57.820 276.580 66.600 276.750 ;
        RECT 71.090 276.610 79.870 276.780 ;
        RECT 84.220 276.630 93.000 276.800 ;
        RECT 98.040 276.740 102.800 276.850 ;
        RECT 13.000 273.180 13.390 273.390 ;
        RECT 26.390 273.370 26.730 276.530 ;
        RECT 39.760 273.400 40.100 276.560 ;
        RECT 52.990 273.400 53.330 276.560 ;
        RECT 58.180 276.530 66.600 276.580 ;
        RECT 71.450 276.560 79.870 276.610 ;
        RECT 84.580 276.580 93.000 276.630 ;
        RECT 13.000 270.260 13.370 273.180 ;
        RECT 26.340 273.160 26.730 273.370 ;
        RECT 39.710 273.190 40.100 273.400 ;
        RECT 52.940 273.190 53.330 273.400 ;
        RECT 66.260 273.370 66.600 276.530 ;
        RECT 79.530 273.400 79.870 276.560 ;
        RECT 92.660 273.420 93.000 276.580 ;
        RECT 12.280 270.230 13.390 270.260 ;
        RECT 26.340 270.240 26.710 273.160 ;
        RECT 39.710 270.270 40.080 273.190 ;
        RECT 52.940 270.270 53.310 273.190 ;
        RECT 66.210 273.160 66.600 273.370 ;
        RECT 79.480 273.190 79.870 273.400 ;
        RECT 92.610 273.210 93.000 273.420 ;
        RECT 38.990 270.240 40.100 270.270 ;
        RECT 52.220 270.240 53.330 270.270 ;
        RECT 66.210 270.240 66.580 273.160 ;
        RECT 79.480 270.270 79.850 273.190 ;
        RECT 92.610 270.290 92.980 273.210 ;
        RECT 102.390 270.560 102.800 276.740 ;
        RECT 150.780 271.450 151.060 277.710 ;
        RECT 150.000 271.430 151.060 271.450 ;
        RECT 118.560 271.370 151.060 271.430 ;
        RECT 118.120 271.200 151.060 271.370 ;
        RECT 118.560 271.150 151.060 271.200 ;
        RECT 118.560 271.140 151.040 271.150 ;
        RECT 118.560 271.120 150.130 271.140 ;
        RECT 101.580 270.500 102.800 270.560 ;
        RECT 97.960 270.440 102.800 270.500 ;
        RECT 78.760 270.240 79.870 270.270 ;
        RECT 91.890 270.260 93.000 270.290 ;
        RECT 97.640 270.270 102.800 270.440 ;
        RECT 5.150 270.190 13.390 270.230 ;
        RECT 25.620 270.210 26.730 270.240 ;
        RECT 4.610 270.020 13.390 270.190 ;
        RECT 18.490 270.170 26.730 270.210 ;
        RECT 31.860 270.200 40.100 270.240 ;
        RECT 45.090 270.200 53.330 270.240 ;
        RECT 65.490 270.210 66.600 270.240 ;
        RECT 5.150 269.970 13.390 270.020 ;
        RECT 17.950 270.000 26.730 270.170 ;
        RECT 31.320 270.030 40.100 270.200 ;
        RECT 44.550 270.030 53.330 270.200 ;
        RECT 58.360 270.170 66.600 270.210 ;
        RECT 71.630 270.200 79.870 270.240 ;
        RECT 84.760 270.220 93.000 270.260 ;
        RECT 12.280 269.910 13.390 269.970 ;
        RECT 18.490 269.950 26.730 270.000 ;
        RECT 31.860 269.980 40.100 270.030 ;
        RECT 45.090 269.980 53.330 270.030 ;
        RECT 57.820 270.000 66.600 270.170 ;
        RECT 71.090 270.030 79.870 270.200 ;
        RECT 84.220 270.050 93.000 270.220 ;
        RECT 97.960 270.210 102.800 270.270 ;
        RECT 102.390 270.180 102.800 270.210 ;
        RECT 25.620 269.890 26.730 269.950 ;
        RECT 38.990 269.920 40.100 269.980 ;
        RECT 52.220 269.920 53.330 269.980 ;
        RECT 58.360 269.950 66.600 270.000 ;
        RECT 71.630 269.980 79.870 270.030 ;
        RECT 84.760 270.000 93.000 270.050 ;
        RECT 65.490 269.890 66.600 269.950 ;
        RECT 78.760 269.920 79.870 269.980 ;
        RECT 91.890 269.940 93.000 270.000 ;
        RECT 294.690 232.520 295.590 284.200 ;
        RECT 379.090 276.020 379.370 290.020 ;
        RECT 385.720 289.790 385.890 290.180 ;
        RECT 595.265 289.855 595.595 290.960 ;
        RECT 595.775 291.250 596.485 291.295 ;
        RECT 596.950 291.250 597.580 291.360 ;
        RECT 595.775 290.910 597.580 291.250 ;
        RECT 596.220 290.890 597.580 290.910 ;
        RECT 596.950 290.510 597.580 290.890 ;
        RECT 634.040 291.320 635.600 291.360 ;
        RECT 634.040 290.870 634.320 291.320 ;
        RECT 379.040 275.800 379.370 276.020 ;
        RECT 385.660 276.010 385.940 289.790 ;
        RECT 631.320 289.670 632.060 290.280 ;
        RECT 633.820 290.190 634.530 290.870 ;
        RECT 636.075 290.305 636.405 291.380 ;
        RECT 610.200 288.470 610.370 288.890 ;
        RECT 610.990 288.470 611.160 288.890 ;
        RECT 611.780 288.470 611.950 288.890 ;
        RECT 612.570 288.470 612.740 288.890 ;
        RECT 613.360 288.470 613.530 288.890 ;
        RECT 617.790 288.440 617.960 288.860 ;
        RECT 618.580 288.440 618.750 288.860 ;
        RECT 619.370 288.440 619.540 288.860 ;
        RECT 620.160 288.440 620.330 288.860 ;
        RECT 620.950 288.440 621.120 288.860 ;
        RECT 600.750 287.690 600.920 288.110 ;
        RECT 601.540 287.690 601.710 288.110 ;
        RECT 602.330 287.690 602.500 288.110 ;
        RECT 603.120 287.690 603.290 288.110 ;
        RECT 603.910 287.690 604.080 288.110 ;
        RECT 615.310 287.960 615.790 288.380 ;
        RECT 627.530 287.820 627.700 288.240 ;
        RECT 628.320 287.820 628.490 288.240 ;
        RECT 629.110 287.820 629.280 288.240 ;
        RECT 629.900 287.820 630.070 288.240 ;
        RECT 630.690 287.820 630.860 288.240 ;
        RECT 591.820 285.440 592.170 287.600 ;
        RECT 637.280 287.450 637.680 291.380 ;
        RECT 640.265 290.395 640.595 291.510 ;
        RECT 641.750 291.170 641.980 291.510 ;
        RECT 643.475 291.430 644.185 291.510 ;
        RECT 644.365 291.610 644.695 292.055 ;
        RECT 645.260 291.610 645.570 291.630 ;
        RECT 644.365 291.430 645.570 291.610 ;
        RECT 641.680 290.850 642.060 291.170 ;
        RECT 644.365 290.375 644.695 291.430 ;
        RECT 645.260 291.280 645.570 291.430 ;
        RECT 820.140 291.375 820.310 291.975 ;
        RECT 819.655 291.205 821.715 291.375 ;
        RECT 694.770 288.550 696.160 290.530 ;
        RECT 819.065 290.475 819.475 291.145 ;
        RECT 819.655 290.295 819.825 291.205 ;
        RECT 821.385 291.025 821.715 291.205 ;
        RECT 819.070 290.125 819.825 290.295 ;
        RECT 819.070 289.795 819.320 290.125 ;
        RECT 820.005 290.110 820.395 291.025 ;
        RECT 821.920 290.720 822.195 293.055 ;
        RECT 832.760 292.130 834.110 293.070 ;
        RECT 839.520 292.805 839.770 293.135 ;
        RECT 840.455 293.120 840.845 294.035 ;
        RECT 842.370 292.805 842.645 296.065 ;
        RECT 855.925 295.465 856.335 296.135 ;
        RECT 856.515 295.285 856.685 296.195 ;
        RECT 858.245 296.015 858.575 296.195 ;
        RECT 855.930 295.115 856.685 295.285 ;
        RECT 855.930 294.785 856.180 295.115 ;
        RECT 856.865 295.100 857.255 296.015 ;
        RECT 858.780 295.760 859.055 298.045 ;
        RECT 858.780 295.500 859.070 295.760 ;
        RECT 858.780 294.785 859.055 295.500 ;
        RECT 845.490 292.735 845.740 293.335 ;
        RECT 845.490 292.565 847.865 292.735 ;
        RECT 832.760 291.830 837.310 292.130 ;
        RECT 845.695 292.080 846.025 292.385 ;
        RECT 843.820 291.890 846.025 292.080 ;
        RECT 832.760 291.630 834.110 291.830 ;
        RECT 821.890 290.350 822.210 290.720 ;
        RECT 821.920 289.795 822.195 290.350 ;
        RECT 825.590 289.205 825.760 289.805 ;
        RECT 827.370 289.310 827.645 290.885 ;
        RECT 830.060 289.755 830.310 290.905 ;
        RECT 832.640 290.275 832.810 290.905 ;
        RECT 834.830 290.275 835.080 290.905 ;
        RECT 832.640 290.105 835.080 290.275 ;
        RECT 832.640 289.935 832.810 290.105 ;
        RECT 832.990 289.755 834.650 289.925 ;
        RECT 830.060 289.585 833.160 289.755 ;
        RECT 824.560 288.975 824.880 289.090 ;
        RECT 825.105 289.035 827.165 289.205 ;
        RECT 824.515 288.305 824.925 288.975 ;
        RECT 825.105 288.125 825.275 289.035 ;
        RECT 826.835 288.855 827.165 289.035 ;
        RECT 827.370 288.970 827.840 289.310 ;
        RECT 824.520 287.955 825.275 288.125 ;
        RECT 639.640 287.450 640.090 287.550 ;
        RECT 610.200 287.000 610.370 287.420 ;
        RECT 610.990 287.000 611.160 287.420 ;
        RECT 611.780 287.000 611.950 287.420 ;
        RECT 612.570 287.000 612.740 287.420 ;
        RECT 613.360 287.000 613.530 287.420 ;
        RECT 614.030 286.950 614.200 287.370 ;
        RECT 615.610 286.950 615.780 287.370 ;
        RECT 617.190 286.950 617.360 287.370 ;
        RECT 617.790 286.970 617.960 287.390 ;
        RECT 618.580 286.970 618.750 287.390 ;
        RECT 619.370 286.970 619.540 287.390 ;
        RECT 620.160 286.970 620.330 287.390 ;
        RECT 620.950 286.970 621.120 287.390 ;
        RECT 637.280 287.260 640.090 287.450 ;
        RECT 637.280 287.250 637.680 287.260 ;
        RECT 600.750 286.220 600.920 286.640 ;
        RECT 601.540 286.220 601.710 286.640 ;
        RECT 602.330 286.220 602.500 286.640 ;
        RECT 603.120 286.220 603.290 286.640 ;
        RECT 603.910 286.220 604.080 286.640 ;
        RECT 608.320 286.530 608.990 286.840 ;
        RECT 622.910 286.420 623.600 286.970 ;
        RECT 639.640 286.860 640.090 287.260 ;
        RECT 643.700 286.920 644.120 287.600 ;
        RECT 821.890 287.380 822.165 287.895 ;
        RECT 824.520 287.625 824.770 287.955 ;
        RECT 825.455 287.940 825.845 288.855 ;
        RECT 827.370 287.625 827.645 288.970 ;
        RECT 830.060 288.745 830.310 289.585 ;
        RECT 830.490 288.925 831.440 289.205 ;
        RECT 831.975 288.925 833.165 289.300 ;
        RECT 831.270 288.745 831.440 288.925 ;
        RECT 833.345 288.745 833.645 288.985 ;
        RECT 830.060 288.575 831.090 288.745 ;
        RECT 831.270 288.655 833.645 288.745 ;
        RECT 831.270 288.575 833.515 288.655 ;
        RECT 830.840 287.645 831.090 288.575 ;
        RECT 833.895 288.475 834.300 289.575 ;
        RECT 834.480 289.145 834.650 289.755 ;
        RECT 834.830 289.325 835.080 290.105 ;
        RECT 834.480 288.815 834.810 289.145 ;
        RECT 833.780 287.645 834.300 288.475 ;
        RECT 836.970 288.690 837.290 291.830 ;
        RECT 842.380 290.360 842.655 290.945 ;
        RECT 843.820 290.360 844.050 291.890 ;
        RECT 845.695 291.835 846.025 291.890 ;
        RECT 846.270 291.655 846.440 292.565 ;
        RECT 847.535 292.385 847.865 292.565 ;
        RECT 846.620 291.835 846.950 292.385 ;
        RECT 848.070 292.330 848.325 294.415 ;
        RECT 849.040 292.330 849.870 292.530 ;
        RECT 848.070 292.140 849.870 292.330 ;
        RECT 846.270 291.155 846.600 291.655 ;
        RECT 848.070 291.155 848.325 292.140 ;
        RECT 849.040 291.780 849.870 292.140 ;
        RECT 858.820 291.850 859.095 292.515 ;
        RECT 861.580 292.465 861.830 293.065 ;
        RECT 861.580 292.295 863.955 292.465 ;
        RECT 861.785 291.850 862.115 292.115 ;
        RECT 858.820 291.670 862.115 291.850 ;
        RECT 857.040 290.835 857.210 291.435 ;
        RECT 856.555 290.665 858.615 290.835 ;
        RECT 855.965 290.370 856.375 290.605 ;
        RECT 842.380 290.170 844.050 290.360 ;
        RECT 840.600 289.265 840.770 289.865 ;
        RECT 840.115 289.095 842.175 289.265 ;
        RECT 839.525 288.690 839.935 289.035 ;
        RECT 836.970 288.470 839.935 288.690 ;
        RECT 836.970 288.360 837.350 288.470 ;
        RECT 839.525 288.365 839.935 288.470 ;
        RECT 836.980 288.040 837.350 288.360 ;
        RECT 840.115 288.185 840.285 289.095 ;
        RECT 841.845 288.915 842.175 289.095 ;
        RECT 821.880 287.050 822.165 287.380 ;
        RECT 627.530 286.350 627.700 286.770 ;
        RECT 628.320 286.350 628.490 286.770 ;
        RECT 629.110 286.350 629.280 286.770 ;
        RECT 629.900 286.350 630.070 286.770 ;
        RECT 630.690 286.350 630.860 286.770 ;
        RECT 639.380 286.060 639.550 286.480 ;
        RECT 643.430 286.110 643.600 286.530 ;
        RECT 820.110 286.215 820.280 286.815 ;
        RECT 819.625 286.045 821.685 286.215 ;
        RECT 606.450 285.480 606.620 285.900 ;
        RECT 607.240 285.480 607.410 285.900 ;
        RECT 608.030 285.480 608.200 285.900 ;
        RECT 608.820 285.480 608.990 285.900 ;
        RECT 609.610 285.480 609.780 285.900 ;
        RECT 610.200 285.530 610.370 285.950 ;
        RECT 610.990 285.530 611.160 285.950 ;
        RECT 611.780 285.530 611.950 285.950 ;
        RECT 612.570 285.530 612.740 285.950 ;
        RECT 613.360 285.530 613.530 285.950 ;
        RECT 614.030 285.480 614.200 285.900 ;
        RECT 615.610 285.480 615.780 285.900 ;
        RECT 617.190 285.480 617.360 285.900 ;
        RECT 617.790 285.500 617.960 285.920 ;
        RECT 618.580 285.500 618.750 285.920 ;
        RECT 619.370 285.500 619.540 285.920 ;
        RECT 620.160 285.500 620.330 285.920 ;
        RECT 620.950 285.500 621.120 285.920 ;
        RECT 621.540 285.480 621.710 285.900 ;
        RECT 622.330 285.480 622.500 285.900 ;
        RECT 623.120 285.480 623.290 285.900 ;
        RECT 623.910 285.480 624.080 285.900 ;
        RECT 624.700 285.480 624.870 285.900 ;
        RECT 819.035 285.880 819.445 285.985 ;
        RECT 819.020 285.400 819.445 285.880 ;
        RECT 819.035 285.315 819.445 285.400 ;
        RECT 819.625 285.135 819.795 286.045 ;
        RECT 821.355 285.865 821.685 286.045 ;
        RECT 601.930 284.540 602.880 285.010 ;
        RECT 819.040 284.965 819.795 285.135 ;
        RECT 819.040 284.635 819.290 284.965 ;
        RECT 819.975 284.950 820.365 285.865 ;
        RECT 821.890 284.635 822.165 287.050 ;
        RECT 836.990 285.760 837.340 288.040 ;
        RECT 839.530 288.015 840.285 288.185 ;
        RECT 839.530 287.685 839.780 288.015 ;
        RECT 840.465 288.000 840.855 288.915 ;
        RECT 842.380 287.685 842.655 290.170 ;
        RECT 843.820 290.140 844.050 290.170 ;
        RECT 854.950 289.950 856.375 290.370 ;
        RECT 854.980 285.760 855.280 289.950 ;
        RECT 855.965 289.935 856.375 289.950 ;
        RECT 856.555 289.755 856.725 290.665 ;
        RECT 858.285 290.485 858.615 290.665 ;
        RECT 855.970 289.585 856.725 289.755 ;
        RECT 855.970 289.255 856.220 289.585 ;
        RECT 856.905 289.570 857.295 290.485 ;
        RECT 858.820 289.255 859.095 291.670 ;
        RECT 861.785 291.565 862.115 291.670 ;
        RECT 862.360 291.385 862.530 292.295 ;
        RECT 863.625 292.115 863.955 292.295 ;
        RECT 862.710 292.110 863.040 292.115 ;
        RECT 862.710 291.790 863.050 292.110 ;
        RECT 864.160 292.090 864.415 294.145 ;
        RECT 865.130 292.090 866.340 292.460 ;
        RECT 864.140 291.890 866.340 292.090 ;
        RECT 862.710 291.565 863.040 291.790 ;
        RECT 862.360 290.885 862.690 291.385 ;
        RECT 864.160 290.885 864.415 291.890 ;
        RECT 865.130 291.740 866.340 291.890 ;
        RECT 836.990 285.360 855.310 285.760 ;
        RECT 857.110 285.435 857.280 286.035 ;
        RECT 591.820 282.280 592.170 284.440 ;
        RECT 679.520 280.835 679.770 281.985 ;
        RECT 682.100 281.355 682.270 281.985 ;
        RECT 684.290 281.355 684.540 281.985 ;
        RECT 682.100 281.185 684.540 281.355 ;
        RECT 682.100 281.015 682.270 281.185 ;
        RECT 682.450 280.835 684.110 281.005 ;
        RECT 679.520 280.665 682.620 280.835 ;
        RECT 679.520 279.825 679.770 280.665 ;
        RECT 679.950 280.005 680.900 280.285 ;
        RECT 680.730 279.825 680.900 280.005 ;
        RECT 682.805 279.825 683.105 280.065 ;
        RECT 679.520 279.655 680.550 279.825 ;
        RECT 680.730 279.735 683.105 279.825 ;
        RECT 680.730 279.655 682.975 279.735 ;
        RECT 632.340 277.530 633.560 278.800 ;
        RECT 680.300 278.725 680.550 279.655 ;
        RECT 683.355 279.555 683.760 280.655 ;
        RECT 683.940 280.225 684.110 280.835 ;
        RECT 684.290 280.405 684.540 281.185 ;
        RECT 696.800 280.845 697.050 281.995 ;
        RECT 699.380 281.365 699.550 281.995 ;
        RECT 701.570 281.365 701.820 281.995 ;
        RECT 699.380 281.195 701.820 281.365 ;
        RECT 699.380 281.025 699.550 281.195 ;
        RECT 699.730 280.845 701.390 281.015 ;
        RECT 696.800 280.675 699.900 280.845 ;
        RECT 683.940 279.895 684.270 280.225 ;
        RECT 696.800 279.835 697.050 280.675 ;
        RECT 697.230 280.015 698.180 280.295 ;
        RECT 698.010 279.835 698.180 280.015 ;
        RECT 700.085 279.940 700.385 280.075 ;
        RECT 700.085 279.835 700.400 279.940 ;
        RECT 696.800 279.665 697.830 279.835 ;
        RECT 698.010 279.700 700.400 279.835 ;
        RECT 698.010 279.665 700.255 279.700 ;
        RECT 683.240 278.725 683.760 279.555 ;
        RECT 697.580 278.735 697.830 279.665 ;
        RECT 700.635 279.565 701.040 280.665 ;
        RECT 701.220 280.235 701.390 280.845 ;
        RECT 701.570 280.415 701.820 281.195 ;
        RECT 714.570 280.845 714.820 281.995 ;
        RECT 717.150 281.365 717.320 281.995 ;
        RECT 719.340 281.365 719.590 281.995 ;
        RECT 717.150 281.195 719.590 281.365 ;
        RECT 717.150 281.025 717.320 281.195 ;
        RECT 717.500 280.845 719.160 281.015 ;
        RECT 714.570 280.675 717.670 280.845 ;
        RECT 701.220 279.905 701.550 280.235 ;
        RECT 714.570 279.835 714.820 280.675 ;
        RECT 715.000 280.015 715.950 280.295 ;
        RECT 715.780 279.835 715.950 280.015 ;
        RECT 717.855 279.835 718.155 280.075 ;
        RECT 714.570 279.665 715.600 279.835 ;
        RECT 715.780 279.745 718.155 279.835 ;
        RECT 715.780 279.710 718.140 279.745 ;
        RECT 715.780 279.665 718.025 279.710 ;
        RECT 700.520 278.735 701.040 279.565 ;
        RECT 715.350 278.735 715.600 279.665 ;
        RECT 718.405 279.565 718.810 280.665 ;
        RECT 718.990 280.235 719.160 280.845 ;
        RECT 719.340 280.415 719.590 281.195 ;
        RECT 731.810 280.845 732.060 281.995 ;
        RECT 734.390 281.365 734.560 281.995 ;
        RECT 736.580 281.365 736.830 281.995 ;
        RECT 734.390 281.195 736.830 281.365 ;
        RECT 734.390 281.025 734.560 281.195 ;
        RECT 734.740 280.845 736.400 281.015 ;
        RECT 731.810 280.675 734.910 280.845 ;
        RECT 718.990 279.905 719.320 280.235 ;
        RECT 731.810 279.835 732.060 280.675 ;
        RECT 732.240 280.015 733.190 280.295 ;
        RECT 733.020 279.835 733.190 280.015 ;
        RECT 735.095 279.835 735.395 280.075 ;
        RECT 731.810 279.665 732.840 279.835 ;
        RECT 733.020 279.745 735.395 279.835 ;
        RECT 733.020 279.740 735.380 279.745 ;
        RECT 733.020 279.665 735.265 279.740 ;
        RECT 718.290 278.735 718.810 279.565 ;
        RECT 732.590 278.735 732.840 279.665 ;
        RECT 735.645 279.565 736.050 280.665 ;
        RECT 736.230 280.235 736.400 280.845 ;
        RECT 736.580 280.415 736.830 281.195 ;
        RECT 749.290 280.855 749.540 282.005 ;
        RECT 751.870 281.375 752.040 282.005 ;
        RECT 754.060 281.375 754.310 282.005 ;
        RECT 800.490 281.625 800.875 283.205 ;
        RECT 751.870 281.205 754.310 281.375 ;
        RECT 751.870 281.035 752.040 281.205 ;
        RECT 752.220 280.855 753.880 281.025 ;
        RECT 749.290 280.685 752.390 280.855 ;
        RECT 736.230 279.905 736.560 280.235 ;
        RECT 749.290 279.845 749.540 280.685 ;
        RECT 749.720 280.025 750.670 280.305 ;
        RECT 750.500 279.845 750.670 280.025 ;
        RECT 752.575 279.845 752.875 280.085 ;
        RECT 749.290 279.675 750.320 279.845 ;
        RECT 750.500 279.755 752.875 279.845 ;
        RECT 750.500 279.700 752.860 279.755 ;
        RECT 750.500 279.675 752.745 279.700 ;
        RECT 735.530 278.735 736.050 279.565 ;
        RECT 750.070 278.745 750.320 279.675 ;
        RECT 753.125 279.575 753.530 280.675 ;
        RECT 753.710 280.245 753.880 280.855 ;
        RECT 754.060 280.425 754.310 281.205 ;
        RECT 799.655 281.000 800.365 281.385 ;
        RECT 800.545 281.270 800.875 281.625 ;
        RECT 819.480 281.715 819.730 282.865 ;
        RECT 822.060 282.235 822.230 282.865 ;
        RECT 824.250 282.235 824.500 282.865 ;
        RECT 822.060 282.065 824.500 282.235 ;
        RECT 822.060 281.895 822.230 282.065 ;
        RECT 822.410 281.715 824.070 281.885 ;
        RECT 802.040 281.270 802.970 281.550 ;
        RECT 800.545 280.910 802.970 281.270 ;
        RECT 753.710 279.915 754.040 280.245 ;
        RECT 800.545 279.945 800.875 280.910 ;
        RECT 802.040 280.560 802.970 280.910 ;
        RECT 819.480 281.545 822.580 281.715 ;
        RECT 819.480 280.705 819.730 281.545 ;
        RECT 821.730 281.260 822.110 281.360 ;
        RECT 819.910 280.885 820.860 281.165 ;
        RECT 821.395 280.885 822.585 281.260 ;
        RECT 820.690 280.850 820.860 280.885 ;
        RECT 820.690 280.705 821.160 280.850 ;
        RECT 822.765 280.705 823.065 280.945 ;
        RECT 819.480 280.535 820.510 280.705 ;
        RECT 820.690 280.615 823.065 280.705 ;
        RECT 820.690 280.535 822.935 280.615 ;
        RECT 820.260 279.605 820.510 280.535 ;
        RECT 823.315 280.435 823.720 281.535 ;
        RECT 823.900 281.105 824.070 281.715 ;
        RECT 824.250 281.285 824.500 282.065 ;
        RECT 823.900 280.775 824.230 281.105 ;
        RECT 829.160 281.095 829.330 281.695 ;
        RECT 825.320 280.830 826.030 281.080 ;
        RECT 828.675 280.925 830.735 281.095 ;
        RECT 825.280 280.620 826.030 280.830 ;
        RECT 828.085 280.730 828.495 280.865 ;
        RECT 823.200 279.605 823.720 280.435 ;
        RECT 825.320 280.360 826.030 280.620 ;
        RECT 828.080 280.270 828.495 280.730 ;
        RECT 828.085 280.195 828.495 280.270 ;
        RECT 828.675 280.015 828.845 280.925 ;
        RECT 830.405 280.745 830.735 280.925 ;
        RECT 828.090 279.845 828.845 280.015 ;
        RECT 753.010 278.745 753.530 279.575 ;
        RECT 828.090 279.515 828.340 279.845 ;
        RECT 829.025 279.830 829.415 280.745 ;
        RECT 830.940 279.515 831.215 282.775 ;
        RECT 833.380 281.625 833.630 282.775 ;
        RECT 835.960 282.145 836.130 282.775 ;
        RECT 838.150 282.145 838.400 282.775 ;
        RECT 835.960 281.975 838.400 282.145 ;
        RECT 835.960 281.805 836.130 281.975 ;
        RECT 836.310 281.625 837.970 281.795 ;
        RECT 833.380 281.455 836.480 281.625 ;
        RECT 833.380 280.615 833.630 281.455 ;
        RECT 833.810 280.795 834.760 281.075 ;
        RECT 835.295 280.795 836.485 281.170 ;
        RECT 834.590 280.615 834.760 280.795 ;
        RECT 836.660 280.615 836.990 280.900 ;
        RECT 833.380 280.445 834.410 280.615 ;
        RECT 834.590 280.580 836.990 280.615 ;
        RECT 834.590 280.525 836.965 280.580 ;
        RECT 834.590 280.445 836.835 280.525 ;
        RECT 834.160 279.515 834.410 280.445 ;
        RECT 837.215 280.345 837.620 281.445 ;
        RECT 837.800 281.015 837.970 281.625 ;
        RECT 838.150 281.195 838.400 281.975 ;
        RECT 840.590 281.015 840.840 282.065 ;
        RECT 841.080 281.510 841.440 281.520 ;
        RECT 841.065 281.195 842.025 281.510 ;
        RECT 842.230 281.015 842.480 282.065 ;
        RECT 843.825 281.195 844.175 282.775 ;
        RECT 843.870 281.180 844.175 281.195 ;
        RECT 846.430 281.625 846.680 282.775 ;
        RECT 849.010 282.145 849.180 282.775 ;
        RECT 851.200 282.145 851.450 282.775 ;
        RECT 849.010 281.975 851.450 282.145 ;
        RECT 849.010 281.805 849.180 281.975 ;
        RECT 849.360 281.625 851.020 281.795 ;
        RECT 846.430 281.455 849.530 281.625 ;
        RECT 837.800 280.685 838.130 281.015 ;
        RECT 840.590 280.845 843.700 281.015 ;
        RECT 837.100 279.515 837.620 280.345 ;
        RECT 838.650 280.340 839.040 280.620 ;
        RECT 838.740 279.530 838.910 280.340 ;
        RECT 840.590 279.845 840.885 280.845 ;
        RECT 843.370 280.685 843.700 280.845 ;
        RECT 843.870 280.890 844.230 281.180 ;
        RECT 841.065 280.570 841.395 280.665 ;
        RECT 841.065 280.300 841.400 280.570 ;
        RECT 841.065 279.830 841.395 280.300 ;
        RECT 841.575 279.830 842.715 280.665 ;
        RECT 838.730 278.120 838.910 279.530 ;
        RECT 843.870 279.515 844.175 280.890 ;
        RECT 846.430 280.615 846.680 281.455 ;
        RECT 846.860 280.795 847.810 281.075 ;
        RECT 848.345 280.795 849.535 281.170 ;
        RECT 849.740 280.855 850.020 281.010 ;
        RECT 847.640 280.615 847.810 280.795 ;
        RECT 849.715 280.615 850.020 280.855 ;
        RECT 846.430 280.445 847.460 280.615 ;
        RECT 847.640 280.590 850.020 280.615 ;
        RECT 847.640 280.525 850.015 280.590 ;
        RECT 847.640 280.445 849.885 280.525 ;
        RECT 847.210 279.515 847.460 280.445 ;
        RECT 850.265 280.345 850.670 281.445 ;
        RECT 850.850 281.015 851.020 281.625 ;
        RECT 851.200 281.195 851.450 281.975 ;
        RECT 850.850 280.685 851.180 281.015 ;
        RECT 850.150 279.515 850.670 280.345 ;
        RECT 854.980 279.370 855.280 285.360 ;
        RECT 856.625 285.265 858.685 285.435 ;
        RECT 856.035 284.535 856.445 285.205 ;
        RECT 856.625 284.355 856.795 285.265 ;
        RECT 858.355 285.085 858.685 285.265 ;
        RECT 856.040 284.185 856.795 284.355 ;
        RECT 856.040 283.855 856.290 284.185 ;
        RECT 856.975 284.170 857.365 285.085 ;
        RECT 858.890 283.855 859.165 287.115 ;
        RECT 861.660 283.415 861.910 284.015 ;
        RECT 861.660 283.245 864.035 283.415 ;
        RECT 861.865 282.990 862.195 283.065 ;
        RECT 861.860 282.710 862.195 282.990 ;
        RECT 861.865 282.515 862.195 282.710 ;
        RECT 862.440 282.335 862.610 283.245 ;
        RECT 863.705 283.065 864.035 283.245 ;
        RECT 862.790 282.515 863.120 283.065 ;
        RECT 864.240 283.040 864.495 285.095 ;
        RECT 865.160 283.040 865.910 283.170 ;
        RECT 864.240 282.840 865.910 283.040 ;
        RECT 862.440 281.835 862.770 282.335 ;
        RECT 864.240 281.835 864.495 282.840 ;
        RECT 865.160 282.670 865.910 282.840 ;
        RECT 857.130 279.975 857.300 280.575 ;
        RECT 856.645 279.805 858.705 279.975 ;
        RECT 856.055 279.370 856.465 279.745 ;
        RECT 854.980 279.080 856.465 279.370 ;
        RECT 854.980 279.030 855.280 279.080 ;
        RECT 856.055 279.075 856.465 279.080 ;
        RECT 851.770 278.120 852.380 278.150 ;
        RECT 838.730 278.070 839.120 278.120 ;
        RECT 839.450 278.080 841.600 278.120 ;
        RECT 842.000 278.080 852.380 278.120 ;
        RECT 839.450 278.070 852.380 278.080 ;
        RECT 838.730 277.830 852.380 278.070 ;
        RECT 851.940 277.530 852.380 277.830 ;
        RECT 852.000 277.510 852.340 277.530 ;
        RECT 603.140 276.230 603.310 276.650 ;
        RECT 604.720 276.230 604.890 276.650 ;
        RECT 607.660 276.240 607.830 276.660 ;
        RECT 609.240 276.240 609.410 276.660 ;
        RECT 612.180 276.240 612.350 276.660 ;
        RECT 613.760 276.240 613.930 276.660 ;
        RECT 616.610 276.220 616.780 276.640 ;
        RECT 618.190 276.220 618.360 276.640 ;
        RECT 620.990 276.230 621.160 276.650 ;
        RECT 622.570 276.230 622.740 276.650 ;
        RECT 625.310 276.220 625.480 276.640 ;
        RECT 626.890 276.220 627.060 276.640 ;
        RECT 379.040 274.810 379.340 275.800 ;
        RECT 385.660 275.570 385.980 276.010 ;
        RECT 385.680 274.830 385.980 275.570 ;
        RECT 385.680 274.810 386.470 274.830 ;
        RECT 379.040 274.500 386.470 274.810 ;
        RECT 603.140 274.760 603.310 275.180 ;
        RECT 604.720 274.760 604.890 275.180 ;
        RECT 607.660 274.770 607.830 275.190 ;
        RECT 609.240 274.770 609.410 275.190 ;
        RECT 612.180 274.770 612.350 275.190 ;
        RECT 613.760 274.770 613.930 275.190 ;
        RECT 616.610 274.750 616.780 275.170 ;
        RECT 618.190 274.750 618.360 275.170 ;
        RECT 620.990 274.760 621.160 275.180 ;
        RECT 622.570 274.760 622.740 275.180 ;
        RECT 625.310 274.750 625.480 275.170 ;
        RECT 626.890 274.750 627.060 275.170 ;
        RECT 379.040 274.470 379.340 274.500 ;
        RECT 385.680 274.460 385.980 274.500 ;
        RECT 595.185 273.065 595.570 274.645 ;
        RECT 613.230 273.810 613.700 274.190 ;
        RECT 616.070 273.770 616.500 274.090 ;
        RECT 620.480 273.910 620.890 274.340 ;
        RECT 635.940 273.515 636.325 275.095 ;
        RECT 640.130 273.605 640.515 275.185 ;
        RECT 679.930 275.175 680.180 276.325 ;
        RECT 682.510 275.695 682.680 276.325 ;
        RECT 684.700 275.695 684.950 276.325 ;
        RECT 682.510 275.525 684.950 275.695 ;
        RECT 682.510 275.355 682.680 275.525 ;
        RECT 682.860 275.175 684.520 275.345 ;
        RECT 635.105 273.260 635.815 273.275 ;
        RECT 594.190 272.730 594.870 272.820 ;
        RECT 595.185 272.730 595.515 273.065 ;
        RECT 633.960 272.890 635.815 273.260 ;
        RECT 635.995 273.190 636.325 273.515 ;
        RECT 639.120 273.365 639.490 273.390 ;
        RECT 636.750 273.190 637.590 273.200 ;
        RECT 635.995 273.150 637.590 273.190 ;
        RECT 635.995 272.910 637.600 273.150 ;
        RECT 639.120 272.980 640.005 273.365 ;
        RECT 640.185 273.250 640.515 273.605 ;
        RECT 644.230 273.585 644.615 275.165 ;
        RECT 679.930 275.005 683.030 275.175 ;
        RECT 679.930 274.165 680.180 275.005 ;
        RECT 680.360 274.345 681.310 274.625 ;
        RECT 681.845 274.345 683.035 274.720 ;
        RECT 681.140 274.165 681.310 274.345 ;
        RECT 683.215 274.165 683.515 274.405 ;
        RECT 679.930 273.995 680.960 274.165 ;
        RECT 681.140 274.075 683.515 274.165 ;
        RECT 681.140 273.995 683.385 274.075 ;
        RECT 643.395 273.250 644.105 273.345 ;
        RECT 640.185 273.040 644.105 273.250 ;
        RECT 639.120 272.940 639.490 272.980 ;
        RECT 594.190 272.490 595.515 272.730 ;
        RECT 594.190 272.420 594.870 272.490 ;
        RECT 595.185 271.385 595.515 272.490 ;
        RECT 595.695 272.780 596.405 272.825 ;
        RECT 596.870 272.780 597.500 272.890 ;
        RECT 595.695 272.440 597.500 272.780 ;
        RECT 596.140 272.420 597.500 272.440 ;
        RECT 596.870 272.040 597.500 272.420 ;
        RECT 633.960 272.850 635.520 272.890 ;
        RECT 633.960 272.400 634.240 272.850 ;
        RECT 379.160 271.160 379.330 271.320 ;
        RECT 379.110 257.160 379.390 271.160 ;
        RECT 385.740 270.930 385.910 271.320 ;
        RECT 631.440 271.070 632.060 271.730 ;
        RECT 633.740 271.720 634.450 272.400 ;
        RECT 635.995 271.835 636.325 272.910 ;
        RECT 379.060 256.940 379.390 257.160 ;
        RECT 385.680 257.150 385.960 270.930 ;
        RECT 610.120 270.000 610.290 270.420 ;
        RECT 610.910 270.000 611.080 270.420 ;
        RECT 611.700 270.000 611.870 270.420 ;
        RECT 612.490 270.000 612.660 270.420 ;
        RECT 613.280 270.000 613.450 270.420 ;
        RECT 617.710 269.970 617.880 270.390 ;
        RECT 618.500 269.970 618.670 270.390 ;
        RECT 619.290 269.970 619.460 270.390 ;
        RECT 620.080 269.970 620.250 270.390 ;
        RECT 620.870 269.970 621.040 270.390 ;
        RECT 591.660 267.180 592.010 269.340 ;
        RECT 600.670 269.220 600.840 269.640 ;
        RECT 601.460 269.220 601.630 269.640 ;
        RECT 602.250 269.220 602.420 269.640 ;
        RECT 603.040 269.220 603.210 269.640 ;
        RECT 603.830 269.220 604.000 269.640 ;
        RECT 615.230 269.490 615.710 269.910 ;
        RECT 627.450 269.350 627.620 269.770 ;
        RECT 628.240 269.350 628.410 269.770 ;
        RECT 629.030 269.350 629.200 269.770 ;
        RECT 629.820 269.350 629.990 269.770 ;
        RECT 630.610 269.350 630.780 269.770 ;
        RECT 637.200 268.980 637.600 272.910 ;
        RECT 640.185 271.925 640.515 273.040 ;
        RECT 641.670 272.700 641.900 273.040 ;
        RECT 643.395 272.960 644.105 273.040 ;
        RECT 644.285 273.140 644.615 273.585 ;
        RECT 645.180 273.140 645.490 273.160 ;
        RECT 644.285 272.960 645.490 273.140 ;
        RECT 680.710 273.065 680.960 273.995 ;
        RECT 683.765 273.895 684.170 274.995 ;
        RECT 684.350 274.565 684.520 275.175 ;
        RECT 684.700 274.745 684.950 275.525 ;
        RECT 687.170 275.135 687.420 276.285 ;
        RECT 689.750 275.655 689.920 276.285 ;
        RECT 691.940 275.655 692.190 276.285 ;
        RECT 689.750 275.485 692.190 275.655 ;
        RECT 689.750 275.315 689.920 275.485 ;
        RECT 690.100 275.135 691.760 275.305 ;
        RECT 687.170 274.965 690.270 275.135 ;
        RECT 684.350 274.235 684.680 274.565 ;
        RECT 687.170 274.125 687.420 274.965 ;
        RECT 687.600 274.305 688.550 274.585 ;
        RECT 689.085 274.305 690.275 274.680 ;
        RECT 688.380 274.125 688.550 274.305 ;
        RECT 690.455 274.125 690.755 274.365 ;
        RECT 687.170 273.955 688.200 274.125 ;
        RECT 688.380 274.035 690.755 274.125 ;
        RECT 688.380 273.955 690.625 274.035 ;
        RECT 683.650 273.065 684.170 273.895 ;
        RECT 687.950 273.025 688.200 273.955 ;
        RECT 691.005 273.855 691.410 274.955 ;
        RECT 691.590 274.525 691.760 275.135 ;
        RECT 691.940 274.705 692.190 275.485 ;
        RECT 697.160 275.195 697.410 276.345 ;
        RECT 699.740 275.715 699.910 276.345 ;
        RECT 701.930 275.715 702.180 276.345 ;
        RECT 699.740 275.545 702.180 275.715 ;
        RECT 699.740 275.375 699.910 275.545 ;
        RECT 700.090 275.195 701.750 275.365 ;
        RECT 697.160 275.025 700.260 275.195 ;
        RECT 691.590 274.195 691.920 274.525 ;
        RECT 697.160 274.185 697.410 275.025 ;
        RECT 697.590 274.365 698.540 274.645 ;
        RECT 698.370 274.185 698.540 274.365 ;
        RECT 700.445 274.185 700.745 274.425 ;
        RECT 697.160 274.015 698.190 274.185 ;
        RECT 698.370 274.095 700.745 274.185 ;
        RECT 698.370 274.015 700.615 274.095 ;
        RECT 690.890 273.025 691.410 273.855 ;
        RECT 697.940 273.085 698.190 274.015 ;
        RECT 700.995 273.915 701.400 275.015 ;
        RECT 701.580 274.585 701.750 275.195 ;
        RECT 701.930 274.765 702.180 275.545 ;
        RECT 704.400 275.155 704.650 276.305 ;
        RECT 706.980 275.675 707.150 276.305 ;
        RECT 709.170 275.675 709.420 276.305 ;
        RECT 706.980 275.505 709.420 275.675 ;
        RECT 706.980 275.335 707.150 275.505 ;
        RECT 707.330 275.155 708.990 275.325 ;
        RECT 704.400 274.985 707.500 275.155 ;
        RECT 701.580 274.255 701.910 274.585 ;
        RECT 704.400 274.145 704.650 274.985 ;
        RECT 704.830 274.325 705.780 274.605 ;
        RECT 706.315 274.325 707.505 274.700 ;
        RECT 705.610 274.145 705.780 274.325 ;
        RECT 707.685 274.145 707.985 274.385 ;
        RECT 704.400 273.975 705.430 274.145 ;
        RECT 705.610 274.055 707.985 274.145 ;
        RECT 705.610 273.975 707.855 274.055 ;
        RECT 700.880 273.085 701.400 273.915 ;
        RECT 705.180 273.045 705.430 273.975 ;
        RECT 708.235 273.875 708.640 274.975 ;
        RECT 708.820 274.545 708.990 275.155 ;
        RECT 709.170 274.725 709.420 275.505 ;
        RECT 714.730 275.295 714.980 276.445 ;
        RECT 717.310 275.815 717.480 276.445 ;
        RECT 719.500 275.815 719.750 276.445 ;
        RECT 717.310 275.645 719.750 275.815 ;
        RECT 717.310 275.475 717.480 275.645 ;
        RECT 717.660 275.295 719.320 275.465 ;
        RECT 714.730 275.125 717.830 275.295 ;
        RECT 708.820 274.215 709.150 274.545 ;
        RECT 714.730 274.285 714.980 275.125 ;
        RECT 715.160 274.465 716.110 274.745 ;
        RECT 715.940 274.285 716.110 274.465 ;
        RECT 718.015 274.285 718.315 274.525 ;
        RECT 714.730 274.115 715.760 274.285 ;
        RECT 715.940 274.195 718.315 274.285 ;
        RECT 715.940 274.115 718.185 274.195 ;
        RECT 708.120 273.045 708.640 273.875 ;
        RECT 715.510 273.185 715.760 274.115 ;
        RECT 718.565 274.015 718.970 275.115 ;
        RECT 719.150 274.685 719.320 275.295 ;
        RECT 719.500 274.865 719.750 275.645 ;
        RECT 721.970 275.255 722.220 276.405 ;
        RECT 724.550 275.775 724.720 276.405 ;
        RECT 726.740 275.775 726.990 276.405 ;
        RECT 724.550 275.605 726.990 275.775 ;
        RECT 724.550 275.435 724.720 275.605 ;
        RECT 724.900 275.255 726.560 275.425 ;
        RECT 721.970 275.085 725.070 275.255 ;
        RECT 719.150 274.355 719.480 274.685 ;
        RECT 721.970 274.245 722.220 275.085 ;
        RECT 722.400 274.425 723.350 274.705 ;
        RECT 723.885 274.425 725.075 274.800 ;
        RECT 723.180 274.245 723.350 274.425 ;
        RECT 725.255 274.245 725.555 274.485 ;
        RECT 721.970 274.075 723.000 274.245 ;
        RECT 723.180 274.155 725.555 274.245 ;
        RECT 723.180 274.075 725.425 274.155 ;
        RECT 718.450 273.185 718.970 274.015 ;
        RECT 722.750 273.145 723.000 274.075 ;
        RECT 725.805 273.975 726.210 275.075 ;
        RECT 726.390 274.645 726.560 275.255 ;
        RECT 726.740 274.825 726.990 275.605 ;
        RECT 731.900 275.325 732.150 276.475 ;
        RECT 734.480 275.845 734.650 276.475 ;
        RECT 736.670 275.845 736.920 276.475 ;
        RECT 734.480 275.675 736.920 275.845 ;
        RECT 734.480 275.505 734.650 275.675 ;
        RECT 734.830 275.325 736.490 275.495 ;
        RECT 731.900 275.155 735.000 275.325 ;
        RECT 726.390 274.315 726.720 274.645 ;
        RECT 731.900 274.315 732.150 275.155 ;
        RECT 732.330 274.495 733.280 274.775 ;
        RECT 733.110 274.315 733.280 274.495 ;
        RECT 735.185 274.315 735.485 274.555 ;
        RECT 731.900 274.145 732.930 274.315 ;
        RECT 733.110 274.225 735.485 274.315 ;
        RECT 733.110 274.145 735.355 274.225 ;
        RECT 725.690 273.145 726.210 273.975 ;
        RECT 732.680 273.215 732.930 274.145 ;
        RECT 735.735 274.045 736.140 275.145 ;
        RECT 736.320 274.715 736.490 275.325 ;
        RECT 736.670 274.895 736.920 275.675 ;
        RECT 739.140 275.285 739.390 276.435 ;
        RECT 741.720 275.805 741.890 276.435 ;
        RECT 743.910 275.805 744.160 276.435 ;
        RECT 741.720 275.635 744.160 275.805 ;
        RECT 741.720 275.465 741.890 275.635 ;
        RECT 742.070 275.285 743.730 275.455 ;
        RECT 739.140 275.115 742.240 275.285 ;
        RECT 736.320 274.385 736.650 274.715 ;
        RECT 739.140 274.275 739.390 275.115 ;
        RECT 739.570 274.455 740.520 274.735 ;
        RECT 741.055 274.455 742.245 274.830 ;
        RECT 740.350 274.275 740.520 274.455 ;
        RECT 742.425 274.275 742.725 274.515 ;
        RECT 739.140 274.105 740.170 274.275 ;
        RECT 740.350 274.185 742.725 274.275 ;
        RECT 740.350 274.105 742.595 274.185 ;
        RECT 735.620 273.215 736.140 274.045 ;
        RECT 739.920 273.175 740.170 274.105 ;
        RECT 742.975 274.005 743.380 275.105 ;
        RECT 743.560 274.675 743.730 275.285 ;
        RECT 743.910 274.855 744.160 275.635 ;
        RECT 749.710 275.385 749.960 276.535 ;
        RECT 752.290 275.905 752.460 276.535 ;
        RECT 754.480 275.905 754.730 276.535 ;
        RECT 752.290 275.735 754.730 275.905 ;
        RECT 752.290 275.565 752.460 275.735 ;
        RECT 752.640 275.385 754.300 275.555 ;
        RECT 749.710 275.215 752.810 275.385 ;
        RECT 743.560 274.345 743.890 274.675 ;
        RECT 749.710 274.375 749.960 275.215 ;
        RECT 750.140 274.555 751.090 274.835 ;
        RECT 750.920 274.375 751.090 274.555 ;
        RECT 752.995 274.375 753.295 274.615 ;
        RECT 749.710 274.205 750.740 274.375 ;
        RECT 750.920 274.285 753.295 274.375 ;
        RECT 750.920 274.205 753.165 274.285 ;
        RECT 742.860 273.175 743.380 274.005 ;
        RECT 750.490 273.275 750.740 274.205 ;
        RECT 753.545 274.105 753.950 275.205 ;
        RECT 754.130 274.775 754.300 275.385 ;
        RECT 754.480 274.955 754.730 275.735 ;
        RECT 756.950 275.345 757.200 276.495 ;
        RECT 759.530 275.865 759.700 276.495 ;
        RECT 761.720 275.865 761.970 276.495 ;
        RECT 759.530 275.695 761.970 275.865 ;
        RECT 759.530 275.525 759.700 275.695 ;
        RECT 759.880 275.345 761.540 275.515 ;
        RECT 756.950 275.175 760.050 275.345 ;
        RECT 754.130 274.445 754.460 274.775 ;
        RECT 756.950 274.335 757.200 275.175 ;
        RECT 758.865 274.515 760.055 274.890 ;
        RECT 756.950 274.165 757.980 274.335 ;
        RECT 753.430 273.275 753.950 274.105 ;
        RECT 757.730 273.235 757.980 274.165 ;
        RECT 760.785 274.065 761.190 275.165 ;
        RECT 761.370 274.735 761.540 275.345 ;
        RECT 761.720 274.915 761.970 275.695 ;
        RECT 852.040 275.360 852.340 277.510 ;
        RECT 782.360 275.045 783.800 275.215 ;
        RECT 761.370 274.405 761.700 274.735 ;
        RECT 760.670 273.235 761.190 274.065 ;
        RECT 781.070 273.935 781.400 274.865 ;
        RECT 782.360 273.935 782.530 275.045 ;
        RECT 781.070 273.765 782.530 273.935 ;
        RECT 641.600 272.380 641.980 272.700 ;
        RECT 644.285 271.905 644.615 272.960 ;
        RECT 645.180 272.810 645.490 272.960 ;
        RECT 645.850 271.320 646.500 272.630 ;
        RECT 781.070 271.905 781.340 273.765 ;
        RECT 782.200 273.265 782.530 273.765 ;
        RECT 782.710 273.560 782.960 274.865 ;
        RECT 783.200 274.250 783.450 274.865 ;
        RECT 783.630 274.600 783.800 275.045 ;
        RECT 784.490 275.045 786.230 275.215 ;
        RECT 784.490 274.600 784.660 275.045 ;
        RECT 783.630 274.430 784.660 274.600 ;
        RECT 784.840 274.250 785.010 274.865 ;
        RECT 785.540 274.610 785.870 274.865 ;
        RECT 783.200 274.080 785.010 274.250 ;
        RECT 785.190 274.080 785.410 274.410 ;
        RECT 784.840 273.900 785.010 274.080 ;
        RECT 784.840 273.730 785.060 273.900 ;
        RECT 782.710 273.330 783.235 273.560 ;
        RECT 782.710 272.405 782.980 273.330 ;
        RECT 784.375 272.600 784.705 273.515 ;
        RECT 782.650 271.905 782.980 272.405 ;
        RECT 784.370 272.250 784.705 272.600 ;
        RECT 784.375 272.220 784.705 272.250 ;
        RECT 784.890 272.735 785.060 273.730 ;
        RECT 785.240 273.560 785.410 274.080 ;
        RECT 785.590 273.910 785.760 274.610 ;
        RECT 786.060 274.455 786.230 275.045 ;
        RECT 787.540 275.045 788.570 275.215 ;
        RECT 787.540 274.455 787.710 275.045 ;
        RECT 786.060 274.410 787.710 274.455 ;
        RECT 785.940 274.285 787.710 274.410 ;
        RECT 785.940 274.090 786.270 274.285 ;
        RECT 787.890 274.105 788.220 274.865 ;
        RECT 788.400 274.685 788.570 275.045 ;
        RECT 788.400 274.515 790.210 274.685 ;
        RECT 786.450 273.935 788.220 274.105 ;
        RECT 786.450 273.910 786.620 273.935 ;
        RECT 785.590 273.740 786.620 273.910 ;
        RECT 789.530 273.755 789.860 274.335 ;
        RECT 785.240 273.330 786.265 273.560 ;
        RECT 785.935 272.835 786.265 273.330 ;
        RECT 786.450 273.055 786.620 273.740 ;
        RECT 786.800 273.585 789.860 273.755 ;
        RECT 786.800 273.235 787.130 273.585 ;
        RECT 786.450 272.885 789.070 273.055 ;
        RECT 784.890 272.235 785.160 272.735 ;
        RECT 786.450 272.655 786.620 272.885 ;
        RECT 785.610 272.485 786.620 272.655 ;
        RECT 789.600 272.735 789.860 273.585 ;
        RECT 790.040 273.165 790.210 274.515 ;
        RECT 790.390 274.255 790.640 275.165 ;
        RECT 790.390 274.085 791.265 274.255 ;
        RECT 790.585 273.345 790.915 273.845 ;
        RECT 791.095 273.765 791.265 274.085 ;
        RECT 792.800 274.115 793.050 274.585 ;
        RECT 792.800 273.945 793.805 274.115 ;
        RECT 791.095 273.595 793.455 273.765 ;
        RECT 790.040 272.995 791.210 273.165 ;
        RECT 785.610 272.235 785.940 272.485 ;
        RECT 789.600 272.025 789.930 272.735 ;
        RECT 790.390 272.195 790.720 272.735 ;
        RECT 790.925 272.495 791.210 272.995 ;
        RECT 791.390 272.195 791.560 273.595 ;
        RECT 793.635 273.415 793.805 273.945 ;
        RECT 791.765 273.245 793.805 273.415 ;
        RECT 791.765 272.855 792.095 273.245 ;
        RECT 790.390 272.025 791.560 272.195 ;
        RECT 793.580 272.405 793.805 273.245 ;
        RECT 794.305 273.415 794.555 274.415 ;
        RECT 794.305 273.085 795.680 273.415 ;
        RECT 794.305 272.905 794.515 273.085 ;
        RECT 794.185 272.405 794.515 272.905 ;
        RECT 793.580 271.905 793.910 272.405 ;
        RECT 795.860 272.075 796.195 275.145 ;
        RECT 801.250 275.035 802.690 275.205 ;
        RECT 799.960 273.925 800.290 274.855 ;
        RECT 801.250 273.925 801.420 275.035 ;
        RECT 799.960 273.755 801.420 273.925 ;
        RECT 799.960 271.895 800.230 273.755 ;
        RECT 801.090 273.255 801.420 273.755 ;
        RECT 801.600 273.550 801.850 274.855 ;
        RECT 802.090 274.240 802.340 274.855 ;
        RECT 802.520 274.590 802.690 275.035 ;
        RECT 803.380 275.035 805.120 275.205 ;
        RECT 803.380 274.590 803.550 275.035 ;
        RECT 802.520 274.420 803.550 274.590 ;
        RECT 803.730 274.240 803.900 274.855 ;
        RECT 804.430 274.600 804.760 274.855 ;
        RECT 802.090 274.070 803.900 274.240 ;
        RECT 804.080 274.070 804.300 274.400 ;
        RECT 803.730 273.890 803.900 274.070 ;
        RECT 803.730 273.720 803.950 273.890 ;
        RECT 801.600 273.320 802.125 273.550 ;
        RECT 801.600 272.395 801.870 273.320 ;
        RECT 801.540 271.895 801.870 272.395 ;
        RECT 803.265 272.210 803.595 273.505 ;
        RECT 803.780 272.725 803.950 273.720 ;
        RECT 804.130 273.550 804.300 274.070 ;
        RECT 804.480 273.900 804.650 274.600 ;
        RECT 804.950 274.445 805.120 275.035 ;
        RECT 806.430 275.035 807.460 275.205 ;
        RECT 806.430 274.445 806.600 275.035 ;
        RECT 804.950 274.400 806.600 274.445 ;
        RECT 804.830 274.275 806.600 274.400 ;
        RECT 804.830 274.080 805.160 274.275 ;
        RECT 806.780 274.095 807.110 274.855 ;
        RECT 807.290 274.675 807.460 275.035 ;
        RECT 807.290 274.505 809.100 274.675 ;
        RECT 805.340 273.925 807.110 274.095 ;
        RECT 805.340 273.900 805.510 273.925 ;
        RECT 804.480 273.730 805.510 273.900 ;
        RECT 808.420 273.745 808.750 274.325 ;
        RECT 804.130 273.320 805.155 273.550 ;
        RECT 804.825 272.825 805.155 273.320 ;
        RECT 805.340 273.045 805.510 273.730 ;
        RECT 805.690 273.575 808.750 273.745 ;
        RECT 805.690 273.225 806.020 273.575 ;
        RECT 805.340 272.875 807.960 273.045 ;
        RECT 803.780 272.225 804.050 272.725 ;
        RECT 805.340 272.645 805.510 272.875 ;
        RECT 804.500 272.475 805.510 272.645 ;
        RECT 808.490 272.725 808.750 273.575 ;
        RECT 808.930 273.155 809.100 274.505 ;
        RECT 809.280 274.245 809.530 275.155 ;
        RECT 809.280 274.075 810.155 274.245 ;
        RECT 809.475 273.335 809.805 273.835 ;
        RECT 809.985 273.755 810.155 274.075 ;
        RECT 811.690 274.105 811.940 274.575 ;
        RECT 811.690 273.935 812.695 274.105 ;
        RECT 809.985 273.585 812.345 273.755 ;
        RECT 808.930 272.985 810.100 273.155 ;
        RECT 804.500 272.225 804.830 272.475 ;
        RECT 808.490 272.015 808.820 272.725 ;
        RECT 809.280 272.185 809.610 272.725 ;
        RECT 809.815 272.485 810.100 272.985 ;
        RECT 810.280 272.185 810.450 273.585 ;
        RECT 812.525 273.405 812.695 273.935 ;
        RECT 810.655 273.235 812.695 273.405 ;
        RECT 810.655 272.845 810.985 273.235 ;
        RECT 809.280 272.015 810.450 272.185 ;
        RECT 812.470 272.395 812.695 273.235 ;
        RECT 813.195 273.405 813.445 274.405 ;
        RECT 813.195 273.075 814.570 273.405 ;
        RECT 813.195 272.895 813.405 273.075 ;
        RECT 813.075 272.395 813.405 272.895 ;
        RECT 812.470 271.895 812.800 272.395 ;
        RECT 814.750 272.065 815.085 275.135 ;
        RECT 820.100 275.005 821.540 275.175 ;
        RECT 818.810 273.895 819.140 274.825 ;
        RECT 820.100 273.895 820.270 275.005 ;
        RECT 818.810 273.725 820.270 273.895 ;
        RECT 818.810 271.865 819.080 273.725 ;
        RECT 819.940 273.225 820.270 273.725 ;
        RECT 820.450 273.520 820.700 274.825 ;
        RECT 820.940 274.210 821.190 274.825 ;
        RECT 821.370 274.560 821.540 275.005 ;
        RECT 822.230 275.005 823.970 275.175 ;
        RECT 822.230 274.560 822.400 275.005 ;
        RECT 821.370 274.390 822.400 274.560 ;
        RECT 822.580 274.210 822.750 274.825 ;
        RECT 823.280 274.570 823.610 274.825 ;
        RECT 820.940 274.040 822.750 274.210 ;
        RECT 822.930 274.040 823.150 274.370 ;
        RECT 822.580 273.860 822.750 274.040 ;
        RECT 822.580 273.690 822.800 273.860 ;
        RECT 820.450 273.290 820.975 273.520 ;
        RECT 820.450 272.365 820.720 273.290 ;
        RECT 820.390 271.865 820.720 272.365 ;
        RECT 822.115 272.180 822.445 273.475 ;
        RECT 822.630 272.695 822.800 273.690 ;
        RECT 822.980 273.520 823.150 274.040 ;
        RECT 823.330 273.870 823.500 274.570 ;
        RECT 823.800 274.415 823.970 275.005 ;
        RECT 825.280 275.005 826.310 275.175 ;
        RECT 825.280 274.415 825.450 275.005 ;
        RECT 823.800 274.370 825.450 274.415 ;
        RECT 823.680 274.245 825.450 274.370 ;
        RECT 823.680 274.050 824.010 274.245 ;
        RECT 825.630 274.065 825.960 274.825 ;
        RECT 826.140 274.645 826.310 275.005 ;
        RECT 826.140 274.475 827.950 274.645 ;
        RECT 824.190 273.895 825.960 274.065 ;
        RECT 824.190 273.870 824.360 273.895 ;
        RECT 823.330 273.700 824.360 273.870 ;
        RECT 827.270 273.715 827.600 274.295 ;
        RECT 822.980 273.290 824.005 273.520 ;
        RECT 823.675 272.795 824.005 273.290 ;
        RECT 824.190 273.015 824.360 273.700 ;
        RECT 824.540 273.545 827.600 273.715 ;
        RECT 824.540 273.195 824.870 273.545 ;
        RECT 824.190 272.845 826.810 273.015 ;
        RECT 822.630 272.195 822.900 272.695 ;
        RECT 824.190 272.615 824.360 272.845 ;
        RECT 823.350 272.445 824.360 272.615 ;
        RECT 827.340 272.695 827.600 273.545 ;
        RECT 827.780 273.125 827.950 274.475 ;
        RECT 828.130 274.215 828.380 275.125 ;
        RECT 828.130 274.045 829.005 274.215 ;
        RECT 828.325 273.305 828.655 273.805 ;
        RECT 828.835 273.725 829.005 274.045 ;
        RECT 830.540 274.075 830.790 274.545 ;
        RECT 830.540 273.905 831.545 274.075 ;
        RECT 828.835 273.555 831.195 273.725 ;
        RECT 827.780 272.955 828.950 273.125 ;
        RECT 823.350 272.195 823.680 272.445 ;
        RECT 827.340 271.985 827.670 272.695 ;
        RECT 828.130 272.155 828.460 272.695 ;
        RECT 828.665 272.455 828.950 272.955 ;
        RECT 829.130 272.155 829.300 273.555 ;
        RECT 831.375 273.375 831.545 273.905 ;
        RECT 829.505 273.205 831.545 273.375 ;
        RECT 829.505 272.815 829.835 273.205 ;
        RECT 828.130 271.985 829.300 272.155 ;
        RECT 831.320 272.365 831.545 273.205 ;
        RECT 832.045 273.375 832.295 274.375 ;
        RECT 832.045 273.045 833.420 273.375 ;
        RECT 832.045 272.865 832.255 273.045 ;
        RECT 831.925 272.365 832.255 272.865 ;
        RECT 831.320 271.865 831.650 272.365 ;
        RECT 833.600 272.035 833.935 275.105 ;
        RECT 838.550 273.405 838.800 274.455 ;
        RECT 839.250 273.900 839.480 273.910 ;
        RECT 839.025 273.585 839.985 273.900 ;
        RECT 840.190 273.405 840.440 274.455 ;
        RECT 841.785 273.585 842.135 275.165 ;
        RECT 851.930 274.830 852.560 275.360 ;
        RECT 855.010 274.620 855.250 279.030 ;
        RECT 856.645 278.895 856.815 279.805 ;
        RECT 858.375 279.625 858.705 279.805 ;
        RECT 856.060 278.725 856.815 278.895 ;
        RECT 856.060 278.395 856.310 278.725 ;
        RECT 856.995 278.710 857.385 279.625 ;
        RECT 858.910 278.395 859.185 281.655 ;
        RECT 865.220 281.200 865.980 282.160 ;
        RECT 838.550 273.235 841.660 273.405 ;
        RECT 838.550 272.235 838.845 273.235 ;
        RECT 841.330 273.075 841.660 273.235 ;
        RECT 839.025 272.530 839.355 273.055 ;
        RECT 839.020 272.240 839.355 272.530 ;
        RECT 839.025 272.220 839.355 272.240 ;
        RECT 839.535 272.220 840.675 273.055 ;
        RECT 841.830 271.905 842.135 273.585 ;
        RECT 848.700 274.310 855.250 274.620 ;
        RECT 848.700 274.290 855.240 274.310 ;
        RECT 845.870 271.225 846.040 271.825 ;
        RECT 845.385 271.055 847.445 271.225 ;
        RECT 844.780 270.995 845.170 271.030 ;
        RECT 639.560 268.980 640.010 269.080 ;
        RECT 610.120 268.530 610.290 268.950 ;
        RECT 610.910 268.530 611.080 268.950 ;
        RECT 611.700 268.530 611.870 268.950 ;
        RECT 612.490 268.530 612.660 268.950 ;
        RECT 613.280 268.530 613.450 268.950 ;
        RECT 613.950 268.480 614.120 268.900 ;
        RECT 615.530 268.480 615.700 268.900 ;
        RECT 617.110 268.480 617.280 268.900 ;
        RECT 617.710 268.500 617.880 268.920 ;
        RECT 618.500 268.500 618.670 268.920 ;
        RECT 619.290 268.500 619.460 268.920 ;
        RECT 620.080 268.500 620.250 268.920 ;
        RECT 620.870 268.500 621.040 268.920 ;
        RECT 637.200 268.790 640.010 268.980 ;
        RECT 637.200 268.780 637.600 268.790 ;
        RECT 600.670 267.750 600.840 268.170 ;
        RECT 601.460 267.750 601.630 268.170 ;
        RECT 602.250 267.750 602.420 268.170 ;
        RECT 603.040 267.750 603.210 268.170 ;
        RECT 603.830 267.750 604.000 268.170 ;
        RECT 608.240 268.060 608.910 268.370 ;
        RECT 622.830 267.950 623.520 268.500 ;
        RECT 639.560 268.390 640.010 268.790 ;
        RECT 643.620 268.450 644.040 269.130 ;
        RECT 681.120 268.965 681.290 269.565 ;
        RECT 680.635 268.795 682.695 268.965 ;
        RECT 627.450 267.880 627.620 268.300 ;
        RECT 628.240 267.880 628.410 268.300 ;
        RECT 629.030 267.880 629.200 268.300 ;
        RECT 629.820 267.880 629.990 268.300 ;
        RECT 630.610 267.880 630.780 268.300 ;
        RECT 680.045 268.065 680.455 268.735 ;
        RECT 639.300 267.590 639.470 268.010 ;
        RECT 643.350 267.640 643.520 268.060 ;
        RECT 680.635 267.885 680.805 268.795 ;
        RECT 682.365 268.615 682.695 268.795 ;
        RECT 680.050 267.715 680.805 267.885 ;
        RECT 606.370 267.010 606.540 267.430 ;
        RECT 607.160 267.010 607.330 267.430 ;
        RECT 607.950 267.010 608.120 267.430 ;
        RECT 608.740 267.010 608.910 267.430 ;
        RECT 609.530 267.010 609.700 267.430 ;
        RECT 610.120 267.060 610.290 267.480 ;
        RECT 610.910 267.060 611.080 267.480 ;
        RECT 611.700 267.060 611.870 267.480 ;
        RECT 612.490 267.060 612.660 267.480 ;
        RECT 613.280 267.060 613.450 267.480 ;
        RECT 613.950 267.010 614.120 267.430 ;
        RECT 615.530 267.010 615.700 267.430 ;
        RECT 617.110 267.010 617.280 267.430 ;
        RECT 617.710 267.030 617.880 267.450 ;
        RECT 618.500 267.030 618.670 267.450 ;
        RECT 619.290 267.030 619.460 267.450 ;
        RECT 620.080 267.030 620.250 267.450 ;
        RECT 620.870 267.030 621.040 267.450 ;
        RECT 621.460 267.010 621.630 267.430 ;
        RECT 622.250 267.010 622.420 267.430 ;
        RECT 623.040 267.010 623.210 267.430 ;
        RECT 623.830 267.010 624.000 267.430 ;
        RECT 624.620 267.010 624.790 267.430 ;
        RECT 680.050 267.385 680.300 267.715 ;
        RECT 680.985 267.700 681.375 268.615 ;
        RECT 682.900 267.385 683.175 270.645 ;
        RECT 686.780 268.975 686.950 269.575 ;
        RECT 686.295 268.805 688.355 268.975 ;
        RECT 685.705 268.075 686.115 268.745 ;
        RECT 686.295 267.895 686.465 268.805 ;
        RECT 688.025 268.625 688.355 268.805 ;
        RECT 688.560 268.910 688.835 270.655 ;
        RECT 691.330 268.995 691.580 269.595 ;
        RECT 685.710 267.725 686.465 267.895 ;
        RECT 686.645 268.430 687.035 268.625 ;
        RECT 688.560 268.520 688.860 268.910 ;
        RECT 691.330 268.825 693.705 268.995 ;
        RECT 686.645 267.850 687.040 268.430 ;
        RECT 685.710 267.395 685.960 267.725 ;
        RECT 686.645 267.710 687.035 267.850 ;
        RECT 688.560 267.395 688.835 268.520 ;
        RECT 691.535 268.360 691.865 268.645 ;
        RECT 691.530 268.095 691.865 268.360 ;
        RECT 691.530 268.090 691.820 268.095 ;
        RECT 692.110 267.915 692.280 268.825 ;
        RECT 693.375 268.645 693.705 268.825 ;
        RECT 692.460 268.095 692.790 268.645 ;
        RECT 692.110 267.415 692.440 267.915 ;
        RECT 693.910 267.415 694.165 270.675 ;
        RECT 698.350 268.985 698.520 269.585 ;
        RECT 697.865 268.815 699.925 268.985 ;
        RECT 697.865 267.905 698.035 268.815 ;
        RECT 699.595 268.635 699.925 268.815 ;
        RECT 697.280 267.735 698.035 267.905 ;
        RECT 697.280 267.405 697.530 267.735 ;
        RECT 698.215 267.720 698.605 268.635 ;
        RECT 700.130 267.405 700.405 270.665 ;
        RECT 704.010 268.995 704.180 269.595 ;
        RECT 703.525 268.825 705.585 268.995 ;
        RECT 702.935 268.095 703.345 268.765 ;
        RECT 703.525 267.915 703.695 268.825 ;
        RECT 705.255 268.645 705.585 268.825 ;
        RECT 705.790 268.930 706.065 270.675 ;
        RECT 708.560 269.015 708.810 269.615 ;
        RECT 702.940 267.745 703.695 267.915 ;
        RECT 703.875 268.450 704.265 268.645 ;
        RECT 705.790 268.540 706.090 268.930 ;
        RECT 708.560 268.845 710.935 269.015 ;
        RECT 703.875 267.870 704.270 268.450 ;
        RECT 702.940 267.415 703.190 267.745 ;
        RECT 703.875 267.730 704.265 267.870 ;
        RECT 705.790 267.415 706.065 268.540 ;
        RECT 708.765 268.380 709.095 268.665 ;
        RECT 708.760 268.115 709.095 268.380 ;
        RECT 708.760 268.110 709.050 268.115 ;
        RECT 709.340 267.935 709.510 268.845 ;
        RECT 710.605 268.665 710.935 268.845 ;
        RECT 709.690 268.115 710.020 268.665 ;
        RECT 709.340 267.435 709.670 267.935 ;
        RECT 711.140 267.435 711.395 270.695 ;
        RECT 715.920 269.085 716.090 269.685 ;
        RECT 715.435 268.915 717.495 269.085 ;
        RECT 715.435 268.005 715.605 268.915 ;
        RECT 717.165 268.735 717.495 268.915 ;
        RECT 714.850 267.835 715.605 268.005 ;
        RECT 714.850 267.505 715.100 267.835 ;
        RECT 715.785 267.820 716.175 268.735 ;
        RECT 717.700 267.505 717.975 270.765 ;
        RECT 721.580 269.095 721.750 269.695 ;
        RECT 721.095 268.925 723.155 269.095 ;
        RECT 720.505 268.195 720.915 268.865 ;
        RECT 721.095 268.015 721.265 268.925 ;
        RECT 722.825 268.745 723.155 268.925 ;
        RECT 723.360 269.030 723.635 270.775 ;
        RECT 726.130 269.115 726.380 269.715 ;
        RECT 720.510 267.845 721.265 268.015 ;
        RECT 721.445 268.550 721.835 268.745 ;
        RECT 723.360 268.640 723.660 269.030 ;
        RECT 726.130 268.945 728.505 269.115 ;
        RECT 721.445 267.970 721.840 268.550 ;
        RECT 720.510 267.515 720.760 267.845 ;
        RECT 721.445 267.830 721.835 267.970 ;
        RECT 723.360 267.515 723.635 268.640 ;
        RECT 726.335 268.480 726.665 268.765 ;
        RECT 726.330 268.215 726.665 268.480 ;
        RECT 726.330 268.210 726.620 268.215 ;
        RECT 726.910 268.035 727.080 268.945 ;
        RECT 728.175 268.765 728.505 268.945 ;
        RECT 727.260 268.215 727.590 268.765 ;
        RECT 726.910 267.535 727.240 268.035 ;
        RECT 728.710 267.535 728.965 270.795 ;
        RECT 733.090 269.115 733.260 269.715 ;
        RECT 732.605 268.945 734.665 269.115 ;
        RECT 732.605 268.035 732.775 268.945 ;
        RECT 734.335 268.765 734.665 268.945 ;
        RECT 732.020 267.865 732.775 268.035 ;
        RECT 732.020 267.535 732.270 267.865 ;
        RECT 732.955 267.850 733.345 268.765 ;
        RECT 734.870 267.535 735.145 270.795 ;
        RECT 738.750 269.125 738.920 269.725 ;
        RECT 738.265 268.955 740.325 269.125 ;
        RECT 737.675 268.225 738.085 268.895 ;
        RECT 738.265 268.045 738.435 268.955 ;
        RECT 739.995 268.775 740.325 268.955 ;
        RECT 740.530 269.060 740.805 270.805 ;
        RECT 743.300 269.145 743.550 269.745 ;
        RECT 737.680 267.875 738.435 268.045 ;
        RECT 738.615 268.580 739.005 268.775 ;
        RECT 740.530 268.670 740.830 269.060 ;
        RECT 743.300 268.975 745.675 269.145 ;
        RECT 738.615 268.000 739.010 268.580 ;
        RECT 737.680 267.545 737.930 267.875 ;
        RECT 738.615 267.860 739.005 268.000 ;
        RECT 740.530 267.545 740.805 268.670 ;
        RECT 743.505 268.510 743.835 268.795 ;
        RECT 743.500 268.245 743.835 268.510 ;
        RECT 743.500 268.240 743.790 268.245 ;
        RECT 744.080 268.065 744.250 268.975 ;
        RECT 745.345 268.795 745.675 268.975 ;
        RECT 744.430 268.245 744.760 268.795 ;
        RECT 744.080 267.565 744.410 268.065 ;
        RECT 745.880 267.565 746.135 270.825 ;
        RECT 750.900 269.175 751.070 269.775 ;
        RECT 750.415 269.005 752.475 269.175 ;
        RECT 750.415 268.095 750.585 269.005 ;
        RECT 752.145 268.825 752.475 269.005 ;
        RECT 749.830 267.925 750.585 268.095 ;
        RECT 749.830 267.595 750.080 267.925 ;
        RECT 750.765 267.910 751.155 268.825 ;
        RECT 752.680 267.595 752.955 270.855 ;
        RECT 756.560 269.185 756.730 269.785 ;
        RECT 756.075 269.015 758.135 269.185 ;
        RECT 755.485 268.285 755.895 268.955 ;
        RECT 756.075 268.105 756.245 269.015 ;
        RECT 757.805 268.835 758.135 269.015 ;
        RECT 758.340 269.120 758.615 270.865 ;
        RECT 761.110 269.205 761.360 269.805 ;
        RECT 755.490 267.935 756.245 268.105 ;
        RECT 758.340 268.730 758.640 269.120 ;
        RECT 761.110 269.035 763.485 269.205 ;
        RECT 755.490 267.605 755.740 267.935 ;
        RECT 758.340 267.605 758.615 268.730 ;
        RECT 761.315 268.570 761.645 268.855 ;
        RECT 761.310 268.305 761.645 268.570 ;
        RECT 761.310 268.300 761.600 268.305 ;
        RECT 761.890 268.125 762.060 269.035 ;
        RECT 763.155 268.855 763.485 269.035 ;
        RECT 762.240 268.305 762.570 268.855 ;
        RECT 761.890 267.625 762.220 268.125 ;
        RECT 763.690 267.625 763.945 270.885 ;
        RECT 844.780 270.710 845.205 270.995 ;
        RECT 844.795 270.325 845.205 270.710 ;
        RECT 845.385 270.145 845.555 271.055 ;
        RECT 847.115 270.875 847.445 271.055 ;
        RECT 847.650 270.940 847.925 272.905 ;
        RECT 848.700 270.940 849.020 274.290 ;
        RECT 852.000 273.090 852.530 273.750 ;
        RECT 857.130 273.435 857.300 274.035 ;
        RECT 856.645 273.265 858.705 273.435 ;
        RECT 856.055 273.090 856.465 273.205 ;
        RECT 851.040 271.335 851.425 272.915 ;
        RECT 852.000 272.830 856.465 273.090 ;
        RECT 856.055 272.535 856.465 272.830 ;
        RECT 856.645 272.355 856.815 273.265 ;
        RECT 858.375 273.085 858.705 273.265 ;
        RECT 856.060 272.185 856.815 272.355 ;
        RECT 856.060 271.855 856.310 272.185 ;
        RECT 856.995 272.170 857.385 273.085 ;
        RECT 858.910 272.410 859.185 275.115 ;
        RECT 860.210 272.410 860.380 272.420 ;
        RECT 858.910 272.230 860.380 272.410 ;
        RECT 858.910 271.855 859.185 272.230 ;
        RECT 849.330 270.940 849.560 270.950 ;
        RECT 850.205 270.940 850.915 271.095 ;
        RECT 844.800 269.975 845.555 270.145 ;
        RECT 844.800 269.645 845.050 269.975 ;
        RECT 845.735 269.960 846.125 270.875 ;
        RECT 847.650 270.730 850.915 270.940 ;
        RECT 847.650 269.645 847.925 270.730 ;
        RECT 839.630 267.925 839.800 268.525 ;
        RECT 839.145 267.755 841.205 267.925 ;
        RECT 782.370 267.485 783.810 267.655 ;
        RECT 591.660 264.020 592.010 266.180 ;
        RECT 601.360 266.090 602.710 266.600 ;
        RECT 781.080 266.375 781.410 267.305 ;
        RECT 782.370 266.375 782.540 267.485 ;
        RECT 781.080 266.205 782.540 266.375 ;
        RECT 781.080 264.345 781.350 266.205 ;
        RECT 782.210 265.705 782.540 266.205 ;
        RECT 782.720 266.000 782.970 267.305 ;
        RECT 783.210 266.690 783.460 267.305 ;
        RECT 783.640 267.040 783.810 267.485 ;
        RECT 784.500 267.485 786.240 267.655 ;
        RECT 784.500 267.040 784.670 267.485 ;
        RECT 783.640 266.870 784.670 267.040 ;
        RECT 784.850 266.690 785.020 267.305 ;
        RECT 785.550 267.050 785.880 267.305 ;
        RECT 783.210 266.520 785.020 266.690 ;
        RECT 785.200 266.520 785.420 266.850 ;
        RECT 784.850 266.340 785.020 266.520 ;
        RECT 784.850 266.170 785.070 266.340 ;
        RECT 782.720 265.770 783.245 266.000 ;
        RECT 782.720 264.845 782.990 265.770 ;
        RECT 782.660 264.345 782.990 264.845 ;
        RECT 784.385 264.660 784.715 265.955 ;
        RECT 784.900 265.175 785.070 266.170 ;
        RECT 785.250 266.000 785.420 266.520 ;
        RECT 785.600 266.350 785.770 267.050 ;
        RECT 786.070 266.895 786.240 267.485 ;
        RECT 787.550 267.485 788.580 267.655 ;
        RECT 787.550 266.895 787.720 267.485 ;
        RECT 786.070 266.850 787.720 266.895 ;
        RECT 785.950 266.725 787.720 266.850 ;
        RECT 785.950 266.530 786.280 266.725 ;
        RECT 787.900 266.545 788.230 267.305 ;
        RECT 788.410 267.125 788.580 267.485 ;
        RECT 788.410 266.955 790.220 267.125 ;
        RECT 786.460 266.375 788.230 266.545 ;
        RECT 786.460 266.350 786.630 266.375 ;
        RECT 785.600 266.180 786.630 266.350 ;
        RECT 789.540 266.195 789.870 266.775 ;
        RECT 785.250 265.770 786.275 266.000 ;
        RECT 785.945 265.275 786.275 265.770 ;
        RECT 786.460 265.495 786.630 266.180 ;
        RECT 786.810 266.025 789.870 266.195 ;
        RECT 786.810 265.675 787.140 266.025 ;
        RECT 786.460 265.325 789.080 265.495 ;
        RECT 784.900 264.675 785.170 265.175 ;
        RECT 786.460 265.095 786.630 265.325 ;
        RECT 785.620 264.925 786.630 265.095 ;
        RECT 789.610 265.175 789.870 266.025 ;
        RECT 790.050 265.605 790.220 266.955 ;
        RECT 790.400 266.695 790.650 267.605 ;
        RECT 790.400 266.525 791.275 266.695 ;
        RECT 790.595 265.785 790.925 266.285 ;
        RECT 791.105 266.205 791.275 266.525 ;
        RECT 792.810 266.555 793.060 267.025 ;
        RECT 792.810 266.385 793.815 266.555 ;
        RECT 791.105 266.035 793.465 266.205 ;
        RECT 790.050 265.435 791.220 265.605 ;
        RECT 785.620 264.675 785.950 264.925 ;
        RECT 789.610 264.465 789.940 265.175 ;
        RECT 790.400 264.635 790.730 265.175 ;
        RECT 790.935 264.935 791.220 265.435 ;
        RECT 791.400 264.635 791.570 266.035 ;
        RECT 793.645 265.855 793.815 266.385 ;
        RECT 791.775 265.685 793.815 265.855 ;
        RECT 791.775 265.295 792.105 265.685 ;
        RECT 790.400 264.465 791.570 264.635 ;
        RECT 793.590 264.845 793.815 265.685 ;
        RECT 794.315 265.855 794.565 266.855 ;
        RECT 794.315 265.525 795.690 265.855 ;
        RECT 794.315 265.345 794.525 265.525 ;
        RECT 794.195 264.845 794.525 265.345 ;
        RECT 793.590 264.345 793.920 264.845 ;
        RECT 795.870 264.515 796.205 267.585 ;
        RECT 800.900 267.545 802.340 267.715 ;
        RECT 799.610 266.435 799.940 267.365 ;
        RECT 800.900 266.435 801.070 267.545 ;
        RECT 799.610 266.265 801.070 266.435 ;
        RECT 799.610 264.405 799.880 266.265 ;
        RECT 800.740 265.765 801.070 266.265 ;
        RECT 801.250 266.060 801.500 267.365 ;
        RECT 801.740 266.750 801.990 267.365 ;
        RECT 802.170 267.100 802.340 267.545 ;
        RECT 803.030 267.545 804.770 267.715 ;
        RECT 803.030 267.100 803.200 267.545 ;
        RECT 802.170 266.930 803.200 267.100 ;
        RECT 803.380 266.750 803.550 267.365 ;
        RECT 804.080 267.110 804.410 267.365 ;
        RECT 801.740 266.580 803.550 266.750 ;
        RECT 803.730 266.580 803.950 266.910 ;
        RECT 803.380 266.400 803.550 266.580 ;
        RECT 803.380 266.230 803.600 266.400 ;
        RECT 801.250 265.830 801.775 266.060 ;
        RECT 801.250 264.905 801.520 265.830 ;
        RECT 801.190 264.405 801.520 264.905 ;
        RECT 802.915 264.720 803.245 266.015 ;
        RECT 803.430 265.235 803.600 266.230 ;
        RECT 803.780 266.060 803.950 266.580 ;
        RECT 804.130 266.410 804.300 267.110 ;
        RECT 804.600 266.955 804.770 267.545 ;
        RECT 806.080 267.545 807.110 267.715 ;
        RECT 806.080 266.955 806.250 267.545 ;
        RECT 804.600 266.910 806.250 266.955 ;
        RECT 804.480 266.785 806.250 266.910 ;
        RECT 804.480 266.590 804.810 266.785 ;
        RECT 806.430 266.605 806.760 267.365 ;
        RECT 806.940 267.185 807.110 267.545 ;
        RECT 806.940 267.015 808.750 267.185 ;
        RECT 804.990 266.435 806.760 266.605 ;
        RECT 804.990 266.410 805.160 266.435 ;
        RECT 804.130 266.240 805.160 266.410 ;
        RECT 808.070 266.255 808.400 266.835 ;
        RECT 803.780 265.830 804.805 266.060 ;
        RECT 804.475 265.335 804.805 265.830 ;
        RECT 804.990 265.555 805.160 266.240 ;
        RECT 805.340 266.085 808.400 266.255 ;
        RECT 805.340 265.735 805.670 266.085 ;
        RECT 804.990 265.385 807.610 265.555 ;
        RECT 803.430 264.735 803.700 265.235 ;
        RECT 804.990 265.155 805.160 265.385 ;
        RECT 804.150 264.985 805.160 265.155 ;
        RECT 808.140 265.235 808.400 266.085 ;
        RECT 808.580 265.665 808.750 267.015 ;
        RECT 808.930 266.755 809.180 267.665 ;
        RECT 808.930 266.585 809.805 266.755 ;
        RECT 809.125 265.845 809.455 266.345 ;
        RECT 809.635 266.265 809.805 266.585 ;
        RECT 811.340 266.615 811.590 267.085 ;
        RECT 811.340 266.445 812.345 266.615 ;
        RECT 809.635 266.095 811.995 266.265 ;
        RECT 808.580 265.495 809.750 265.665 ;
        RECT 804.150 264.735 804.480 264.985 ;
        RECT 808.140 264.525 808.470 265.235 ;
        RECT 808.930 264.695 809.260 265.235 ;
        RECT 809.465 264.995 809.750 265.495 ;
        RECT 809.930 264.695 810.100 266.095 ;
        RECT 812.175 265.915 812.345 266.445 ;
        RECT 810.305 265.745 812.345 265.915 ;
        RECT 810.305 265.355 810.635 265.745 ;
        RECT 808.930 264.525 810.100 264.695 ;
        RECT 812.120 264.905 812.345 265.745 ;
        RECT 812.845 265.915 813.095 266.915 ;
        RECT 812.845 265.585 814.220 265.915 ;
        RECT 812.845 265.405 813.055 265.585 ;
        RECT 812.725 264.905 813.055 265.405 ;
        RECT 812.120 264.405 812.450 264.905 ;
        RECT 814.400 264.575 814.735 267.645 ;
        RECT 838.555 267.630 838.965 267.695 ;
        RECT 838.530 267.360 838.965 267.630 ;
        RECT 838.555 267.025 838.965 267.360 ;
        RECT 839.145 266.845 839.315 267.755 ;
        RECT 840.875 267.575 841.205 267.755 ;
        RECT 838.560 266.675 839.315 266.845 ;
        RECT 838.560 266.345 838.810 266.675 ;
        RECT 839.495 266.660 839.885 267.575 ;
        RECT 841.410 266.345 841.685 269.605 ;
        RECT 849.330 265.900 849.560 270.730 ;
        RECT 850.205 270.710 850.915 270.730 ;
        RECT 851.095 270.920 851.425 271.335 ;
        RECT 852.460 270.920 852.940 271.090 ;
        RECT 851.095 270.720 852.940 270.920 ;
        RECT 851.095 269.655 851.425 270.720 ;
        RECT 852.460 270.510 852.940 270.720 ;
        RECT 860.210 269.630 860.380 272.230 ;
        RECT 861.650 270.045 861.900 270.645 ;
        RECT 861.650 269.875 864.025 270.045 ;
        RECT 861.855 269.630 862.185 269.695 ;
        RECT 860.210 269.500 862.185 269.630 ;
        RECT 860.220 269.450 862.185 269.500 ;
        RECT 860.220 269.440 860.890 269.450 ;
        RECT 861.855 269.145 862.185 269.450 ;
        RECT 862.430 268.965 862.600 269.875 ;
        RECT 863.695 269.695 864.025 269.875 ;
        RECT 862.780 269.145 863.110 269.695 ;
        RECT 864.230 269.650 864.485 271.725 ;
        RECT 865.380 269.650 866.770 270.030 ;
        RECT 864.230 269.420 866.770 269.650 ;
        RECT 862.430 268.465 862.760 268.965 ;
        RECT 864.230 268.465 864.485 269.420 ;
        RECT 865.380 268.840 866.770 269.420 ;
        RECT 858.990 267.720 859.265 268.445 ;
        RECT 857.210 266.765 857.380 267.365 ;
        RECT 858.980 267.330 859.265 267.720 ;
        RECT 856.725 266.595 858.785 266.765 ;
        RECT 856.135 266.250 856.545 266.535 ;
        RECT 854.710 266.020 856.545 266.250 ;
        RECT 853.610 265.900 854.060 265.960 ;
        RECT 849.330 265.890 854.060 265.900 ;
        RECT 849.310 265.630 854.060 265.890 ;
        RECT 632.160 259.980 633.650 260.970 ;
        RECT 679.500 259.305 679.750 260.455 ;
        RECT 682.080 259.825 682.250 260.455 ;
        RECT 684.270 259.825 684.520 260.455 ;
        RECT 682.080 259.655 684.520 259.825 ;
        RECT 682.080 259.485 682.250 259.655 ;
        RECT 682.430 259.305 684.090 259.475 ;
        RECT 679.500 259.135 682.600 259.305 ;
        RECT 602.990 258.500 603.160 258.920 ;
        RECT 604.570 258.500 604.740 258.920 ;
        RECT 607.510 258.510 607.680 258.930 ;
        RECT 609.090 258.510 609.260 258.930 ;
        RECT 612.030 258.510 612.200 258.930 ;
        RECT 613.610 258.510 613.780 258.930 ;
        RECT 616.460 258.490 616.630 258.910 ;
        RECT 618.040 258.490 618.210 258.910 ;
        RECT 620.840 258.500 621.010 258.920 ;
        RECT 622.420 258.500 622.590 258.920 ;
        RECT 625.160 258.490 625.330 258.910 ;
        RECT 626.740 258.490 626.910 258.910 ;
        RECT 679.500 258.295 679.750 259.135 ;
        RECT 679.930 258.475 680.880 258.755 ;
        RECT 680.710 258.295 680.880 258.475 ;
        RECT 682.785 258.295 683.085 258.535 ;
        RECT 679.500 258.125 680.530 258.295 ;
        RECT 680.710 258.205 683.085 258.295 ;
        RECT 680.710 258.125 682.955 258.205 ;
        RECT 379.060 255.950 379.360 256.940 ;
        RECT 385.680 256.710 386.000 257.150 ;
        RECT 602.990 257.030 603.160 257.450 ;
        RECT 604.570 257.030 604.740 257.450 ;
        RECT 607.510 257.040 607.680 257.460 ;
        RECT 609.090 257.040 609.260 257.460 ;
        RECT 612.030 257.040 612.200 257.460 ;
        RECT 613.610 257.040 613.780 257.460 ;
        RECT 616.460 257.020 616.630 257.440 ;
        RECT 618.040 257.020 618.210 257.440 ;
        RECT 620.840 257.030 621.010 257.450 ;
        RECT 622.420 257.030 622.590 257.450 ;
        RECT 625.160 257.020 625.330 257.440 ;
        RECT 626.740 257.020 626.910 257.440 ;
        RECT 385.700 255.970 386.000 256.710 ;
        RECT 385.700 255.950 386.490 255.970 ;
        RECT 379.060 255.640 386.490 255.950 ;
        RECT 379.060 255.610 379.360 255.640 ;
        RECT 379.670 243.450 381.280 255.640 ;
        RECT 385.700 255.600 386.000 255.640 ;
        RECT 595.035 255.335 595.420 256.915 ;
        RECT 613.080 256.080 613.550 256.460 ;
        RECT 615.920 256.040 616.350 256.360 ;
        RECT 620.330 256.180 620.740 256.610 ;
        RECT 635.790 255.785 636.175 257.365 ;
        RECT 639.980 255.875 640.365 257.455 ;
        RECT 634.955 255.530 635.665 255.545 ;
        RECT 386.610 253.990 388.450 255.270 ;
        RECT 594.040 255.000 594.720 255.090 ;
        RECT 595.035 255.000 595.365 255.335 ;
        RECT 633.810 255.160 635.665 255.530 ;
        RECT 635.845 255.460 636.175 255.785 ;
        RECT 638.970 255.635 639.340 255.660 ;
        RECT 636.600 255.460 637.440 255.470 ;
        RECT 635.845 255.420 637.440 255.460 ;
        RECT 635.845 255.180 637.450 255.420 ;
        RECT 638.970 255.250 639.855 255.635 ;
        RECT 640.035 255.520 640.365 255.875 ;
        RECT 644.080 255.855 644.465 257.435 ;
        RECT 680.280 257.195 680.530 258.125 ;
        RECT 683.335 258.025 683.740 259.125 ;
        RECT 683.920 258.695 684.090 259.305 ;
        RECT 684.270 258.875 684.520 259.655 ;
        RECT 696.780 259.315 697.030 260.465 ;
        RECT 699.360 259.835 699.530 260.465 ;
        RECT 701.550 259.835 701.800 260.465 ;
        RECT 699.360 259.665 701.800 259.835 ;
        RECT 699.360 259.495 699.530 259.665 ;
        RECT 699.710 259.315 701.370 259.485 ;
        RECT 696.780 259.145 699.880 259.315 ;
        RECT 683.920 258.365 684.250 258.695 ;
        RECT 696.780 258.305 697.030 259.145 ;
        RECT 697.210 258.485 698.160 258.765 ;
        RECT 697.990 258.305 698.160 258.485 ;
        RECT 700.065 258.410 700.365 258.545 ;
        RECT 700.065 258.305 700.380 258.410 ;
        RECT 696.780 258.135 697.810 258.305 ;
        RECT 697.990 258.170 700.380 258.305 ;
        RECT 697.990 258.135 700.235 258.170 ;
        RECT 683.220 257.195 683.740 258.025 ;
        RECT 697.560 257.205 697.810 258.135 ;
        RECT 700.615 258.035 701.020 259.135 ;
        RECT 701.200 258.705 701.370 259.315 ;
        RECT 701.550 258.885 701.800 259.665 ;
        RECT 714.550 259.315 714.800 260.465 ;
        RECT 717.130 259.835 717.300 260.465 ;
        RECT 719.320 259.835 719.570 260.465 ;
        RECT 717.130 259.665 719.570 259.835 ;
        RECT 717.130 259.495 717.300 259.665 ;
        RECT 717.480 259.315 719.140 259.485 ;
        RECT 714.550 259.145 717.650 259.315 ;
        RECT 701.200 258.375 701.530 258.705 ;
        RECT 714.550 258.305 714.800 259.145 ;
        RECT 714.980 258.485 715.930 258.765 ;
        RECT 715.760 258.305 715.930 258.485 ;
        RECT 717.835 258.305 718.135 258.545 ;
        RECT 714.550 258.135 715.580 258.305 ;
        RECT 715.760 258.215 718.135 258.305 ;
        RECT 715.760 258.180 718.120 258.215 ;
        RECT 715.760 258.135 718.005 258.180 ;
        RECT 700.500 257.205 701.020 258.035 ;
        RECT 715.330 257.205 715.580 258.135 ;
        RECT 718.385 258.035 718.790 259.135 ;
        RECT 718.970 258.705 719.140 259.315 ;
        RECT 719.320 258.885 719.570 259.665 ;
        RECT 731.790 259.315 732.040 260.465 ;
        RECT 734.370 259.835 734.540 260.465 ;
        RECT 736.560 259.835 736.810 260.465 ;
        RECT 734.370 259.665 736.810 259.835 ;
        RECT 734.370 259.495 734.540 259.665 ;
        RECT 734.720 259.315 736.380 259.485 ;
        RECT 731.790 259.145 734.890 259.315 ;
        RECT 718.970 258.375 719.300 258.705 ;
        RECT 731.790 258.305 732.040 259.145 ;
        RECT 732.220 258.485 733.170 258.765 ;
        RECT 733.000 258.305 733.170 258.485 ;
        RECT 735.075 258.305 735.375 258.545 ;
        RECT 731.790 258.135 732.820 258.305 ;
        RECT 733.000 258.215 735.375 258.305 ;
        RECT 733.000 258.210 735.360 258.215 ;
        RECT 733.000 258.135 735.245 258.210 ;
        RECT 718.270 257.205 718.790 258.035 ;
        RECT 732.570 257.205 732.820 258.135 ;
        RECT 735.625 258.035 736.030 259.135 ;
        RECT 736.210 258.705 736.380 259.315 ;
        RECT 736.560 258.885 736.810 259.665 ;
        RECT 749.270 259.325 749.520 260.475 ;
        RECT 751.850 259.845 752.020 260.475 ;
        RECT 754.040 259.845 754.290 260.475 ;
        RECT 751.850 259.675 754.290 259.845 ;
        RECT 751.850 259.505 752.020 259.675 ;
        RECT 752.200 259.325 753.860 259.495 ;
        RECT 749.270 259.155 752.370 259.325 ;
        RECT 736.210 258.375 736.540 258.705 ;
        RECT 749.270 258.315 749.520 259.155 ;
        RECT 749.700 258.495 750.650 258.775 ;
        RECT 750.480 258.315 750.650 258.495 ;
        RECT 752.555 258.315 752.855 258.555 ;
        RECT 749.270 258.145 750.300 258.315 ;
        RECT 750.480 258.225 752.855 258.315 ;
        RECT 750.480 258.170 752.840 258.225 ;
        RECT 750.480 258.145 752.725 258.170 ;
        RECT 735.510 257.205 736.030 258.035 ;
        RECT 750.050 257.215 750.300 258.145 ;
        RECT 753.105 258.045 753.510 259.145 ;
        RECT 753.690 258.715 753.860 259.325 ;
        RECT 754.040 258.895 754.290 259.675 ;
        RECT 753.690 258.385 754.020 258.715 ;
        RECT 752.990 257.215 753.510 258.045 ;
        RECT 643.245 255.520 643.955 255.615 ;
        RECT 640.035 255.310 643.955 255.520 ;
        RECT 638.970 255.210 639.340 255.250 ;
        RECT 594.040 254.760 595.365 255.000 ;
        RECT 594.040 254.690 594.720 254.760 ;
        RECT 595.035 253.655 595.365 254.760 ;
        RECT 595.545 255.050 596.255 255.095 ;
        RECT 596.720 255.050 597.350 255.160 ;
        RECT 595.545 254.710 597.350 255.050 ;
        RECT 595.990 254.690 597.350 254.710 ;
        RECT 596.720 254.310 597.350 254.690 ;
        RECT 633.810 255.120 635.370 255.160 ;
        RECT 633.810 254.670 634.090 255.120 ;
        RECT 631.290 253.410 631.990 254.040 ;
        RECT 633.590 253.990 634.300 254.670 ;
        RECT 635.845 254.105 636.175 255.180 ;
        RECT 609.970 252.270 610.140 252.690 ;
        RECT 610.760 252.270 610.930 252.690 ;
        RECT 611.550 252.270 611.720 252.690 ;
        RECT 612.340 252.270 612.510 252.690 ;
        RECT 613.130 252.270 613.300 252.690 ;
        RECT 617.560 252.240 617.730 252.660 ;
        RECT 618.350 252.240 618.520 252.660 ;
        RECT 619.140 252.240 619.310 252.660 ;
        RECT 619.930 252.240 620.100 252.660 ;
        RECT 620.720 252.240 620.890 252.660 ;
        RECT 600.520 251.490 600.690 251.910 ;
        RECT 601.310 251.490 601.480 251.910 ;
        RECT 602.100 251.490 602.270 251.910 ;
        RECT 602.890 251.490 603.060 251.910 ;
        RECT 603.680 251.490 603.850 251.910 ;
        RECT 615.080 251.760 615.560 252.180 ;
        RECT 627.300 251.620 627.470 252.040 ;
        RECT 628.090 251.620 628.260 252.040 ;
        RECT 628.880 251.620 629.050 252.040 ;
        RECT 629.670 251.620 629.840 252.040 ;
        RECT 630.460 251.620 630.630 252.040 ;
        RECT 637.050 251.250 637.450 255.180 ;
        RECT 640.035 254.195 640.365 255.310 ;
        RECT 641.520 254.970 641.750 255.310 ;
        RECT 643.245 255.230 643.955 255.310 ;
        RECT 644.135 255.410 644.465 255.855 ;
        RECT 645.030 255.410 645.340 255.430 ;
        RECT 644.135 255.230 645.340 255.410 ;
        RECT 641.450 254.650 641.830 254.970 ;
        RECT 644.135 254.175 644.465 255.230 ;
        RECT 645.030 255.080 645.340 255.230 ;
        RECT 679.910 253.645 680.160 254.795 ;
        RECT 682.490 254.165 682.660 254.795 ;
        RECT 684.680 254.165 684.930 254.795 ;
        RECT 682.490 253.995 684.930 254.165 ;
        RECT 682.490 253.825 682.660 253.995 ;
        RECT 682.840 253.645 684.500 253.815 ;
        RECT 679.910 253.475 683.010 253.645 ;
        RECT 679.910 252.635 680.160 253.475 ;
        RECT 680.340 252.815 681.290 253.095 ;
        RECT 681.120 252.635 681.290 252.815 ;
        RECT 683.195 252.635 683.495 252.875 ;
        RECT 679.910 252.465 680.940 252.635 ;
        RECT 681.120 252.545 683.495 252.635 ;
        RECT 681.120 252.465 683.365 252.545 ;
        RECT 680.690 251.535 680.940 252.465 ;
        RECT 683.745 252.365 684.150 253.465 ;
        RECT 684.330 253.035 684.500 253.645 ;
        RECT 684.680 253.215 684.930 253.995 ;
        RECT 687.150 253.605 687.400 254.755 ;
        RECT 689.730 254.125 689.900 254.755 ;
        RECT 691.920 254.125 692.170 254.755 ;
        RECT 689.730 253.955 692.170 254.125 ;
        RECT 689.730 253.785 689.900 253.955 ;
        RECT 690.080 253.605 691.740 253.775 ;
        RECT 687.150 253.435 690.250 253.605 ;
        RECT 684.330 252.705 684.660 253.035 ;
        RECT 687.150 252.595 687.400 253.435 ;
        RECT 687.580 252.775 688.530 253.055 ;
        RECT 689.065 252.775 690.255 253.150 ;
        RECT 688.360 252.595 688.530 252.775 ;
        RECT 690.435 252.595 690.735 252.835 ;
        RECT 687.150 252.425 688.180 252.595 ;
        RECT 688.360 252.505 690.735 252.595 ;
        RECT 688.360 252.425 690.605 252.505 ;
        RECT 683.630 251.535 684.150 252.365 ;
        RECT 687.930 251.495 688.180 252.425 ;
        RECT 690.985 252.325 691.390 253.425 ;
        RECT 691.570 252.995 691.740 253.605 ;
        RECT 691.920 253.175 692.170 253.955 ;
        RECT 697.140 253.665 697.390 254.815 ;
        RECT 699.720 254.185 699.890 254.815 ;
        RECT 701.910 254.185 702.160 254.815 ;
        RECT 699.720 254.015 702.160 254.185 ;
        RECT 699.720 253.845 699.890 254.015 ;
        RECT 700.070 253.665 701.730 253.835 ;
        RECT 697.140 253.495 700.240 253.665 ;
        RECT 691.570 252.665 691.900 252.995 ;
        RECT 697.140 252.655 697.390 253.495 ;
        RECT 697.570 252.835 698.520 253.115 ;
        RECT 698.350 252.655 698.520 252.835 ;
        RECT 700.425 252.655 700.725 252.895 ;
        RECT 697.140 252.485 698.170 252.655 ;
        RECT 698.350 252.565 700.725 252.655 ;
        RECT 698.350 252.485 700.595 252.565 ;
        RECT 690.870 251.495 691.390 252.325 ;
        RECT 697.920 251.555 698.170 252.485 ;
        RECT 700.975 252.385 701.380 253.485 ;
        RECT 701.560 253.055 701.730 253.665 ;
        RECT 701.910 253.235 702.160 254.015 ;
        RECT 704.380 253.625 704.630 254.775 ;
        RECT 706.960 254.145 707.130 254.775 ;
        RECT 709.150 254.145 709.400 254.775 ;
        RECT 706.960 253.975 709.400 254.145 ;
        RECT 706.960 253.805 707.130 253.975 ;
        RECT 707.310 253.625 708.970 253.795 ;
        RECT 704.380 253.455 707.480 253.625 ;
        RECT 701.560 252.725 701.890 253.055 ;
        RECT 704.380 252.615 704.630 253.455 ;
        RECT 704.810 252.795 705.760 253.075 ;
        RECT 706.295 252.795 707.485 253.170 ;
        RECT 705.590 252.615 705.760 252.795 ;
        RECT 707.665 252.615 707.965 252.855 ;
        RECT 704.380 252.445 705.410 252.615 ;
        RECT 705.590 252.525 707.965 252.615 ;
        RECT 705.590 252.445 707.835 252.525 ;
        RECT 700.860 251.555 701.380 252.385 ;
        RECT 705.160 251.515 705.410 252.445 ;
        RECT 708.215 252.345 708.620 253.445 ;
        RECT 708.800 253.015 708.970 253.625 ;
        RECT 709.150 253.195 709.400 253.975 ;
        RECT 714.710 253.765 714.960 254.915 ;
        RECT 717.290 254.285 717.460 254.915 ;
        RECT 719.480 254.285 719.730 254.915 ;
        RECT 717.290 254.115 719.730 254.285 ;
        RECT 717.290 253.945 717.460 254.115 ;
        RECT 717.640 253.765 719.300 253.935 ;
        RECT 714.710 253.595 717.810 253.765 ;
        RECT 708.800 252.685 709.130 253.015 ;
        RECT 714.710 252.755 714.960 253.595 ;
        RECT 715.140 252.935 716.090 253.215 ;
        RECT 715.920 252.755 716.090 252.935 ;
        RECT 717.995 252.755 718.295 252.995 ;
        RECT 714.710 252.585 715.740 252.755 ;
        RECT 715.920 252.665 718.295 252.755 ;
        RECT 715.920 252.585 718.165 252.665 ;
        RECT 708.100 251.515 708.620 252.345 ;
        RECT 715.490 251.655 715.740 252.585 ;
        RECT 718.545 252.485 718.950 253.585 ;
        RECT 719.130 253.155 719.300 253.765 ;
        RECT 719.480 253.335 719.730 254.115 ;
        RECT 721.950 253.725 722.200 254.875 ;
        RECT 724.530 254.245 724.700 254.875 ;
        RECT 726.720 254.245 726.970 254.875 ;
        RECT 724.530 254.075 726.970 254.245 ;
        RECT 724.530 253.905 724.700 254.075 ;
        RECT 724.880 253.725 726.540 253.895 ;
        RECT 721.950 253.555 725.050 253.725 ;
        RECT 719.130 252.825 719.460 253.155 ;
        RECT 721.950 252.715 722.200 253.555 ;
        RECT 722.380 252.895 723.330 253.175 ;
        RECT 723.865 252.895 725.055 253.270 ;
        RECT 723.160 252.715 723.330 252.895 ;
        RECT 725.235 252.715 725.535 252.955 ;
        RECT 721.950 252.545 722.980 252.715 ;
        RECT 723.160 252.625 725.535 252.715 ;
        RECT 723.160 252.545 725.405 252.625 ;
        RECT 718.430 251.655 718.950 252.485 ;
        RECT 722.730 251.615 722.980 252.545 ;
        RECT 725.785 252.445 726.190 253.545 ;
        RECT 726.370 253.115 726.540 253.725 ;
        RECT 726.720 253.295 726.970 254.075 ;
        RECT 731.880 253.795 732.130 254.945 ;
        RECT 734.460 254.315 734.630 254.945 ;
        RECT 736.650 254.315 736.900 254.945 ;
        RECT 734.460 254.145 736.900 254.315 ;
        RECT 734.460 253.975 734.630 254.145 ;
        RECT 734.810 253.795 736.470 253.965 ;
        RECT 731.880 253.625 734.980 253.795 ;
        RECT 726.370 252.785 726.700 253.115 ;
        RECT 731.880 252.785 732.130 253.625 ;
        RECT 732.310 252.965 733.260 253.245 ;
        RECT 733.090 252.785 733.260 252.965 ;
        RECT 735.165 252.785 735.465 253.025 ;
        RECT 731.880 252.615 732.910 252.785 ;
        RECT 733.090 252.695 735.465 252.785 ;
        RECT 733.090 252.615 735.335 252.695 ;
        RECT 725.670 251.615 726.190 252.445 ;
        RECT 732.660 251.685 732.910 252.615 ;
        RECT 735.715 252.515 736.120 253.615 ;
        RECT 736.300 253.185 736.470 253.795 ;
        RECT 736.650 253.365 736.900 254.145 ;
        RECT 739.120 253.755 739.370 254.905 ;
        RECT 741.700 254.275 741.870 254.905 ;
        RECT 743.890 254.275 744.140 254.905 ;
        RECT 741.700 254.105 744.140 254.275 ;
        RECT 741.700 253.935 741.870 254.105 ;
        RECT 742.050 253.755 743.710 253.925 ;
        RECT 739.120 253.585 742.220 253.755 ;
        RECT 736.300 252.855 736.630 253.185 ;
        RECT 739.120 252.745 739.370 253.585 ;
        RECT 739.550 252.925 740.500 253.205 ;
        RECT 741.035 252.925 742.225 253.300 ;
        RECT 740.330 252.745 740.500 252.925 ;
        RECT 742.405 252.745 742.705 252.985 ;
        RECT 739.120 252.575 740.150 252.745 ;
        RECT 740.330 252.655 742.705 252.745 ;
        RECT 740.330 252.575 742.575 252.655 ;
        RECT 735.600 251.685 736.120 252.515 ;
        RECT 739.900 251.645 740.150 252.575 ;
        RECT 742.955 252.475 743.360 253.575 ;
        RECT 743.540 253.145 743.710 253.755 ;
        RECT 743.890 253.325 744.140 254.105 ;
        RECT 749.690 253.855 749.940 255.005 ;
        RECT 752.270 254.375 752.440 255.005 ;
        RECT 754.460 254.375 754.710 255.005 ;
        RECT 752.270 254.205 754.710 254.375 ;
        RECT 752.270 254.035 752.440 254.205 ;
        RECT 752.620 253.855 754.280 254.025 ;
        RECT 749.690 253.685 752.790 253.855 ;
        RECT 743.540 252.815 743.870 253.145 ;
        RECT 749.690 252.845 749.940 253.685 ;
        RECT 750.120 253.025 751.070 253.305 ;
        RECT 750.900 252.845 751.070 253.025 ;
        RECT 752.975 252.845 753.275 253.085 ;
        RECT 749.690 252.675 750.720 252.845 ;
        RECT 750.900 252.755 753.275 252.845 ;
        RECT 750.900 252.675 753.145 252.755 ;
        RECT 742.840 251.645 743.360 252.475 ;
        RECT 750.470 251.745 750.720 252.675 ;
        RECT 753.525 252.575 753.930 253.675 ;
        RECT 754.110 253.245 754.280 253.855 ;
        RECT 754.460 253.425 754.710 254.205 ;
        RECT 756.930 253.815 757.180 254.965 ;
        RECT 759.510 254.335 759.680 254.965 ;
        RECT 761.700 254.335 761.950 254.965 ;
        RECT 759.510 254.165 761.950 254.335 ;
        RECT 759.510 253.995 759.680 254.165 ;
        RECT 759.860 253.815 761.520 253.985 ;
        RECT 756.930 253.645 760.030 253.815 ;
        RECT 754.110 252.915 754.440 253.245 ;
        RECT 756.930 252.805 757.180 253.645 ;
        RECT 758.845 252.985 760.035 253.360 ;
        RECT 756.930 252.635 757.960 252.805 ;
        RECT 753.410 251.745 753.930 252.575 ;
        RECT 757.710 251.705 757.960 252.635 ;
        RECT 760.765 252.535 761.170 253.635 ;
        RECT 761.350 253.205 761.520 253.815 ;
        RECT 761.700 253.385 761.950 254.165 ;
        RECT 761.350 252.875 761.680 253.205 ;
        RECT 760.650 251.705 761.170 252.535 ;
        RECT 639.410 251.250 639.860 251.350 ;
        RECT 609.970 250.800 610.140 251.220 ;
        RECT 610.760 250.800 610.930 251.220 ;
        RECT 611.550 250.800 611.720 251.220 ;
        RECT 612.340 250.800 612.510 251.220 ;
        RECT 613.130 250.800 613.300 251.220 ;
        RECT 613.800 250.750 613.970 251.170 ;
        RECT 615.380 250.750 615.550 251.170 ;
        RECT 616.960 250.750 617.130 251.170 ;
        RECT 617.560 250.770 617.730 251.190 ;
        RECT 618.350 250.770 618.520 251.190 ;
        RECT 619.140 250.770 619.310 251.190 ;
        RECT 619.930 250.770 620.100 251.190 ;
        RECT 620.720 250.770 620.890 251.190 ;
        RECT 637.050 251.060 639.860 251.250 ;
        RECT 637.050 251.050 637.450 251.060 ;
        RECT 591.430 248.380 591.780 250.540 ;
        RECT 600.520 250.020 600.690 250.440 ;
        RECT 601.310 250.020 601.480 250.440 ;
        RECT 602.100 250.020 602.270 250.440 ;
        RECT 602.890 250.020 603.060 250.440 ;
        RECT 603.680 250.020 603.850 250.440 ;
        RECT 608.090 250.330 608.760 250.640 ;
        RECT 622.680 250.220 623.370 250.770 ;
        RECT 639.410 250.660 639.860 251.060 ;
        RECT 643.470 250.720 643.890 251.400 ;
        RECT 849.310 251.180 849.640 265.630 ;
        RECT 853.610 265.530 854.060 265.630 ;
        RECT 854.710 254.450 855.260 266.020 ;
        RECT 856.135 265.865 856.545 266.020 ;
        RECT 856.725 265.685 856.895 266.595 ;
        RECT 858.455 266.415 858.785 266.595 ;
        RECT 856.140 265.515 856.895 265.685 ;
        RECT 856.140 265.185 856.390 265.515 ;
        RECT 857.075 265.500 857.465 266.415 ;
        RECT 858.990 265.185 859.265 267.330 ;
        RECT 857.080 257.455 857.250 258.055 ;
        RECT 856.595 257.285 858.655 257.455 ;
        RECT 856.005 256.555 856.415 257.225 ;
        RECT 856.595 256.375 856.765 257.285 ;
        RECT 858.325 257.105 858.655 257.285 ;
        RECT 856.010 256.205 856.765 256.375 ;
        RECT 856.010 255.875 856.260 256.205 ;
        RECT 856.945 256.190 857.335 257.105 ;
        RECT 858.860 257.050 859.135 259.135 ;
        RECT 858.850 256.540 859.135 257.050 ;
        RECT 858.860 255.875 859.135 256.540 ;
        RECT 861.590 254.965 861.840 255.565 ;
        RECT 861.590 254.795 863.965 254.965 ;
        RECT 854.630 253.820 855.420 254.450 ;
        RECT 861.795 254.310 862.125 254.615 ;
        RECT 860.410 254.190 862.125 254.310 ;
        RECT 860.400 254.080 862.125 254.190 ;
        RECT 858.920 252.900 859.195 253.365 ;
        RECT 860.400 252.900 860.610 254.080 ;
        RECT 861.795 254.065 862.125 254.080 ;
        RECT 862.370 253.885 862.540 254.795 ;
        RECT 863.635 254.615 863.965 254.795 ;
        RECT 864.170 254.690 864.425 256.645 ;
        RECT 865.550 254.690 866.900 254.760 ;
        RECT 862.720 254.610 863.050 254.615 ;
        RECT 862.720 254.310 863.060 254.610 ;
        RECT 864.160 254.450 866.900 254.690 ;
        RECT 862.720 254.065 863.050 254.310 ;
        RECT 862.370 253.385 862.700 253.885 ;
        RECT 864.170 253.385 864.425 254.450 ;
        RECT 866.540 253.710 866.890 254.450 ;
        RECT 866.340 252.920 867.280 253.710 ;
        RECT 858.920 252.660 860.610 252.900 ;
        RECT 857.140 251.685 857.310 252.285 ;
        RECT 856.655 251.515 858.715 251.685 ;
        RECT 856.065 251.180 856.475 251.455 ;
        RECT 849.300 250.900 856.475 251.180 ;
        RECT 849.310 250.880 849.640 250.900 ;
        RECT 856.065 250.785 856.475 250.900 ;
        RECT 856.655 250.605 856.825 251.515 ;
        RECT 858.385 251.335 858.715 251.515 ;
        RECT 627.300 250.150 627.470 250.570 ;
        RECT 628.090 250.150 628.260 250.570 ;
        RECT 628.880 250.150 629.050 250.570 ;
        RECT 629.670 250.150 629.840 250.570 ;
        RECT 630.460 250.150 630.630 250.570 ;
        RECT 856.070 250.435 856.825 250.605 ;
        RECT 639.150 249.860 639.320 250.280 ;
        RECT 643.200 249.910 643.370 250.330 ;
        RECT 856.070 250.105 856.320 250.435 ;
        RECT 857.005 250.420 857.395 251.335 ;
        RECT 858.920 250.105 859.195 252.660 ;
        RECT 606.220 249.280 606.390 249.700 ;
        RECT 607.010 249.280 607.180 249.700 ;
        RECT 607.800 249.280 607.970 249.700 ;
        RECT 608.590 249.280 608.760 249.700 ;
        RECT 609.380 249.280 609.550 249.700 ;
        RECT 609.970 249.330 610.140 249.750 ;
        RECT 610.760 249.330 610.930 249.750 ;
        RECT 611.550 249.330 611.720 249.750 ;
        RECT 612.340 249.330 612.510 249.750 ;
        RECT 613.130 249.330 613.300 249.750 ;
        RECT 613.800 249.280 613.970 249.700 ;
        RECT 615.380 249.280 615.550 249.700 ;
        RECT 616.960 249.280 617.130 249.700 ;
        RECT 617.560 249.300 617.730 249.720 ;
        RECT 618.350 249.300 618.520 249.720 ;
        RECT 619.140 249.300 619.310 249.720 ;
        RECT 619.930 249.300 620.100 249.720 ;
        RECT 620.720 249.300 620.890 249.720 ;
        RECT 621.310 249.280 621.480 249.700 ;
        RECT 622.100 249.280 622.270 249.700 ;
        RECT 622.890 249.280 623.060 249.700 ;
        RECT 623.680 249.280 623.850 249.700 ;
        RECT 624.470 249.280 624.640 249.700 ;
        RECT 681.100 247.435 681.270 248.035 ;
        RECT 680.615 247.265 682.675 247.435 ;
        RECT 680.615 246.355 680.785 247.265 ;
        RECT 682.345 247.085 682.675 247.265 ;
        RECT 680.030 246.185 680.785 246.355 ;
        RECT 680.030 245.855 680.280 246.185 ;
        RECT 680.965 246.170 681.355 247.085 ;
        RECT 682.880 245.855 683.155 249.115 ;
        RECT 686.760 247.445 686.930 248.045 ;
        RECT 686.275 247.275 688.335 247.445 ;
        RECT 685.685 246.545 686.095 247.215 ;
        RECT 686.275 246.365 686.445 247.275 ;
        RECT 688.005 247.095 688.335 247.275 ;
        RECT 688.540 247.380 688.815 249.125 ;
        RECT 691.310 247.465 691.560 248.065 ;
        RECT 685.690 246.195 686.445 246.365 ;
        RECT 686.625 246.900 687.015 247.095 ;
        RECT 688.540 246.990 688.840 247.380 ;
        RECT 691.310 247.295 693.685 247.465 ;
        RECT 686.625 246.320 687.020 246.900 ;
        RECT 685.690 245.865 685.940 246.195 ;
        RECT 686.625 246.180 687.015 246.320 ;
        RECT 688.540 245.865 688.815 246.990 ;
        RECT 691.515 246.830 691.845 247.115 ;
        RECT 691.510 246.565 691.845 246.830 ;
        RECT 691.510 246.560 691.800 246.565 ;
        RECT 692.090 246.385 692.260 247.295 ;
        RECT 693.355 247.115 693.685 247.295 ;
        RECT 692.440 246.565 692.770 247.115 ;
        RECT 692.090 245.885 692.420 246.385 ;
        RECT 693.890 245.885 694.145 249.145 ;
        RECT 698.330 247.455 698.500 248.055 ;
        RECT 697.845 247.285 699.905 247.455 ;
        RECT 697.845 246.375 698.015 247.285 ;
        RECT 699.575 247.105 699.905 247.285 ;
        RECT 697.260 246.205 698.015 246.375 ;
        RECT 697.260 245.875 697.510 246.205 ;
        RECT 698.195 246.190 698.585 247.105 ;
        RECT 700.110 245.875 700.385 249.135 ;
        RECT 703.990 247.465 704.160 248.065 ;
        RECT 703.505 247.295 705.565 247.465 ;
        RECT 702.915 246.565 703.325 247.235 ;
        RECT 703.505 246.385 703.675 247.295 ;
        RECT 705.235 247.115 705.565 247.295 ;
        RECT 705.770 247.400 706.045 249.145 ;
        RECT 708.540 247.485 708.790 248.085 ;
        RECT 702.920 246.215 703.675 246.385 ;
        RECT 703.855 246.920 704.245 247.115 ;
        RECT 705.770 247.010 706.070 247.400 ;
        RECT 708.540 247.315 710.915 247.485 ;
        RECT 703.855 246.340 704.250 246.920 ;
        RECT 702.920 245.885 703.170 246.215 ;
        RECT 703.855 246.200 704.245 246.340 ;
        RECT 705.770 245.885 706.045 247.010 ;
        RECT 708.745 246.850 709.075 247.135 ;
        RECT 708.740 246.585 709.075 246.850 ;
        RECT 708.740 246.580 709.030 246.585 ;
        RECT 709.320 246.405 709.490 247.315 ;
        RECT 710.585 247.135 710.915 247.315 ;
        RECT 709.670 246.585 710.000 247.135 ;
        RECT 709.320 245.905 709.650 246.405 ;
        RECT 711.120 245.905 711.375 249.165 ;
        RECT 715.900 247.555 716.070 248.155 ;
        RECT 715.415 247.385 717.475 247.555 ;
        RECT 715.415 246.475 715.585 247.385 ;
        RECT 717.145 247.205 717.475 247.385 ;
        RECT 714.830 246.305 715.585 246.475 ;
        RECT 714.830 245.975 715.080 246.305 ;
        RECT 715.765 246.290 716.155 247.205 ;
        RECT 717.680 245.975 717.955 249.235 ;
        RECT 721.560 247.565 721.730 248.165 ;
        RECT 721.075 247.395 723.135 247.565 ;
        RECT 720.485 246.665 720.895 247.335 ;
        RECT 721.075 246.485 721.245 247.395 ;
        RECT 722.805 247.215 723.135 247.395 ;
        RECT 723.340 247.500 723.615 249.245 ;
        RECT 726.110 247.585 726.360 248.185 ;
        RECT 720.490 246.315 721.245 246.485 ;
        RECT 721.425 247.020 721.815 247.215 ;
        RECT 723.340 247.110 723.640 247.500 ;
        RECT 726.110 247.415 728.485 247.585 ;
        RECT 721.425 246.440 721.820 247.020 ;
        RECT 720.490 245.985 720.740 246.315 ;
        RECT 721.425 246.300 721.815 246.440 ;
        RECT 723.340 245.985 723.615 247.110 ;
        RECT 726.315 246.950 726.645 247.235 ;
        RECT 726.310 246.685 726.645 246.950 ;
        RECT 726.310 246.680 726.600 246.685 ;
        RECT 726.890 246.505 727.060 247.415 ;
        RECT 728.155 247.235 728.485 247.415 ;
        RECT 727.240 246.685 727.570 247.235 ;
        RECT 726.890 246.005 727.220 246.505 ;
        RECT 728.690 246.005 728.945 249.265 ;
        RECT 733.070 247.585 733.240 248.185 ;
        RECT 732.585 247.415 734.645 247.585 ;
        RECT 732.585 246.505 732.755 247.415 ;
        RECT 734.315 247.235 734.645 247.415 ;
        RECT 732.000 246.335 732.755 246.505 ;
        RECT 732.000 246.005 732.250 246.335 ;
        RECT 732.935 246.320 733.325 247.235 ;
        RECT 734.850 246.005 735.125 249.265 ;
        RECT 738.730 247.595 738.900 248.195 ;
        RECT 738.245 247.425 740.305 247.595 ;
        RECT 737.655 246.695 738.065 247.365 ;
        RECT 738.245 246.515 738.415 247.425 ;
        RECT 739.975 247.245 740.305 247.425 ;
        RECT 740.510 247.530 740.785 249.275 ;
        RECT 743.280 247.615 743.530 248.215 ;
        RECT 737.660 246.345 738.415 246.515 ;
        RECT 738.595 247.050 738.985 247.245 ;
        RECT 740.510 247.140 740.810 247.530 ;
        RECT 743.280 247.445 745.655 247.615 ;
        RECT 738.595 246.470 738.990 247.050 ;
        RECT 737.660 246.015 737.910 246.345 ;
        RECT 738.595 246.330 738.985 246.470 ;
        RECT 740.510 246.015 740.785 247.140 ;
        RECT 743.485 246.980 743.815 247.265 ;
        RECT 743.480 246.715 743.815 246.980 ;
        RECT 743.480 246.710 743.770 246.715 ;
        RECT 744.060 246.535 744.230 247.445 ;
        RECT 745.325 247.265 745.655 247.445 ;
        RECT 744.410 246.715 744.740 247.265 ;
        RECT 744.060 246.035 744.390 246.535 ;
        RECT 745.860 246.035 746.115 249.295 ;
        RECT 750.880 247.645 751.050 248.245 ;
        RECT 750.395 247.475 752.455 247.645 ;
        RECT 750.395 246.565 750.565 247.475 ;
        RECT 752.125 247.295 752.455 247.475 ;
        RECT 749.810 246.395 750.565 246.565 ;
        RECT 749.810 246.065 750.060 246.395 ;
        RECT 750.745 246.380 751.135 247.295 ;
        RECT 752.660 246.065 752.935 249.325 ;
        RECT 756.540 247.655 756.710 248.255 ;
        RECT 756.055 247.485 758.115 247.655 ;
        RECT 755.465 246.755 755.875 247.425 ;
        RECT 756.055 246.575 756.225 247.485 ;
        RECT 757.785 247.305 758.115 247.485 ;
        RECT 758.320 247.590 758.595 249.335 ;
        RECT 761.090 247.675 761.340 248.275 ;
        RECT 755.470 246.405 756.225 246.575 ;
        RECT 758.320 247.200 758.620 247.590 ;
        RECT 761.090 247.505 763.465 247.675 ;
        RECT 755.470 246.075 755.720 246.405 ;
        RECT 758.320 246.075 758.595 247.200 ;
        RECT 761.295 247.040 761.625 247.325 ;
        RECT 761.290 246.775 761.625 247.040 ;
        RECT 761.290 246.770 761.580 246.775 ;
        RECT 761.870 246.595 762.040 247.505 ;
        RECT 763.135 247.325 763.465 247.505 ;
        RECT 762.220 246.775 762.550 247.325 ;
        RECT 761.870 246.095 762.200 246.595 ;
        RECT 763.670 246.095 763.925 249.355 ;
        RECT 378.670 241.130 381.980 243.450 ;
        RECT 330.920 232.520 333.480 232.620 ;
        RECT 294.690 231.710 333.480 232.520 ;
        RECT 330.920 231.240 333.480 231.710 ;
        RECT 331.210 217.660 332.110 231.240 ;
        RECT 338.660 218.070 340.190 218.140 ;
        RECT 331.210 217.130 332.240 217.660 ;
        RECT 331.340 216.350 332.240 217.130 ;
        RECT 338.660 216.980 341.140 218.070 ;
        RECT 338.050 216.370 338.360 216.390 ;
        RECT 338.010 216.350 338.360 216.370 ;
        RECT 344.520 216.350 344.990 216.370 ;
        RECT 331.340 215.970 344.990 216.350 ;
        RECT 331.340 215.730 332.240 215.970 ;
        RECT 331.360 214.830 331.770 215.730 ;
        RECT 331.460 201.340 331.750 214.830 ;
        RECT 338.010 214.770 338.360 215.970 ;
        RECT 338.010 201.360 338.300 214.770 ;
        RECT 344.520 214.460 344.990 215.970 ;
        RECT 344.590 201.380 344.880 214.460 ;
        RECT 331.510 200.730 331.680 201.340 ;
        RECT 338.090 200.730 338.260 201.360 ;
        RECT 344.670 200.730 344.840 201.380 ;
        RECT 402.070 196.240 402.840 196.960 ;
        RECT 404.230 196.950 405.700 197.910 ;
        RECT 409.010 196.240 409.320 196.290 ;
        RECT 415.510 196.240 415.820 196.390 ;
        RECT 402.070 195.970 415.930 196.240 ;
        RECT 402.070 195.770 402.840 195.970 ;
        RECT 402.350 195.230 402.660 195.770 ;
        RECT 402.350 195.000 402.680 195.230 ;
        RECT 409.010 195.120 409.320 195.970 ;
        RECT 415.510 195.400 415.820 195.970 ;
        RECT 402.430 177.590 402.660 195.000 ;
        RECT 409.020 177.670 409.250 195.120 ;
        RECT 415.510 195.040 415.850 195.400 ;
        RECT 415.620 177.750 415.850 195.040 ;
        RECT 402.480 177.150 402.650 177.590 ;
        RECT 409.060 177.150 409.230 177.670 ;
        RECT 415.640 177.150 415.810 177.750 ;
      LAYER mcon ;
        RECT 379.300 369.765 379.470 369.935 ;
        RECT 379.300 369.405 379.470 369.575 ;
        RECT 385.880 369.765 386.050 369.935 ;
        RECT 385.880 369.405 386.050 369.575 ;
        RECT 379.160 365.195 379.330 365.365 ;
        RECT 379.160 364.835 379.330 365.005 ;
        RECT 379.160 361.725 379.330 361.895 ;
        RECT 379.160 361.365 379.330 361.535 ;
        RECT 379.160 358.255 379.330 358.425 ;
        RECT 379.160 357.895 379.330 358.065 ;
        RECT 379.160 354.785 379.330 354.955 ;
        RECT 379.160 354.425 379.330 354.595 ;
        RECT 379.160 351.315 379.330 351.485 ;
        RECT 385.740 365.195 385.910 365.365 ;
        RECT 385.740 364.835 385.910 365.005 ;
        RECT 385.740 361.725 385.910 361.895 ;
        RECT 385.740 361.365 385.910 361.535 ;
        RECT 385.740 358.255 385.910 358.425 ;
        RECT 385.740 357.895 385.910 358.065 ;
        RECT 385.740 354.785 385.910 354.955 ;
        RECT 385.740 354.425 385.910 354.595 ;
        RECT 653.075 352.535 653.245 352.705 ;
        RECT 653.075 352.175 653.245 352.345 ;
        RECT 385.740 351.315 385.910 351.485 ;
        RECT 379.160 350.955 379.330 351.125 ;
        RECT 385.740 350.955 385.910 351.125 ;
        RECT 662.985 352.800 663.155 352.970 ;
        RECT 668.265 352.800 668.435 352.970 ;
        RECT 670.665 352.800 670.835 352.970 ;
        RECT 669.230 351.885 669.400 352.055 ;
        RECT 672.105 352.585 672.275 352.755 ;
        RECT 675.810 351.805 675.980 351.975 ;
        RECT 681.035 352.760 681.205 352.930 ;
        RECT 686.315 352.760 686.485 352.930 ;
        RECT 688.715 352.760 688.885 352.930 ;
        RECT 687.330 351.885 687.500 352.055 ;
        RECT 690.160 352.530 690.330 352.700 ;
        RECT 693.420 351.885 693.590 352.055 ;
        RECT 698.625 352.780 698.795 352.950 ;
        RECT 703.905 352.780 704.075 352.950 ;
        RECT 706.305 352.780 706.475 352.950 ;
        RECT 704.875 351.915 705.045 352.085 ;
        RECT 707.775 352.650 707.945 352.820 ;
        RECT 711.235 351.845 711.405 352.015 ;
        RECT 716.475 352.780 716.645 352.950 ;
        RECT 721.755 352.780 721.925 352.950 ;
        RECT 724.155 352.780 724.325 352.950 ;
        RECT 722.755 351.835 722.925 352.005 ;
        RECT 725.595 352.550 725.765 352.720 ;
        RECT 729.505 351.815 729.675 351.985 ;
        RECT 734.735 352.780 734.905 352.950 ;
        RECT 740.015 352.780 740.185 352.950 ;
        RECT 742.415 352.780 742.585 352.950 ;
        RECT 741.000 351.905 741.170 352.075 ;
        RECT 743.865 352.605 744.035 352.775 ;
        RECT 747.270 351.815 747.440 351.985 ;
        RECT 752.505 352.750 752.675 352.920 ;
        RECT 757.785 352.750 757.955 352.920 ;
        RECT 760.185 352.750 760.355 352.920 ;
        RECT 758.770 351.640 758.940 351.810 ;
        RECT 761.625 352.605 761.795 352.775 ;
        RECT 765.300 351.695 765.470 351.865 ;
        RECT 770.545 352.670 770.715 352.840 ;
        RECT 775.825 352.670 775.995 352.840 ;
        RECT 778.225 352.670 778.395 352.840 ;
        RECT 776.795 351.805 776.965 351.975 ;
        RECT 779.640 352.530 779.810 352.700 ;
        RECT 783.475 351.685 783.645 351.855 ;
        RECT 788.705 352.710 788.875 352.880 ;
        RECT 793.985 352.710 794.155 352.880 ;
        RECT 796.385 352.710 796.555 352.880 ;
        RECT 794.945 351.695 795.115 351.865 ;
        RECT 797.805 352.590 797.975 352.760 ;
        RECT 801.855 351.705 802.025 351.875 ;
        RECT 807.085 352.720 807.255 352.890 ;
        RECT 812.365 352.720 812.535 352.890 ;
        RECT 814.765 352.720 814.935 352.890 ;
        RECT 813.345 351.740 813.515 351.910 ;
        RECT 816.185 352.615 816.355 352.785 ;
        RECT 818.590 351.710 819.480 352.240 ;
        RECT 656.110 349.645 656.640 350.175 ;
        RECT 820.665 351.660 820.835 351.830 ;
        RECT 825.885 352.700 826.055 352.870 ;
        RECT 829.060 351.780 829.230 351.950 ;
        RECT 831.165 352.700 831.335 352.870 ;
        RECT 833.565 352.700 833.735 352.870 ;
        RECT 835.005 352.625 835.175 352.795 ;
        RECT 839.120 353.320 839.290 353.490 ;
        RECT 836.175 351.315 836.705 351.845 ;
        RECT 832.135 348.125 834.105 349.375 ;
        RECT 837.460 347.340 838.710 348.230 ;
        RECT 379.140 346.315 379.310 346.485 ;
        RECT 379.140 345.955 379.310 346.125 ;
        RECT 379.140 342.845 379.310 343.015 ;
        RECT 379.140 342.485 379.310 342.655 ;
        RECT 379.140 339.375 379.310 339.545 ;
        RECT 379.140 339.015 379.310 339.185 ;
        RECT 379.140 335.905 379.310 336.075 ;
        RECT 379.140 335.545 379.310 335.715 ;
        RECT 379.140 332.435 379.310 332.605 ;
        RECT 385.720 346.315 385.890 346.485 ;
        RECT 385.720 345.955 385.890 346.125 ;
        RECT 780.295 343.435 780.825 344.685 ;
        RECT 785.840 343.705 786.010 343.875 ;
        RECT 799.285 344.630 799.455 344.800 ;
        RECT 804.565 344.630 804.735 344.800 ;
        RECT 806.965 344.630 807.135 344.800 ;
        RECT 805.525 343.810 805.695 343.980 ;
        RECT 813.415 345.295 813.585 345.465 ;
        RECT 813.435 343.700 813.605 343.870 ;
        RECT 818.645 344.540 818.815 344.710 ;
        RECT 823.925 344.540 824.095 344.710 ;
        RECT 826.325 344.540 826.495 344.710 ;
        RECT 824.910 343.660 825.080 343.830 ;
        RECT 870.645 345.835 871.895 347.805 ;
        RECT 385.720 342.845 385.890 343.015 ;
        RECT 385.720 342.485 385.890 342.655 ;
        RECT 385.720 339.375 385.890 339.545 ;
        RECT 385.720 339.015 385.890 339.185 ;
        RECT 385.720 335.905 385.890 336.075 ;
        RECT 385.720 335.545 385.890 335.715 ;
        RECT 632.285 333.710 633.175 334.240 ;
        RECT 853.655 338.820 853.825 338.990 ;
        RECT 854.015 338.820 854.185 338.990 ;
        RECT 852.620 337.645 852.790 337.815 ;
        RECT 855.200 337.645 855.370 337.815 ;
        RECT 852.620 336.175 852.790 336.345 ;
        RECT 855.200 336.175 855.370 336.345 ;
        RECT 852.620 334.705 852.790 334.875 ;
        RECT 855.200 334.705 855.370 334.875 ;
        RECT 852.620 333.235 852.790 333.405 ;
        RECT 855.200 333.235 855.370 333.405 ;
        RECT 385.720 332.435 385.890 332.605 ;
        RECT 379.140 332.075 379.310 332.245 ;
        RECT 385.720 332.075 385.890 332.245 ;
        RECT 603.420 332.175 603.590 332.345 ;
        RECT 605.000 332.175 605.170 332.345 ;
        RECT 607.940 332.185 608.110 332.355 ;
        RECT 609.520 332.185 609.690 332.355 ;
        RECT 612.460 332.185 612.630 332.355 ;
        RECT 614.040 332.185 614.210 332.355 ;
        RECT 616.890 332.165 617.060 332.335 ;
        RECT 618.470 332.165 618.640 332.335 ;
        RECT 621.270 332.175 621.440 332.345 ;
        RECT 622.850 332.175 623.020 332.345 ;
        RECT 625.590 332.165 625.760 332.335 ;
        RECT 627.170 332.165 627.340 332.335 ;
        RECT 603.420 330.705 603.590 330.875 ;
        RECT 605.000 330.705 605.170 330.875 ;
        RECT 607.940 330.715 608.110 330.885 ;
        RECT 609.520 330.715 609.690 330.885 ;
        RECT 612.460 330.715 612.630 330.885 ;
        RECT 614.040 330.715 614.210 330.885 ;
        RECT 616.890 330.695 617.060 330.865 ;
        RECT 618.470 330.695 618.640 330.865 ;
        RECT 621.270 330.705 621.440 330.875 ;
        RECT 622.850 330.705 623.020 330.875 ;
        RECT 625.590 330.695 625.760 330.865 ;
        RECT 627.170 330.695 627.340 330.865 ;
        RECT 613.650 329.765 613.820 329.935 ;
        RECT 616.480 329.680 616.650 329.850 ;
        RECT 620.865 329.845 621.035 330.015 ;
        RECT 639.500 328.900 639.670 329.070 ;
        RECT 666.255 330.920 666.425 331.090 ;
        RECT 663.415 329.835 663.585 330.005 ;
        RECT 594.545 328.355 594.715 328.525 ;
        RECT 594.905 328.355 595.075 328.525 ;
        RECT 379.140 327.465 379.310 327.635 ;
        RECT 379.140 327.105 379.310 327.275 ;
        RECT 379.140 323.995 379.310 324.165 ;
        RECT 379.140 323.635 379.310 323.805 ;
        RECT 209.210 320.835 210.100 321.365 ;
        RECT 379.140 320.525 379.310 320.695 ;
        RECT 379.140 320.165 379.310 320.335 ;
        RECT 212.115 319.320 212.285 319.490 ;
        RECT 212.475 319.320 212.645 319.490 ;
        RECT 215.585 319.320 215.755 319.490 ;
        RECT 215.945 319.320 216.115 319.490 ;
        RECT 219.055 319.320 219.225 319.490 ;
        RECT 219.415 319.320 219.585 319.490 ;
        RECT 222.525 319.320 222.695 319.490 ;
        RECT 222.885 319.320 223.055 319.490 ;
        RECT 225.995 319.320 226.165 319.490 ;
        RECT 226.355 319.320 226.525 319.490 ;
        RECT 232.155 319.310 232.325 319.480 ;
        RECT 232.515 319.310 232.685 319.480 ;
        RECT 235.625 319.310 235.795 319.480 ;
        RECT 235.985 319.310 236.155 319.480 ;
        RECT 239.095 319.310 239.265 319.480 ;
        RECT 239.455 319.310 239.625 319.480 ;
        RECT 242.565 319.310 242.735 319.480 ;
        RECT 242.925 319.310 243.095 319.480 ;
        RECT 246.035 319.310 246.205 319.480 ;
        RECT 246.395 319.310 246.565 319.480 ;
        RECT 252.215 319.310 252.385 319.480 ;
        RECT 252.575 319.310 252.745 319.480 ;
        RECT 255.685 319.310 255.855 319.480 ;
        RECT 256.045 319.310 256.215 319.480 ;
        RECT 259.155 319.310 259.325 319.480 ;
        RECT 259.515 319.310 259.685 319.480 ;
        RECT 262.625 319.310 262.795 319.480 ;
        RECT 262.985 319.310 263.155 319.480 ;
        RECT 266.095 319.310 266.265 319.480 ;
        RECT 266.455 319.310 266.625 319.480 ;
        RECT 272.265 319.310 272.435 319.480 ;
        RECT 272.625 319.310 272.795 319.480 ;
        RECT 275.735 319.310 275.905 319.480 ;
        RECT 276.095 319.310 276.265 319.480 ;
        RECT 279.205 319.310 279.375 319.480 ;
        RECT 279.565 319.310 279.735 319.480 ;
        RECT 282.675 319.310 282.845 319.480 ;
        RECT 283.035 319.310 283.205 319.480 ;
        RECT 286.145 319.310 286.315 319.480 ;
        RECT 286.505 319.310 286.675 319.480 ;
        RECT 379.140 317.055 379.310 317.225 ;
        RECT 379.140 316.695 379.310 316.865 ;
        RECT 379.140 313.585 379.310 313.755 ;
        RECT 385.720 327.465 385.890 327.635 ;
        RECT 385.720 327.105 385.890 327.275 ;
        RECT 597.200 328.020 597.730 328.550 ;
        RECT 634.110 327.615 634.640 328.145 ;
        RECT 631.760 327.175 631.930 327.345 ;
        RECT 632.120 327.175 632.290 327.345 ;
        RECT 610.400 325.945 610.570 326.115 ;
        RECT 611.190 325.945 611.360 326.115 ;
        RECT 611.980 325.945 612.150 326.115 ;
        RECT 612.770 325.945 612.940 326.115 ;
        RECT 613.560 325.945 613.730 326.115 ;
        RECT 617.990 325.915 618.160 326.085 ;
        RECT 618.780 325.915 618.950 326.085 ;
        RECT 619.570 325.915 619.740 326.085 ;
        RECT 620.360 325.915 620.530 326.085 ;
        RECT 621.150 325.915 621.320 326.085 ;
        RECT 600.950 325.165 601.120 325.335 ;
        RECT 601.740 325.165 601.910 325.335 ;
        RECT 602.530 325.165 602.700 325.335 ;
        RECT 603.320 325.165 603.490 325.335 ;
        RECT 604.110 325.165 604.280 325.335 ;
        RECT 615.640 325.425 615.810 325.595 ;
        RECT 627.730 325.295 627.900 325.465 ;
        RECT 628.520 325.295 628.690 325.465 ;
        RECT 629.310 325.295 629.480 325.465 ;
        RECT 630.100 325.295 630.270 325.465 ;
        RECT 630.890 325.295 631.060 325.465 ;
        RECT 664.370 329.525 664.540 329.695 ;
        RECT 668.965 329.840 669.135 330.010 ;
        RECT 669.985 329.580 670.155 329.750 ;
        RECT 682.430 330.680 682.600 330.850 ;
        RECT 677.635 330.150 677.805 330.320 ;
        RECT 676.185 329.840 676.355 330.010 ;
        RECT 682.310 329.660 682.480 329.830 ;
        RECT 683.255 329.460 683.425 329.630 ;
        RECT 688.630 329.815 688.800 329.985 ;
        RECT 641.985 328.275 642.155 328.445 ;
        RECT 645.530 328.720 645.700 328.890 ;
        RECT 610.400 324.475 610.570 324.645 ;
        RECT 611.190 324.475 611.360 324.645 ;
        RECT 611.980 324.475 612.150 324.645 ;
        RECT 612.770 324.475 612.940 324.645 ;
        RECT 613.560 324.475 613.730 324.645 ;
        RECT 614.230 324.425 614.400 324.595 ;
        RECT 615.810 324.425 615.980 324.595 ;
        RECT 617.390 324.425 617.560 324.595 ;
        RECT 617.990 324.445 618.160 324.615 ;
        RECT 618.780 324.445 618.950 324.615 ;
        RECT 619.570 324.445 619.740 324.615 ;
        RECT 620.360 324.445 620.530 324.615 ;
        RECT 621.150 324.445 621.320 324.615 ;
        RECT 639.975 324.505 640.145 324.675 ;
        RECT 385.720 323.995 385.890 324.165 ;
        RECT 385.720 323.635 385.890 323.805 ;
        RECT 600.950 323.695 601.120 323.865 ;
        RECT 601.740 323.695 601.910 323.865 ;
        RECT 602.530 323.695 602.700 323.865 ;
        RECT 603.320 323.695 603.490 323.865 ;
        RECT 608.770 323.965 608.940 324.135 ;
        RECT 644.010 324.555 644.180 324.725 ;
        RECT 623.370 323.960 623.540 324.130 ;
        RECT 604.110 323.695 604.280 323.865 ;
        RECT 627.730 323.825 627.900 323.995 ;
        RECT 628.520 323.825 628.690 323.995 ;
        RECT 629.310 323.825 629.480 323.995 ;
        RECT 630.100 323.825 630.270 323.995 ;
        RECT 630.890 323.825 631.060 323.995 ;
        RECT 639.580 323.535 639.750 323.705 ;
        RECT 643.630 323.585 643.800 323.755 ;
        RECT 657.710 323.660 658.240 324.190 ;
        RECT 606.650 322.955 606.820 323.125 ;
        RECT 607.440 322.955 607.610 323.125 ;
        RECT 608.230 322.955 608.400 323.125 ;
        RECT 609.020 322.955 609.190 323.125 ;
        RECT 609.810 322.955 609.980 323.125 ;
        RECT 610.400 323.005 610.570 323.175 ;
        RECT 611.190 323.005 611.360 323.175 ;
        RECT 611.980 323.005 612.150 323.175 ;
        RECT 612.770 323.005 612.940 323.175 ;
        RECT 613.560 323.005 613.730 323.175 ;
        RECT 614.230 322.955 614.400 323.125 ;
        RECT 615.810 322.955 615.980 323.125 ;
        RECT 617.390 322.955 617.560 323.125 ;
        RECT 617.990 322.975 618.160 323.145 ;
        RECT 618.780 322.975 618.950 323.145 ;
        RECT 619.570 322.975 619.740 323.145 ;
        RECT 620.360 322.975 620.530 323.145 ;
        RECT 621.150 322.975 621.320 323.145 ;
        RECT 621.740 322.955 621.910 323.125 ;
        RECT 622.530 322.955 622.700 323.125 ;
        RECT 623.320 322.955 623.490 323.125 ;
        RECT 624.110 322.955 624.280 323.125 ;
        RECT 624.900 322.955 625.070 323.125 ;
        RECT 660.330 323.540 660.860 324.070 ;
        RECT 662.495 323.635 663.025 324.165 ;
        RECT 665.665 323.845 665.835 324.015 ;
        RECT 667.245 323.870 667.415 324.040 ;
        RECT 667.605 323.870 667.775 324.040 ;
        RECT 665.665 323.485 665.835 323.655 ;
        RECT 669.360 323.505 669.530 323.675 ;
        RECT 670.015 323.655 670.545 324.185 ;
        RECT 671.850 323.935 672.020 324.105 ;
        RECT 671.850 323.575 672.020 323.745 ;
        RECT 677.440 324.435 677.610 324.605 ;
        RECT 679.685 324.800 679.855 324.970 ;
        RECT 673.850 323.430 674.020 323.600 ;
        RECT 676.890 323.575 677.060 323.745 ;
        RECT 678.210 323.065 678.380 323.235 ;
        RECT 682.230 323.620 682.400 323.790 ;
        RECT 683.175 323.200 683.345 323.370 ;
        RECT 688.640 323.155 688.810 323.325 ;
        RECT 385.720 320.525 385.890 320.695 ;
        RECT 385.720 320.165 385.890 320.335 ;
        RECT 591.920 322.205 592.090 322.375 ;
        RECT 591.920 321.845 592.090 322.015 ;
        RECT 602.540 321.980 602.710 322.150 ;
        RECT 591.920 321.485 592.090 321.655 ;
        RECT 591.920 321.125 592.090 321.295 ;
        RECT 591.920 320.765 592.090 320.935 ;
        RECT 591.920 320.405 592.090 320.575 ;
        RECT 385.720 317.055 385.890 317.225 ;
        RECT 662.140 318.565 662.310 318.735 ;
        RECT 664.850 318.850 665.020 319.020 ;
        RECT 670.255 319.115 670.425 319.285 ;
        RECT 662.070 317.705 662.240 317.875 ;
        RECT 663.010 317.205 663.180 317.375 ;
        RECT 385.720 316.695 385.890 316.865 ;
        RECT 667.445 318.140 667.615 318.310 ;
        RECT 632.700 315.605 633.230 316.135 ;
        RECT 603.270 314.005 603.440 314.175 ;
        RECT 604.850 314.005 605.020 314.175 ;
        RECT 607.790 314.015 607.960 314.185 ;
        RECT 609.370 314.015 609.540 314.185 ;
        RECT 612.310 314.015 612.480 314.185 ;
        RECT 613.890 314.015 614.060 314.185 ;
        RECT 616.740 313.995 616.910 314.165 ;
        RECT 618.320 313.995 618.490 314.165 ;
        RECT 621.120 314.005 621.290 314.175 ;
        RECT 622.700 314.005 622.870 314.175 ;
        RECT 625.440 313.995 625.610 314.165 ;
        RECT 627.020 313.995 627.190 314.165 ;
        RECT 385.720 313.585 385.890 313.755 ;
        RECT 379.140 313.225 379.310 313.395 ;
        RECT 212.115 312.740 212.285 312.910 ;
        RECT 212.475 312.740 212.645 312.910 ;
        RECT 215.585 312.740 215.755 312.910 ;
        RECT 215.945 312.740 216.115 312.910 ;
        RECT 219.055 312.740 219.225 312.910 ;
        RECT 219.415 312.740 219.585 312.910 ;
        RECT 222.525 312.740 222.695 312.910 ;
        RECT 222.885 312.740 223.055 312.910 ;
        RECT 225.995 312.740 226.165 312.910 ;
        RECT 226.355 312.740 226.525 312.910 ;
        RECT 232.155 312.730 232.325 312.900 ;
        RECT 232.515 312.730 232.685 312.900 ;
        RECT 235.625 312.730 235.795 312.900 ;
        RECT 235.985 312.730 236.155 312.900 ;
        RECT 239.095 312.730 239.265 312.900 ;
        RECT 239.455 312.730 239.625 312.900 ;
        RECT 242.565 312.730 242.735 312.900 ;
        RECT 242.925 312.730 243.095 312.900 ;
        RECT 246.035 312.730 246.205 312.900 ;
        RECT 246.395 312.730 246.565 312.900 ;
        RECT 252.215 312.730 252.385 312.900 ;
        RECT 252.575 312.730 252.745 312.900 ;
        RECT 255.685 312.730 255.855 312.900 ;
        RECT 256.045 312.730 256.215 312.900 ;
        RECT 259.155 312.730 259.325 312.900 ;
        RECT 259.515 312.730 259.685 312.900 ;
        RECT 262.625 312.730 262.795 312.900 ;
        RECT 262.985 312.730 263.155 312.900 ;
        RECT 266.095 312.730 266.265 312.900 ;
        RECT 266.455 312.730 266.625 312.900 ;
        RECT 272.265 312.730 272.435 312.900 ;
        RECT 272.625 312.730 272.795 312.900 ;
        RECT 275.735 312.730 275.905 312.900 ;
        RECT 276.095 312.730 276.265 312.900 ;
        RECT 279.205 312.730 279.375 312.900 ;
        RECT 279.565 312.730 279.735 312.900 ;
        RECT 282.675 312.730 282.845 312.900 ;
        RECT 283.035 312.730 283.205 312.900 ;
        RECT 286.145 312.730 286.315 312.900 ;
        RECT 286.505 312.730 286.675 312.900 ;
        RECT 385.720 313.225 385.890 313.395 ;
        RECT 668.380 317.660 668.550 317.830 ;
        RECT 672.875 318.100 673.045 318.270 ;
        RECT 673.815 317.720 673.985 317.890 ;
        RECT 679.585 317.820 679.755 317.990 ;
        RECT 684.485 317.315 684.655 317.485 ;
        RECT 691.930 317.940 692.100 318.110 ;
        RECT 694.220 318.015 694.390 318.185 ;
        RECT 603.270 312.535 603.440 312.705 ;
        RECT 604.850 312.535 605.020 312.705 ;
        RECT 607.790 312.545 607.960 312.715 ;
        RECT 609.370 312.545 609.540 312.715 ;
        RECT 612.310 312.545 612.480 312.715 ;
        RECT 613.890 312.545 614.060 312.715 ;
        RECT 616.740 312.525 616.910 312.695 ;
        RECT 618.320 312.525 618.490 312.695 ;
        RECT 621.120 312.535 621.290 312.705 ;
        RECT 622.700 312.535 622.870 312.705 ;
        RECT 625.440 312.525 625.610 312.695 ;
        RECT 627.020 312.525 627.190 312.695 ;
        RECT 613.500 311.595 613.670 311.765 ;
        RECT 616.330 311.510 616.500 311.680 ;
        RECT 620.715 311.675 620.885 311.845 ;
        RECT 639.350 310.730 639.520 310.900 ;
        RECT 594.395 310.185 594.565 310.355 ;
        RECT 594.755 310.185 594.925 310.355 ;
        RECT 379.140 308.645 379.310 308.815 ;
        RECT 597.050 309.850 597.580 310.380 ;
        RECT 633.960 309.445 634.490 309.975 ;
        RECT 379.140 308.285 379.310 308.455 ;
        RECT 212.115 306.160 212.285 306.330 ;
        RECT 212.475 306.160 212.645 306.330 ;
        RECT 215.585 306.160 215.755 306.330 ;
        RECT 215.945 306.160 216.115 306.330 ;
        RECT 219.055 306.160 219.225 306.330 ;
        RECT 219.415 306.160 219.585 306.330 ;
        RECT 222.525 306.160 222.695 306.330 ;
        RECT 222.885 306.160 223.055 306.330 ;
        RECT 225.995 306.160 226.165 306.330 ;
        RECT 226.355 306.160 226.525 306.330 ;
        RECT 232.155 306.150 232.325 306.320 ;
        RECT 232.515 306.150 232.685 306.320 ;
        RECT 235.625 306.150 235.795 306.320 ;
        RECT 235.985 306.150 236.155 306.320 ;
        RECT 239.095 306.150 239.265 306.320 ;
        RECT 239.455 306.150 239.625 306.320 ;
        RECT 242.565 306.150 242.735 306.320 ;
        RECT 242.925 306.150 243.095 306.320 ;
        RECT 246.035 306.150 246.205 306.320 ;
        RECT 246.395 306.150 246.565 306.320 ;
        RECT 252.215 306.150 252.385 306.320 ;
        RECT 252.575 306.150 252.745 306.320 ;
        RECT 255.685 306.150 255.855 306.320 ;
        RECT 256.045 306.150 256.215 306.320 ;
        RECT 259.155 306.150 259.325 306.320 ;
        RECT 259.515 306.150 259.685 306.320 ;
        RECT 262.625 306.150 262.795 306.320 ;
        RECT 262.985 306.150 263.155 306.320 ;
        RECT 266.095 306.150 266.265 306.320 ;
        RECT 266.455 306.150 266.625 306.320 ;
        RECT 272.265 306.150 272.435 306.320 ;
        RECT 272.625 306.150 272.795 306.320 ;
        RECT 275.735 306.150 275.905 306.320 ;
        RECT 276.095 306.150 276.265 306.320 ;
        RECT 279.205 306.150 279.375 306.320 ;
        RECT 279.565 306.150 279.735 306.320 ;
        RECT 282.675 306.150 282.845 306.320 ;
        RECT 283.035 306.150 283.205 306.320 ;
        RECT 286.145 306.150 286.315 306.320 ;
        RECT 286.505 306.150 286.675 306.320 ;
        RECT 289.080 303.030 289.610 305.360 ;
        RECT 379.140 305.175 379.310 305.345 ;
        RECT 379.140 304.815 379.310 304.985 ;
        RECT 379.140 301.705 379.310 301.875 ;
        RECT 379.140 301.345 379.310 301.515 ;
        RECT 212.075 298.330 212.245 298.500 ;
        RECT 212.435 298.330 212.605 298.500 ;
        RECT 215.545 298.330 215.715 298.500 ;
        RECT 215.905 298.330 216.075 298.500 ;
        RECT 219.015 298.330 219.185 298.500 ;
        RECT 219.375 298.330 219.545 298.500 ;
        RECT 222.485 298.330 222.655 298.500 ;
        RECT 222.845 298.330 223.015 298.500 ;
        RECT 225.955 298.330 226.125 298.500 ;
        RECT 226.315 298.330 226.485 298.500 ;
        RECT 232.045 298.330 232.215 298.500 ;
        RECT 232.405 298.330 232.575 298.500 ;
        RECT 235.515 298.330 235.685 298.500 ;
        RECT 235.875 298.330 236.045 298.500 ;
        RECT 238.985 298.330 239.155 298.500 ;
        RECT 239.345 298.330 239.515 298.500 ;
        RECT 242.455 298.330 242.625 298.500 ;
        RECT 242.815 298.330 242.985 298.500 ;
        RECT 245.925 298.330 246.095 298.500 ;
        RECT 246.285 298.330 246.455 298.500 ;
        RECT 252.155 298.330 252.325 298.500 ;
        RECT 252.515 298.330 252.685 298.500 ;
        RECT 255.625 298.330 255.795 298.500 ;
        RECT 255.985 298.330 256.155 298.500 ;
        RECT 259.095 298.330 259.265 298.500 ;
        RECT 259.455 298.330 259.625 298.500 ;
        RECT 262.565 298.330 262.735 298.500 ;
        RECT 262.925 298.330 263.095 298.500 ;
        RECT 266.035 298.330 266.205 298.500 ;
        RECT 266.395 298.330 266.565 298.500 ;
        RECT 272.265 298.330 272.435 298.500 ;
        RECT 272.625 298.330 272.795 298.500 ;
        RECT 275.735 298.330 275.905 298.500 ;
        RECT 276.095 298.330 276.265 298.500 ;
        RECT 279.205 298.330 279.375 298.500 ;
        RECT 279.565 298.330 279.735 298.500 ;
        RECT 282.675 298.330 282.845 298.500 ;
        RECT 283.035 298.330 283.205 298.500 ;
        RECT 286.145 298.330 286.315 298.500 ;
        RECT 286.505 298.330 286.675 298.500 ;
        RECT 97.885 296.590 98.055 296.760 ;
        RECT 98.245 296.590 98.415 296.760 ;
        RECT 101.355 296.590 101.525 296.760 ;
        RECT 101.715 296.590 101.885 296.760 ;
        RECT 4.855 296.340 5.025 296.510 ;
        RECT 5.215 296.340 5.385 296.510 ;
        RECT 8.325 296.340 8.495 296.510 ;
        RECT 8.685 296.340 8.855 296.510 ;
        RECT 11.795 296.340 11.965 296.510 ;
        RECT 12.155 296.340 12.325 296.510 ;
        RECT 18.195 296.320 18.365 296.490 ;
        RECT 18.555 296.320 18.725 296.490 ;
        RECT 21.665 296.320 21.835 296.490 ;
        RECT 22.025 296.320 22.195 296.490 ;
        RECT 25.135 296.320 25.305 296.490 ;
        RECT 25.495 296.320 25.665 296.490 ;
        RECT 31.565 296.350 31.735 296.520 ;
        RECT 31.925 296.350 32.095 296.520 ;
        RECT 35.035 296.350 35.205 296.520 ;
        RECT 35.395 296.350 35.565 296.520 ;
        RECT 38.505 296.350 38.675 296.520 ;
        RECT 38.865 296.350 39.035 296.520 ;
        RECT 44.795 296.350 44.965 296.520 ;
        RECT 45.155 296.350 45.325 296.520 ;
        RECT 48.265 296.350 48.435 296.520 ;
        RECT 48.625 296.350 48.795 296.520 ;
        RECT 51.735 296.350 51.905 296.520 ;
        RECT 52.095 296.350 52.265 296.520 ;
        RECT 58.065 296.320 58.235 296.490 ;
        RECT 58.425 296.320 58.595 296.490 ;
        RECT 61.535 296.320 61.705 296.490 ;
        RECT 61.895 296.320 62.065 296.490 ;
        RECT 65.005 296.320 65.175 296.490 ;
        RECT 65.365 296.320 65.535 296.490 ;
        RECT 71.335 296.350 71.505 296.520 ;
        RECT 71.695 296.350 71.865 296.520 ;
        RECT 74.805 296.350 74.975 296.520 ;
        RECT 75.165 296.350 75.335 296.520 ;
        RECT 78.275 296.350 78.445 296.520 ;
        RECT 78.635 296.350 78.805 296.520 ;
        RECT 84.465 296.370 84.635 296.540 ;
        RECT 84.825 296.370 84.995 296.540 ;
        RECT 87.935 296.370 88.105 296.540 ;
        RECT 88.295 296.370 88.465 296.540 ;
        RECT 91.405 296.370 91.575 296.540 ;
        RECT 91.765 296.370 91.935 296.540 ;
        RECT 4.855 289.760 5.025 289.930 ;
        RECT 5.215 289.760 5.385 289.930 ;
        RECT 8.325 289.760 8.495 289.930 ;
        RECT 8.685 289.760 8.855 289.930 ;
        RECT 11.795 289.760 11.965 289.930 ;
        RECT 12.155 289.760 12.325 289.930 ;
        RECT 379.140 298.235 379.310 298.405 ;
        RECT 379.140 297.875 379.310 298.045 ;
        RECT 379.140 294.765 379.310 294.935 ;
        RECT 385.720 308.645 385.890 308.815 ;
        RECT 631.810 308.750 632.340 309.280 ;
        RECT 385.720 308.285 385.890 308.455 ;
        RECT 610.250 307.775 610.420 307.945 ;
        RECT 611.040 307.775 611.210 307.945 ;
        RECT 611.830 307.775 612.000 307.945 ;
        RECT 612.620 307.775 612.790 307.945 ;
        RECT 613.410 307.775 613.580 307.945 ;
        RECT 617.840 307.745 618.010 307.915 ;
        RECT 618.630 307.745 618.800 307.915 ;
        RECT 619.420 307.745 619.590 307.915 ;
        RECT 620.210 307.745 620.380 307.915 ;
        RECT 621.000 307.745 621.170 307.915 ;
        RECT 600.800 306.995 600.970 307.165 ;
        RECT 601.590 306.995 601.760 307.165 ;
        RECT 602.380 306.995 602.550 307.165 ;
        RECT 603.170 306.995 603.340 307.165 ;
        RECT 603.960 306.995 604.130 307.165 ;
        RECT 615.490 307.255 615.660 307.425 ;
        RECT 627.580 307.125 627.750 307.295 ;
        RECT 628.370 307.125 628.540 307.295 ;
        RECT 629.160 307.125 629.330 307.295 ;
        RECT 629.950 307.125 630.120 307.295 ;
        RECT 630.740 307.125 630.910 307.295 ;
        RECT 641.835 310.105 642.005 310.275 ;
        RECT 645.380 310.550 645.550 310.720 ;
        RECT 666.260 307.930 667.510 309.180 ;
        RECT 385.720 305.175 385.890 305.345 ;
        RECT 385.720 304.815 385.890 304.985 ;
        RECT 591.940 306.100 592.110 306.270 ;
        RECT 610.250 306.305 610.420 306.475 ;
        RECT 611.040 306.305 611.210 306.475 ;
        RECT 611.830 306.305 612.000 306.475 ;
        RECT 612.620 306.305 612.790 306.475 ;
        RECT 613.410 306.305 613.580 306.475 ;
        RECT 614.080 306.255 614.250 306.425 ;
        RECT 615.660 306.255 615.830 306.425 ;
        RECT 617.240 306.255 617.410 306.425 ;
        RECT 617.840 306.275 618.010 306.445 ;
        RECT 618.630 306.275 618.800 306.445 ;
        RECT 619.420 306.275 619.590 306.445 ;
        RECT 620.210 306.275 620.380 306.445 ;
        RECT 621.000 306.275 621.170 306.445 ;
        RECT 639.825 306.335 639.995 306.505 ;
        RECT 591.940 305.740 592.110 305.910 ;
        RECT 591.940 305.380 592.110 305.550 ;
        RECT 600.800 305.525 600.970 305.695 ;
        RECT 601.590 305.525 601.760 305.695 ;
        RECT 602.380 305.525 602.550 305.695 ;
        RECT 603.170 305.525 603.340 305.695 ;
        RECT 608.620 305.795 608.790 305.965 ;
        RECT 643.860 306.385 644.030 306.555 ;
        RECT 623.220 305.790 623.390 305.960 ;
        RECT 603.960 305.525 604.130 305.695 ;
        RECT 627.580 305.655 627.750 305.825 ;
        RECT 628.370 305.655 628.540 305.825 ;
        RECT 629.160 305.655 629.330 305.825 ;
        RECT 629.950 305.655 630.120 305.825 ;
        RECT 630.740 305.655 630.910 305.825 ;
        RECT 639.430 305.365 639.600 305.535 ;
        RECT 643.480 305.415 643.650 305.585 ;
        RECT 591.940 305.020 592.110 305.190 ;
        RECT 591.940 304.660 592.110 304.830 ;
        RECT 606.500 304.785 606.670 304.955 ;
        RECT 607.290 304.785 607.460 304.955 ;
        RECT 608.080 304.785 608.250 304.955 ;
        RECT 608.870 304.785 609.040 304.955 ;
        RECT 609.660 304.785 609.830 304.955 ;
        RECT 610.250 304.835 610.420 305.005 ;
        RECT 611.040 304.835 611.210 305.005 ;
        RECT 611.830 304.835 612.000 305.005 ;
        RECT 612.620 304.835 612.790 305.005 ;
        RECT 613.410 304.835 613.580 305.005 ;
        RECT 614.080 304.785 614.250 304.955 ;
        RECT 615.660 304.785 615.830 304.955 ;
        RECT 617.240 304.785 617.410 304.955 ;
        RECT 617.840 304.805 618.010 304.975 ;
        RECT 618.630 304.805 618.800 304.975 ;
        RECT 619.420 304.805 619.590 304.975 ;
        RECT 620.210 304.805 620.380 304.975 ;
        RECT 621.000 304.805 621.170 304.975 ;
        RECT 621.590 304.785 621.760 304.955 ;
        RECT 622.380 304.785 622.550 304.955 ;
        RECT 623.170 304.785 623.340 304.955 ;
        RECT 623.960 304.785 624.130 304.955 ;
        RECT 624.750 304.785 624.920 304.955 ;
        RECT 591.940 304.300 592.110 304.470 ;
        RECT 602.170 303.900 602.340 304.070 ;
        RECT 602.530 303.900 602.700 304.070 ;
        RECT 385.720 301.705 385.890 301.875 ;
        RECT 385.720 301.345 385.890 301.515 ;
        RECT 591.940 302.945 592.110 303.115 ;
        RECT 591.940 302.585 592.110 302.755 ;
        RECT 591.940 302.225 592.110 302.395 ;
        RECT 798.555 305.980 798.725 306.150 ;
        RECT 797.120 305.340 797.290 305.510 ;
        RECT 799.965 305.000 800.135 305.170 ;
        RECT 800.955 305.980 801.125 306.150 ;
        RECT 806.235 305.980 806.405 306.150 ;
        RECT 811.500 306.715 811.670 306.885 ;
        RECT 811.505 305.660 811.675 305.830 ;
        RECT 814.900 306.015 815.070 306.185 ;
        RECT 816.315 305.980 816.485 306.150 ;
        RECT 817.725 305.470 817.895 305.640 ;
        RECT 818.715 305.980 818.885 306.150 ;
        RECT 823.995 305.980 824.165 306.150 ;
        RECT 834.200 306.715 834.370 306.885 ;
        RECT 829.215 305.875 829.385 306.045 ;
        RECT 834.270 305.495 834.440 305.665 ;
        RECT 837.595 305.935 837.765 306.105 ;
        RECT 838.930 305.640 839.100 305.810 ;
        RECT 839.485 305.525 839.655 305.695 ;
        RECT 842.915 305.695 843.085 305.865 ;
        RECT 852.620 331.765 852.790 331.935 ;
        RECT 855.200 331.765 855.370 331.935 ;
        RECT 870.830 331.345 871.720 331.875 ;
        RECT 865.720 330.770 865.890 330.940 ;
        RECT 866.080 330.770 866.250 330.940 ;
        RECT 866.440 330.770 866.610 330.940 ;
        RECT 852.620 330.295 852.790 330.465 ;
        RECT 855.200 330.295 855.370 330.465 ;
        RECT 869.930 330.125 870.100 330.295 ;
        RECT 871.220 330.125 871.390 330.295 ;
        RECT 872.510 330.125 872.680 330.295 ;
        RECT 864.740 329.575 864.910 329.745 ;
        RECT 866.030 329.575 866.200 329.745 ;
        RECT 867.320 329.575 867.490 329.745 ;
        RECT 852.620 328.825 852.790 328.995 ;
        RECT 855.200 328.825 855.370 328.995 ;
        RECT 869.930 328.655 870.100 328.825 ;
        RECT 871.220 328.655 871.390 328.825 ;
        RECT 872.510 328.655 872.680 328.825 ;
        RECT 864.740 328.105 864.910 328.275 ;
        RECT 866.030 328.105 866.200 328.275 ;
        RECT 867.320 328.105 867.490 328.275 ;
        RECT 852.620 327.355 852.790 327.525 ;
        RECT 855.200 327.355 855.370 327.525 ;
        RECT 859.460 327.545 859.630 327.715 ;
        RECT 862.040 327.545 862.210 327.715 ;
        RECT 869.930 327.185 870.100 327.355 ;
        RECT 871.220 327.185 871.390 327.355 ;
        RECT 872.510 327.185 872.680 327.355 ;
        RECT 864.740 326.635 864.910 326.805 ;
        RECT 866.030 326.635 866.200 326.805 ;
        RECT 867.320 326.635 867.490 326.805 ;
        RECT 852.620 325.885 852.790 326.055 ;
        RECT 855.200 325.885 855.370 326.055 ;
        RECT 859.460 326.075 859.630 326.245 ;
        RECT 862.040 326.075 862.210 326.245 ;
        RECT 869.930 325.715 870.100 325.885 ;
        RECT 871.220 325.715 871.390 325.885 ;
        RECT 872.510 325.715 872.680 325.885 ;
        RECT 864.740 325.165 864.910 325.335 ;
        RECT 866.030 325.165 866.200 325.335 ;
        RECT 867.320 325.165 867.490 325.335 ;
        RECT 852.620 324.415 852.790 324.585 ;
        RECT 855.200 324.415 855.370 324.585 ;
        RECT 859.460 324.605 859.630 324.775 ;
        RECT 862.040 324.605 862.210 324.775 ;
        RECT 869.930 324.245 870.100 324.415 ;
        RECT 871.220 324.245 871.390 324.415 ;
        RECT 872.510 324.245 872.680 324.415 ;
        RECT 864.740 323.695 864.910 323.865 ;
        RECT 866.030 323.695 866.200 323.865 ;
        RECT 867.320 323.695 867.490 323.865 ;
        RECT 852.620 322.945 852.790 323.115 ;
        RECT 855.200 322.945 855.370 323.115 ;
        RECT 859.460 323.135 859.630 323.305 ;
        RECT 862.040 323.135 862.210 323.305 ;
        RECT 852.620 321.475 852.790 321.645 ;
        RECT 855.200 321.475 855.370 321.645 ;
        RECT 859.460 321.665 859.630 321.835 ;
        RECT 862.040 321.665 862.210 321.835 ;
        RECT 874.400 321.615 874.570 321.785 ;
        RECT 869.970 320.565 870.140 320.735 ;
        RECT 852.620 320.005 852.790 320.175 ;
        RECT 855.200 320.005 855.370 320.175 ;
        RECT 859.460 320.195 859.630 320.365 ;
        RECT 873.220 320.505 873.390 320.675 ;
        RECT 875.800 320.505 875.970 320.675 ;
        RECT 862.040 320.195 862.210 320.365 ;
        RECT 869.970 319.095 870.140 319.265 ;
        RECT 852.620 318.535 852.790 318.705 ;
        RECT 855.200 318.535 855.370 318.705 ;
        RECT 859.460 318.725 859.630 318.895 ;
        RECT 873.220 319.035 873.390 319.205 ;
        RECT 875.800 319.035 875.970 319.205 ;
        RECT 862.040 318.725 862.210 318.895 ;
        RECT 869.970 317.625 870.140 317.795 ;
        RECT 852.620 317.065 852.790 317.235 ;
        RECT 855.200 317.065 855.370 317.235 ;
        RECT 859.460 317.255 859.630 317.425 ;
        RECT 873.220 317.565 873.390 317.735 ;
        RECT 875.800 317.565 875.970 317.735 ;
        RECT 862.040 317.255 862.210 317.425 ;
        RECT 869.970 316.155 870.140 316.325 ;
        RECT 852.620 315.595 852.790 315.765 ;
        RECT 855.200 315.595 855.370 315.765 ;
        RECT 859.460 315.785 859.630 315.955 ;
        RECT 873.220 316.095 873.390 316.265 ;
        RECT 875.800 316.095 875.970 316.265 ;
        RECT 862.040 315.785 862.210 315.955 ;
        RECT 869.970 314.685 870.140 314.855 ;
        RECT 852.620 314.125 852.790 314.295 ;
        RECT 855.200 314.125 855.370 314.295 ;
        RECT 859.460 314.315 859.630 314.485 ;
        RECT 873.220 314.625 873.390 314.795 ;
        RECT 875.800 314.625 875.970 314.795 ;
        RECT 862.040 314.315 862.210 314.485 ;
        RECT 832.870 305.005 833.040 305.175 ;
        RECT 591.940 301.865 592.110 302.035 ;
        RECT 591.940 301.505 592.110 301.675 ;
        RECT 591.940 301.145 592.110 301.315 ;
        RECT 696.505 300.900 697.395 302.150 ;
        RECT 385.720 298.235 385.890 298.405 ;
        RECT 385.720 297.875 385.890 298.045 ;
        RECT 632.585 296.300 633.475 296.830 ;
        RECT 682.135 296.920 682.305 297.090 ;
        RECT 680.700 296.405 680.870 296.575 ;
        RECT 683.555 295.830 683.725 296.000 ;
        RECT 684.535 296.920 684.705 297.090 ;
        RECT 689.815 296.920 689.985 297.090 ;
        RECT 695.065 297.135 695.235 297.305 ;
        RECT 699.625 296.880 699.795 297.050 ;
        RECT 698.230 296.355 698.400 296.525 ;
        RECT 701.035 295.880 701.205 296.050 ;
        RECT 702.025 296.880 702.195 297.050 ;
        RECT 707.305 296.880 707.475 297.050 ;
        RECT 712.550 297.500 712.720 297.670 ;
        RECT 712.550 297.140 712.720 297.310 ;
        RECT 717.235 296.940 717.405 297.110 ;
        RECT 715.800 296.405 715.970 296.575 ;
        RECT 719.635 296.940 719.805 297.110 ;
        RECT 724.915 296.940 725.085 297.110 ;
        RECT 730.140 297.470 730.310 297.640 ;
        RECT 730.140 297.110 730.310 297.280 ;
        RECT 734.935 296.890 735.105 297.060 ;
        RECT 733.520 296.375 733.690 296.545 ;
        RECT 737.335 296.890 737.505 297.060 ;
        RECT 742.615 296.890 742.785 297.060 ;
        RECT 747.855 297.575 748.025 297.745 ;
        RECT 747.855 297.215 748.025 297.385 ;
        RECT 752.675 296.880 752.845 297.050 ;
        RECT 751.250 296.355 751.420 296.525 ;
        RECT 755.075 296.880 755.245 297.050 ;
        RECT 760.355 296.880 760.525 297.050 ;
        RECT 765.585 297.505 765.755 297.675 ;
        RECT 765.585 297.145 765.755 297.315 ;
        RECT 385.720 294.765 385.890 294.935 ;
        RECT 379.140 294.405 379.310 294.575 ;
        RECT 603.220 294.825 603.390 294.995 ;
        RECT 604.800 294.825 604.970 294.995 ;
        RECT 607.740 294.835 607.910 295.005 ;
        RECT 609.320 294.835 609.490 295.005 ;
        RECT 612.260 294.835 612.430 295.005 ;
        RECT 613.840 294.835 614.010 295.005 ;
        RECT 616.690 294.815 616.860 294.985 ;
        RECT 618.270 294.815 618.440 294.985 ;
        RECT 621.070 294.825 621.240 294.995 ;
        RECT 622.650 294.825 622.820 294.995 ;
        RECT 625.390 294.815 625.560 294.985 ;
        RECT 626.970 294.815 627.140 294.985 ;
        RECT 385.720 294.405 385.890 294.575 ;
        RECT 856.050 295.565 856.220 295.735 ;
        RECT 856.990 295.210 857.160 295.380 ;
        RECT 858.845 295.545 859.015 295.715 ;
        RECT 603.220 293.355 603.390 293.525 ;
        RECT 604.800 293.355 604.970 293.525 ;
        RECT 607.740 293.365 607.910 293.535 ;
        RECT 609.320 293.365 609.490 293.535 ;
        RECT 612.260 293.365 612.430 293.535 ;
        RECT 613.840 293.365 614.010 293.535 ;
        RECT 616.690 293.345 616.860 293.515 ;
        RECT 618.270 293.345 618.440 293.515 ;
        RECT 621.070 293.355 621.240 293.525 ;
        RECT 622.650 293.355 622.820 293.525 ;
        RECT 625.390 293.345 625.560 293.515 ;
        RECT 626.970 293.345 627.140 293.515 ;
        RECT 212.075 291.750 212.245 291.920 ;
        RECT 212.435 291.750 212.605 291.920 ;
        RECT 215.545 291.750 215.715 291.920 ;
        RECT 215.905 291.750 216.075 291.920 ;
        RECT 219.015 291.750 219.185 291.920 ;
        RECT 219.375 291.750 219.545 291.920 ;
        RECT 222.485 291.750 222.655 291.920 ;
        RECT 222.845 291.750 223.015 291.920 ;
        RECT 225.955 291.750 226.125 291.920 ;
        RECT 226.315 291.750 226.485 291.920 ;
        RECT 232.045 291.750 232.215 291.920 ;
        RECT 232.405 291.750 232.575 291.920 ;
        RECT 235.515 291.750 235.685 291.920 ;
        RECT 235.875 291.750 236.045 291.920 ;
        RECT 238.985 291.750 239.155 291.920 ;
        RECT 239.345 291.750 239.515 291.920 ;
        RECT 242.455 291.750 242.625 291.920 ;
        RECT 242.815 291.750 242.985 291.920 ;
        RECT 245.925 291.750 246.095 291.920 ;
        RECT 246.285 291.750 246.455 291.920 ;
        RECT 252.155 291.750 252.325 291.920 ;
        RECT 252.515 291.750 252.685 291.920 ;
        RECT 255.625 291.750 255.795 291.920 ;
        RECT 255.985 291.750 256.155 291.920 ;
        RECT 259.095 291.750 259.265 291.920 ;
        RECT 259.455 291.750 259.625 291.920 ;
        RECT 262.565 291.750 262.735 291.920 ;
        RECT 262.925 291.750 263.095 291.920 ;
        RECT 266.035 291.750 266.205 291.920 ;
        RECT 266.395 291.750 266.565 291.920 ;
        RECT 272.265 291.750 272.435 291.920 ;
        RECT 272.625 291.750 272.795 291.920 ;
        RECT 275.735 291.750 275.905 291.920 ;
        RECT 276.095 291.750 276.265 291.920 ;
        RECT 279.205 291.750 279.375 291.920 ;
        RECT 279.565 291.750 279.735 291.920 ;
        RECT 282.675 291.750 282.845 291.920 ;
        RECT 283.035 291.750 283.205 291.920 ;
        RECT 286.145 291.750 286.315 291.920 ;
        RECT 286.505 291.750 286.675 291.920 ;
        RECT 97.885 290.010 98.055 290.180 ;
        RECT 98.245 290.010 98.415 290.180 ;
        RECT 101.355 290.010 101.525 290.180 ;
        RECT 101.715 290.010 101.885 290.180 ;
        RECT 18.195 289.740 18.365 289.910 ;
        RECT 18.555 289.740 18.725 289.910 ;
        RECT 21.665 289.740 21.835 289.910 ;
        RECT 22.025 289.740 22.195 289.910 ;
        RECT 25.135 289.740 25.305 289.910 ;
        RECT 25.495 289.740 25.665 289.910 ;
        RECT 31.565 289.770 31.735 289.940 ;
        RECT 31.925 289.770 32.095 289.940 ;
        RECT 35.035 289.770 35.205 289.940 ;
        RECT 35.395 289.770 35.565 289.940 ;
        RECT 38.505 289.770 38.675 289.940 ;
        RECT 38.865 289.770 39.035 289.940 ;
        RECT 44.795 289.770 44.965 289.940 ;
        RECT 45.155 289.770 45.325 289.940 ;
        RECT 48.265 289.770 48.435 289.940 ;
        RECT 48.625 289.770 48.795 289.940 ;
        RECT 51.735 289.770 51.905 289.940 ;
        RECT 52.095 289.770 52.265 289.940 ;
        RECT 58.065 289.740 58.235 289.910 ;
        RECT 58.425 289.740 58.595 289.910 ;
        RECT 61.535 289.740 61.705 289.910 ;
        RECT 61.895 289.740 62.065 289.910 ;
        RECT 65.005 289.740 65.175 289.910 ;
        RECT 65.365 289.740 65.535 289.910 ;
        RECT 71.335 289.770 71.505 289.940 ;
        RECT 71.695 289.770 71.865 289.940 ;
        RECT 74.805 289.770 74.975 289.940 ;
        RECT 75.165 289.770 75.335 289.940 ;
        RECT 78.275 289.770 78.445 289.940 ;
        RECT 78.635 289.770 78.805 289.940 ;
        RECT 84.465 289.790 84.635 289.960 ;
        RECT 84.825 289.790 84.995 289.960 ;
        RECT 87.935 289.790 88.105 289.960 ;
        RECT 88.295 289.790 88.465 289.960 ;
        RECT 91.405 289.790 91.575 289.960 ;
        RECT 91.765 289.790 91.935 289.960 ;
        RECT 4.855 283.180 5.025 283.350 ;
        RECT 5.215 283.180 5.385 283.350 ;
        RECT 8.325 283.180 8.495 283.350 ;
        RECT 8.685 283.180 8.855 283.350 ;
        RECT 11.795 283.180 11.965 283.350 ;
        RECT 12.155 283.180 12.325 283.350 ;
        RECT 613.450 292.415 613.620 292.585 ;
        RECT 616.280 292.330 616.450 292.500 ;
        RECT 620.665 292.495 620.835 292.665 ;
        RECT 836.140 293.645 836.310 293.815 ;
        RECT 639.300 291.550 639.470 291.720 ;
        RECT 836.140 293.285 836.310 293.455 ;
        RECT 842.425 294.255 842.595 294.425 ;
        RECT 840.565 293.385 840.735 293.555 ;
        RECT 594.345 291.005 594.515 291.175 ;
        RECT 594.705 291.005 594.875 291.175 ;
        RECT 379.140 289.765 379.310 289.935 ;
        RECT 379.140 289.405 379.310 289.575 ;
        RECT 212.075 285.170 212.245 285.340 ;
        RECT 212.435 285.170 212.605 285.340 ;
        RECT 215.545 285.170 215.715 285.340 ;
        RECT 215.905 285.170 216.075 285.340 ;
        RECT 219.015 285.170 219.185 285.340 ;
        RECT 219.375 285.170 219.545 285.340 ;
        RECT 222.485 285.170 222.655 285.340 ;
        RECT 222.845 285.170 223.015 285.340 ;
        RECT 225.955 285.170 226.125 285.340 ;
        RECT 226.315 285.170 226.485 285.340 ;
        RECT 232.045 285.170 232.215 285.340 ;
        RECT 232.405 285.170 232.575 285.340 ;
        RECT 235.515 285.170 235.685 285.340 ;
        RECT 235.875 285.170 236.045 285.340 ;
        RECT 238.985 285.170 239.155 285.340 ;
        RECT 239.345 285.170 239.515 285.340 ;
        RECT 242.455 285.170 242.625 285.340 ;
        RECT 242.815 285.170 242.985 285.340 ;
        RECT 245.925 285.170 246.095 285.340 ;
        RECT 246.285 285.170 246.455 285.340 ;
        RECT 252.155 285.170 252.325 285.340 ;
        RECT 252.515 285.170 252.685 285.340 ;
        RECT 255.625 285.170 255.795 285.340 ;
        RECT 255.985 285.170 256.155 285.340 ;
        RECT 259.095 285.170 259.265 285.340 ;
        RECT 259.455 285.170 259.625 285.340 ;
        RECT 262.565 285.170 262.735 285.340 ;
        RECT 262.925 285.170 263.095 285.340 ;
        RECT 266.035 285.170 266.205 285.340 ;
        RECT 266.395 285.170 266.565 285.340 ;
        RECT 272.265 285.170 272.435 285.340 ;
        RECT 272.625 285.170 272.795 285.340 ;
        RECT 275.735 285.170 275.905 285.340 ;
        RECT 276.095 285.170 276.265 285.340 ;
        RECT 279.205 285.170 279.375 285.340 ;
        RECT 279.565 285.170 279.735 285.340 ;
        RECT 282.675 285.170 282.845 285.340 ;
        RECT 283.035 285.170 283.205 285.340 ;
        RECT 286.145 285.170 286.315 285.340 ;
        RECT 286.505 285.170 286.675 285.340 ;
        RECT 294.505 284.335 295.755 286.305 ;
        RECT 379.140 286.295 379.310 286.465 ;
        RECT 379.140 285.935 379.310 286.105 ;
        RECT 97.885 283.430 98.055 283.600 ;
        RECT 98.245 283.430 98.415 283.600 ;
        RECT 101.355 283.430 101.525 283.600 ;
        RECT 101.715 283.430 101.885 283.600 ;
        RECT 18.195 283.160 18.365 283.330 ;
        RECT 18.555 283.160 18.725 283.330 ;
        RECT 21.665 283.160 21.835 283.330 ;
        RECT 22.025 283.160 22.195 283.330 ;
        RECT 25.135 283.160 25.305 283.330 ;
        RECT 25.495 283.160 25.665 283.330 ;
        RECT 31.565 283.190 31.735 283.360 ;
        RECT 31.925 283.190 32.095 283.360 ;
        RECT 35.035 283.190 35.205 283.360 ;
        RECT 35.395 283.190 35.565 283.360 ;
        RECT 38.505 283.190 38.675 283.360 ;
        RECT 38.865 283.190 39.035 283.360 ;
        RECT 44.795 283.190 44.965 283.360 ;
        RECT 45.155 283.190 45.325 283.360 ;
        RECT 48.265 283.190 48.435 283.360 ;
        RECT 48.625 283.190 48.795 283.360 ;
        RECT 51.735 283.190 51.905 283.360 ;
        RECT 52.095 283.190 52.265 283.360 ;
        RECT 58.065 283.160 58.235 283.330 ;
        RECT 58.425 283.160 58.595 283.330 ;
        RECT 61.535 283.160 61.705 283.330 ;
        RECT 61.895 283.160 62.065 283.330 ;
        RECT 65.005 283.160 65.175 283.330 ;
        RECT 65.365 283.160 65.535 283.330 ;
        RECT 71.335 283.190 71.505 283.360 ;
        RECT 71.695 283.190 71.865 283.360 ;
        RECT 74.805 283.190 74.975 283.360 ;
        RECT 75.165 283.190 75.335 283.360 ;
        RECT 78.275 283.190 78.445 283.360 ;
        RECT 78.635 283.190 78.805 283.360 ;
        RECT 84.465 283.210 84.635 283.380 ;
        RECT 84.825 283.210 84.995 283.380 ;
        RECT 87.935 283.210 88.105 283.380 ;
        RECT 88.295 283.210 88.465 283.380 ;
        RECT 91.405 283.210 91.575 283.380 ;
        RECT 91.765 283.210 91.935 283.380 ;
        RECT 4.855 276.600 5.025 276.770 ;
        RECT 5.215 276.600 5.385 276.770 ;
        RECT 8.325 276.600 8.495 276.770 ;
        RECT 8.685 276.600 8.855 276.770 ;
        RECT 11.795 276.600 11.965 276.770 ;
        RECT 12.155 276.600 12.325 276.770 ;
        RECT 118.365 277.780 118.535 277.950 ;
        RECT 118.725 277.780 118.895 277.950 ;
        RECT 121.835 277.780 122.005 277.950 ;
        RECT 122.195 277.780 122.365 277.950 ;
        RECT 125.305 277.780 125.475 277.950 ;
        RECT 125.665 277.780 125.835 277.950 ;
        RECT 128.775 277.780 128.945 277.950 ;
        RECT 129.135 277.780 129.305 277.950 ;
        RECT 132.245 277.780 132.415 277.950 ;
        RECT 132.605 277.780 132.775 277.950 ;
        RECT 135.715 277.780 135.885 277.950 ;
        RECT 136.075 277.780 136.245 277.950 ;
        RECT 139.185 277.780 139.355 277.950 ;
        RECT 139.545 277.780 139.715 277.950 ;
        RECT 142.655 277.780 142.825 277.950 ;
        RECT 143.015 277.780 143.185 277.950 ;
        RECT 146.125 277.780 146.295 277.950 ;
        RECT 146.485 277.780 146.655 277.950 ;
        RECT 149.595 277.780 149.765 277.950 ;
        RECT 149.955 277.780 150.125 277.950 ;
        RECT 97.885 276.850 98.055 277.020 ;
        RECT 98.245 276.850 98.415 277.020 ;
        RECT 101.355 276.850 101.525 277.020 ;
        RECT 101.715 276.850 101.885 277.020 ;
        RECT 18.195 276.580 18.365 276.750 ;
        RECT 18.555 276.580 18.725 276.750 ;
        RECT 21.665 276.580 21.835 276.750 ;
        RECT 22.025 276.580 22.195 276.750 ;
        RECT 25.135 276.580 25.305 276.750 ;
        RECT 25.495 276.580 25.665 276.750 ;
        RECT 31.565 276.610 31.735 276.780 ;
        RECT 31.925 276.610 32.095 276.780 ;
        RECT 35.035 276.610 35.205 276.780 ;
        RECT 35.395 276.610 35.565 276.780 ;
        RECT 38.505 276.610 38.675 276.780 ;
        RECT 38.865 276.610 39.035 276.780 ;
        RECT 44.795 276.610 44.965 276.780 ;
        RECT 45.155 276.610 45.325 276.780 ;
        RECT 48.265 276.610 48.435 276.780 ;
        RECT 48.625 276.610 48.795 276.780 ;
        RECT 51.735 276.610 51.905 276.780 ;
        RECT 52.095 276.610 52.265 276.780 ;
        RECT 58.065 276.580 58.235 276.750 ;
        RECT 58.425 276.580 58.595 276.750 ;
        RECT 61.535 276.580 61.705 276.750 ;
        RECT 61.895 276.580 62.065 276.750 ;
        RECT 65.005 276.580 65.175 276.750 ;
        RECT 65.365 276.580 65.535 276.750 ;
        RECT 71.335 276.610 71.505 276.780 ;
        RECT 71.695 276.610 71.865 276.780 ;
        RECT 74.805 276.610 74.975 276.780 ;
        RECT 75.165 276.610 75.335 276.780 ;
        RECT 78.275 276.610 78.445 276.780 ;
        RECT 78.635 276.610 78.805 276.780 ;
        RECT 84.465 276.630 84.635 276.800 ;
        RECT 84.825 276.630 84.995 276.800 ;
        RECT 87.935 276.630 88.105 276.800 ;
        RECT 88.295 276.630 88.465 276.800 ;
        RECT 91.405 276.630 91.575 276.800 ;
        RECT 91.765 276.630 91.935 276.800 ;
        RECT 118.365 271.200 118.535 271.370 ;
        RECT 118.725 271.200 118.895 271.370 ;
        RECT 121.835 271.200 122.005 271.370 ;
        RECT 122.195 271.200 122.365 271.370 ;
        RECT 125.305 271.200 125.475 271.370 ;
        RECT 125.665 271.200 125.835 271.370 ;
        RECT 128.775 271.200 128.945 271.370 ;
        RECT 129.135 271.200 129.305 271.370 ;
        RECT 132.245 271.200 132.415 271.370 ;
        RECT 132.605 271.200 132.775 271.370 ;
        RECT 135.715 271.200 135.885 271.370 ;
        RECT 136.075 271.200 136.245 271.370 ;
        RECT 139.185 271.200 139.355 271.370 ;
        RECT 139.545 271.200 139.715 271.370 ;
        RECT 142.655 271.200 142.825 271.370 ;
        RECT 143.015 271.200 143.185 271.370 ;
        RECT 146.125 271.200 146.295 271.370 ;
        RECT 146.485 271.200 146.655 271.370 ;
        RECT 149.595 271.200 149.765 271.370 ;
        RECT 149.955 271.200 150.125 271.370 ;
        RECT 97.885 270.270 98.055 270.440 ;
        RECT 98.245 270.270 98.415 270.440 ;
        RECT 101.355 270.270 101.525 270.440 ;
        RECT 101.715 270.270 101.885 270.440 ;
        RECT 4.855 270.020 5.025 270.190 ;
        RECT 5.215 270.020 5.385 270.190 ;
        RECT 8.325 270.020 8.495 270.190 ;
        RECT 8.685 270.020 8.855 270.190 ;
        RECT 11.795 270.020 11.965 270.190 ;
        RECT 12.155 270.020 12.325 270.190 ;
        RECT 18.195 270.000 18.365 270.170 ;
        RECT 18.555 270.000 18.725 270.170 ;
        RECT 21.665 270.000 21.835 270.170 ;
        RECT 22.025 270.000 22.195 270.170 ;
        RECT 25.135 270.000 25.305 270.170 ;
        RECT 25.495 270.000 25.665 270.170 ;
        RECT 31.565 270.030 31.735 270.200 ;
        RECT 31.925 270.030 32.095 270.200 ;
        RECT 35.035 270.030 35.205 270.200 ;
        RECT 35.395 270.030 35.565 270.200 ;
        RECT 38.505 270.030 38.675 270.200 ;
        RECT 38.865 270.030 39.035 270.200 ;
        RECT 44.795 270.030 44.965 270.200 ;
        RECT 45.155 270.030 45.325 270.200 ;
        RECT 48.265 270.030 48.435 270.200 ;
        RECT 48.625 270.030 48.795 270.200 ;
        RECT 51.735 270.030 51.905 270.200 ;
        RECT 52.095 270.030 52.265 270.200 ;
        RECT 58.065 270.000 58.235 270.170 ;
        RECT 58.425 270.000 58.595 270.170 ;
        RECT 61.535 270.000 61.705 270.170 ;
        RECT 61.895 270.000 62.065 270.170 ;
        RECT 65.005 270.000 65.175 270.170 ;
        RECT 65.365 270.000 65.535 270.170 ;
        RECT 71.335 270.030 71.505 270.200 ;
        RECT 71.695 270.030 71.865 270.200 ;
        RECT 74.805 270.030 74.975 270.200 ;
        RECT 75.165 270.030 75.335 270.200 ;
        RECT 78.275 270.030 78.445 270.200 ;
        RECT 78.635 270.030 78.805 270.200 ;
        RECT 84.465 270.050 84.635 270.220 ;
        RECT 84.825 270.050 84.995 270.220 ;
        RECT 87.935 270.050 88.105 270.220 ;
        RECT 88.295 270.050 88.465 270.220 ;
        RECT 91.405 270.050 91.575 270.220 ;
        RECT 91.765 270.050 91.935 270.220 ;
        RECT 379.140 282.825 379.310 282.995 ;
        RECT 379.140 282.465 379.310 282.635 ;
        RECT 379.140 279.355 379.310 279.525 ;
        RECT 379.140 278.995 379.310 279.165 ;
        RECT 379.140 275.885 379.310 276.055 ;
        RECT 385.720 289.765 385.890 289.935 ;
        RECT 597.000 290.670 597.530 291.200 ;
        RECT 633.910 290.265 634.440 290.795 ;
        RECT 631.435 289.880 631.605 290.050 ;
        RECT 631.795 289.880 631.965 290.050 ;
        RECT 385.720 289.405 385.890 289.575 ;
        RECT 610.200 288.595 610.370 288.765 ;
        RECT 610.990 288.595 611.160 288.765 ;
        RECT 611.780 288.595 611.950 288.765 ;
        RECT 612.570 288.595 612.740 288.765 ;
        RECT 613.360 288.595 613.530 288.765 ;
        RECT 617.790 288.565 617.960 288.735 ;
        RECT 618.580 288.565 618.750 288.735 ;
        RECT 619.370 288.565 619.540 288.735 ;
        RECT 620.160 288.565 620.330 288.735 ;
        RECT 620.950 288.565 621.120 288.735 ;
        RECT 600.750 287.815 600.920 287.985 ;
        RECT 601.540 287.815 601.710 287.985 ;
        RECT 602.330 287.815 602.500 287.985 ;
        RECT 603.120 287.815 603.290 287.985 ;
        RECT 603.910 287.815 604.080 287.985 ;
        RECT 615.440 288.075 615.610 288.245 ;
        RECT 627.530 287.945 627.700 288.115 ;
        RECT 628.320 287.945 628.490 288.115 ;
        RECT 629.110 287.945 629.280 288.115 ;
        RECT 629.900 287.945 630.070 288.115 ;
        RECT 630.690 287.945 630.860 288.115 ;
        RECT 385.720 286.295 385.890 286.465 ;
        RECT 385.720 285.935 385.890 286.105 ;
        RECT 591.910 287.330 592.080 287.500 ;
        RECT 641.785 290.925 641.955 291.095 ;
        RECT 645.330 291.370 645.500 291.540 ;
        RECT 819.185 290.805 819.355 290.975 ;
        RECT 694.840 288.555 696.090 290.525 ;
        RECT 820.115 290.580 820.285 290.750 ;
        RECT 832.810 291.725 834.060 292.975 ;
        RECT 821.965 290.450 822.135 290.620 ;
        RECT 824.635 288.820 824.805 288.990 ;
        RECT 827.575 289.055 827.745 289.225 ;
        RECT 825.560 288.050 825.730 288.220 ;
        RECT 591.910 286.970 592.080 287.140 ;
        RECT 610.200 287.125 610.370 287.295 ;
        RECT 610.990 287.125 611.160 287.295 ;
        RECT 611.780 287.125 611.950 287.295 ;
        RECT 612.570 287.125 612.740 287.295 ;
        RECT 613.360 287.125 613.530 287.295 ;
        RECT 614.030 287.075 614.200 287.245 ;
        RECT 615.610 287.075 615.780 287.245 ;
        RECT 617.190 287.075 617.360 287.245 ;
        RECT 617.790 287.095 617.960 287.265 ;
        RECT 618.580 287.095 618.750 287.265 ;
        RECT 619.370 287.095 619.540 287.265 ;
        RECT 620.160 287.095 620.330 287.265 ;
        RECT 620.950 287.095 621.120 287.265 ;
        RECT 639.775 287.155 639.945 287.325 ;
        RECT 591.910 286.610 592.080 286.780 ;
        RECT 591.910 286.250 592.080 286.420 ;
        RECT 600.750 286.345 600.920 286.515 ;
        RECT 601.540 286.345 601.710 286.515 ;
        RECT 602.330 286.345 602.500 286.515 ;
        RECT 603.120 286.345 603.290 286.515 ;
        RECT 608.570 286.615 608.740 286.785 ;
        RECT 832.105 289.035 832.275 289.205 ;
        RECT 833.420 288.735 833.590 288.905 ;
        RECT 834.070 288.575 834.240 288.745 ;
        RECT 846.705 292.165 846.875 292.335 ;
        RECT 849.190 291.890 849.720 292.420 ;
        RECT 643.810 287.205 643.980 287.375 ;
        RECT 821.930 287.130 822.100 287.300 ;
        RECT 623.170 286.610 623.340 286.780 ;
        RECT 603.910 286.345 604.080 286.515 ;
        RECT 627.530 286.475 627.700 286.645 ;
        RECT 628.320 286.475 628.490 286.645 ;
        RECT 629.110 286.475 629.280 286.645 ;
        RECT 629.900 286.475 630.070 286.645 ;
        RECT 630.690 286.475 630.860 286.645 ;
        RECT 639.380 286.185 639.550 286.355 ;
        RECT 643.430 286.235 643.600 286.405 ;
        RECT 591.910 285.890 592.080 286.060 ;
        RECT 591.910 285.530 592.080 285.700 ;
        RECT 606.450 285.605 606.620 285.775 ;
        RECT 607.240 285.605 607.410 285.775 ;
        RECT 608.030 285.605 608.200 285.775 ;
        RECT 608.820 285.605 608.990 285.775 ;
        RECT 609.610 285.605 609.780 285.775 ;
        RECT 610.200 285.655 610.370 285.825 ;
        RECT 610.990 285.655 611.160 285.825 ;
        RECT 611.780 285.655 611.950 285.825 ;
        RECT 612.570 285.655 612.740 285.825 ;
        RECT 613.360 285.655 613.530 285.825 ;
        RECT 614.030 285.605 614.200 285.775 ;
        RECT 615.610 285.605 615.780 285.775 ;
        RECT 617.190 285.605 617.360 285.775 ;
        RECT 617.790 285.625 617.960 285.795 ;
        RECT 618.580 285.625 618.750 285.795 ;
        RECT 619.370 285.625 619.540 285.795 ;
        RECT 620.160 285.625 620.330 285.795 ;
        RECT 620.950 285.625 621.120 285.795 ;
        RECT 621.540 285.605 621.710 285.775 ;
        RECT 622.330 285.605 622.500 285.775 ;
        RECT 623.120 285.605 623.290 285.775 ;
        RECT 623.910 285.605 624.080 285.775 ;
        RECT 624.700 285.605 624.870 285.775 ;
        RECT 819.140 285.555 819.310 285.725 ;
        RECT 602.145 284.695 602.315 284.865 ;
        RECT 602.505 284.695 602.675 284.865 ;
        RECT 820.085 285.250 820.255 285.420 ;
        RECT 840.580 288.250 840.750 288.420 ;
        RECT 857.030 289.740 857.200 289.910 ;
        RECT 862.810 291.865 862.980 292.035 ;
        RECT 865.290 291.835 866.180 292.365 ;
        RECT 385.720 282.825 385.890 282.995 ;
        RECT 385.720 282.465 385.890 282.635 ;
        RECT 591.910 284.175 592.080 284.345 ;
        RECT 591.910 283.815 592.080 283.985 ;
        RECT 591.910 283.455 592.080 283.625 ;
        RECT 591.910 283.095 592.080 283.265 ;
        RECT 591.910 282.735 592.080 282.905 ;
        RECT 591.910 282.375 592.080 282.545 ;
        RECT 680.075 280.075 680.245 280.245 ;
        RECT 385.720 279.355 385.890 279.525 ;
        RECT 385.720 278.995 385.890 279.165 ;
        RECT 700.170 279.735 700.340 279.905 ;
        RECT 683.350 279.250 683.520 279.420 ;
        RECT 717.935 279.730 718.105 279.900 ;
        RECT 700.610 279.215 700.780 279.385 ;
        RECT 735.175 279.760 735.345 279.930 ;
        RECT 718.410 279.225 718.580 279.395 ;
        RECT 752.655 279.720 752.825 279.890 ;
        RECT 735.650 279.235 735.820 279.405 ;
        RECT 799.755 281.095 799.925 281.265 ;
        RECT 802.060 280.610 802.950 281.500 ;
        RECT 821.835 281.130 822.005 281.300 ;
        RECT 820.915 280.630 821.085 280.800 ;
        RECT 823.425 280.615 823.595 280.785 ;
        RECT 825.410 280.455 825.940 280.985 ;
        RECT 828.180 280.415 828.350 280.585 ;
        RECT 831.000 280.965 831.170 281.135 ;
        RECT 829.135 280.405 829.305 280.575 ;
        RECT 829.135 280.045 829.305 280.215 ;
        RECT 835.410 280.905 835.580 281.075 ;
        RECT 836.740 280.655 836.910 280.825 ;
        RECT 841.175 281.280 841.345 281.450 ;
        RECT 837.325 280.410 837.495 280.580 ;
        RECT 838.760 280.395 838.930 280.565 ;
        RECT 843.975 280.950 844.145 281.120 ;
        RECT 841.150 280.350 841.320 280.520 ;
        RECT 842.055 280.005 842.225 280.175 ;
        RECT 753.115 279.205 753.285 279.375 ;
        RECT 632.680 277.725 633.210 278.615 ;
        RECT 848.445 280.900 848.615 281.070 ;
        RECT 849.795 280.715 849.965 280.885 ;
        RECT 850.385 280.495 850.555 280.665 ;
        RECT 856.110 284.730 856.280 284.900 ;
        RECT 857.095 284.240 857.265 284.410 ;
        RECT 858.940 284.415 859.110 284.585 ;
        RECT 861.880 282.765 862.050 282.935 ;
        RECT 862.860 282.580 863.030 282.750 ;
        RECT 865.270 282.835 865.440 283.005 ;
        RECT 865.630 282.835 865.800 283.005 ;
        RECT 865.335 281.235 865.865 282.125 ;
        RECT 858.960 280.685 859.130 280.855 ;
        RECT 603.140 276.355 603.310 276.525 ;
        RECT 604.720 276.355 604.890 276.525 ;
        RECT 607.660 276.365 607.830 276.535 ;
        RECT 609.240 276.365 609.410 276.535 ;
        RECT 612.180 276.365 612.350 276.535 ;
        RECT 613.760 276.365 613.930 276.535 ;
        RECT 616.610 276.345 616.780 276.515 ;
        RECT 618.190 276.345 618.360 276.515 ;
        RECT 620.990 276.355 621.160 276.525 ;
        RECT 622.570 276.355 622.740 276.525 ;
        RECT 625.310 276.345 625.480 276.515 ;
        RECT 626.890 276.345 627.060 276.515 ;
        RECT 385.720 275.885 385.890 276.055 ;
        RECT 379.140 275.525 379.310 275.695 ;
        RECT 385.720 275.525 385.890 275.695 ;
        RECT 603.140 274.885 603.310 275.055 ;
        RECT 604.720 274.885 604.890 275.055 ;
        RECT 607.660 274.895 607.830 275.065 ;
        RECT 609.240 274.895 609.410 275.065 ;
        RECT 612.180 274.895 612.350 275.065 ;
        RECT 613.760 274.895 613.930 275.065 ;
        RECT 616.610 274.875 616.780 275.045 ;
        RECT 618.190 274.875 618.360 275.045 ;
        RECT 620.990 274.885 621.160 275.055 ;
        RECT 622.570 274.885 622.740 275.055 ;
        RECT 625.310 274.875 625.480 275.045 ;
        RECT 626.890 274.875 627.060 275.045 ;
        RECT 613.370 273.945 613.540 274.115 ;
        RECT 616.200 273.860 616.370 274.030 ;
        RECT 620.585 274.025 620.755 274.195 ;
        RECT 639.220 273.080 639.390 273.250 ;
        RECT 681.885 274.510 682.055 274.680 ;
        RECT 683.255 274.130 683.425 274.300 ;
        RECT 683.885 274.400 684.055 274.570 ;
        RECT 594.265 272.535 594.435 272.705 ;
        RECT 594.625 272.535 594.795 272.705 ;
        RECT 596.920 272.200 597.450 272.730 ;
        RECT 633.830 271.795 634.360 272.325 ;
        RECT 631.675 271.325 631.845 271.495 ;
        RECT 379.160 270.905 379.330 271.075 ;
        RECT 379.160 270.545 379.330 270.715 ;
        RECT 379.160 267.435 379.330 267.605 ;
        RECT 379.160 267.075 379.330 267.245 ;
        RECT 379.160 263.965 379.330 264.135 ;
        RECT 379.160 263.605 379.330 263.775 ;
        RECT 379.160 260.495 379.330 260.665 ;
        RECT 379.160 260.135 379.330 260.305 ;
        RECT 379.160 257.025 379.330 257.195 ;
        RECT 385.740 270.905 385.910 271.075 ;
        RECT 385.740 270.545 385.910 270.715 ;
        RECT 610.120 270.125 610.290 270.295 ;
        RECT 610.910 270.125 611.080 270.295 ;
        RECT 611.700 270.125 611.870 270.295 ;
        RECT 612.490 270.125 612.660 270.295 ;
        RECT 613.280 270.125 613.450 270.295 ;
        RECT 617.710 270.095 617.880 270.265 ;
        RECT 618.500 270.095 618.670 270.265 ;
        RECT 619.290 270.095 619.460 270.265 ;
        RECT 620.080 270.095 620.250 270.265 ;
        RECT 620.870 270.095 621.040 270.265 ;
        RECT 600.670 269.345 600.840 269.515 ;
        RECT 385.740 267.435 385.910 267.605 ;
        RECT 385.740 267.075 385.910 267.245 ;
        RECT 591.750 269.070 591.920 269.240 ;
        RECT 601.460 269.345 601.630 269.515 ;
        RECT 602.250 269.345 602.420 269.515 ;
        RECT 603.040 269.345 603.210 269.515 ;
        RECT 603.830 269.345 604.000 269.515 ;
        RECT 615.360 269.605 615.530 269.775 ;
        RECT 627.450 269.475 627.620 269.645 ;
        RECT 628.240 269.475 628.410 269.645 ;
        RECT 629.030 269.475 629.200 269.645 ;
        RECT 629.820 269.475 629.990 269.645 ;
        RECT 630.610 269.475 630.780 269.645 ;
        RECT 641.705 272.455 641.875 272.625 ;
        RECT 645.250 272.900 645.420 273.070 ;
        RECT 689.195 274.410 689.365 274.580 ;
        RECT 690.535 274.120 690.705 274.290 ;
        RECT 691.105 274.090 691.275 274.260 ;
        RECT 700.485 274.150 700.655 274.320 ;
        RECT 701.115 274.420 701.285 274.590 ;
        RECT 706.425 274.430 706.595 274.600 ;
        RECT 707.765 274.140 707.935 274.310 ;
        RECT 708.335 274.110 708.505 274.280 ;
        RECT 718.055 274.250 718.225 274.420 ;
        RECT 718.685 274.520 718.855 274.690 ;
        RECT 723.995 274.530 724.165 274.700 ;
        RECT 725.335 274.240 725.505 274.410 ;
        RECT 725.905 274.210 726.075 274.380 ;
        RECT 735.225 274.280 735.395 274.450 ;
        RECT 735.855 274.550 736.025 274.720 ;
        RECT 741.165 274.560 741.335 274.730 ;
        RECT 742.505 274.270 742.675 274.440 ;
        RECT 743.075 274.240 743.245 274.410 ;
        RECT 753.035 274.340 753.205 274.510 ;
        RECT 753.665 274.610 753.835 274.780 ;
        RECT 758.975 274.620 759.145 274.790 ;
        RECT 760.885 274.300 761.055 274.470 ;
        RECT 783.035 273.360 783.205 273.530 ;
        RECT 784.450 272.340 784.620 272.510 ;
        RECT 785.435 273.360 785.605 273.530 ;
        RECT 790.715 273.360 790.885 273.530 ;
        RECT 795.955 274.075 796.125 274.245 ;
        RECT 795.955 273.715 796.125 273.885 ;
        RECT 801.925 273.350 802.095 273.520 ;
        RECT 803.355 272.380 803.525 272.550 ;
        RECT 804.325 273.350 804.495 273.520 ;
        RECT 814.835 274.410 815.005 274.580 ;
        RECT 809.605 273.350 809.775 273.520 ;
        RECT 814.835 274.050 815.005 274.220 ;
        RECT 820.775 273.320 820.945 273.490 ;
        RECT 822.195 272.385 822.365 272.555 ;
        RECT 823.175 273.320 823.345 273.490 ;
        RECT 828.455 273.320 828.625 273.490 ;
        RECT 833.690 274.205 833.860 274.375 ;
        RECT 833.690 273.845 833.860 274.015 ;
        RECT 839.280 273.685 839.450 273.855 ;
        RECT 851.980 274.830 852.510 275.360 ;
        RECT 857.105 278.990 857.275 279.160 ;
        RECT 841.910 273.265 842.080 273.435 ;
        RECT 839.085 272.300 839.255 272.470 ;
        RECT 839.930 272.855 840.100 273.025 ;
        RECT 841.910 272.905 842.080 273.075 ;
        RECT 591.750 268.710 591.920 268.880 ;
        RECT 610.120 268.655 610.290 268.825 ;
        RECT 610.910 268.655 611.080 268.825 ;
        RECT 611.700 268.655 611.870 268.825 ;
        RECT 612.490 268.655 612.660 268.825 ;
        RECT 613.280 268.655 613.450 268.825 ;
        RECT 613.950 268.605 614.120 268.775 ;
        RECT 591.750 268.350 591.920 268.520 ;
        RECT 615.530 268.605 615.700 268.775 ;
        RECT 617.110 268.605 617.280 268.775 ;
        RECT 617.710 268.625 617.880 268.795 ;
        RECT 618.500 268.625 618.670 268.795 ;
        RECT 619.290 268.625 619.460 268.795 ;
        RECT 620.080 268.625 620.250 268.795 ;
        RECT 620.870 268.625 621.040 268.795 ;
        RECT 639.695 268.685 639.865 268.855 ;
        RECT 591.750 267.990 591.920 268.160 ;
        RECT 591.750 267.630 591.920 267.800 ;
        RECT 600.670 267.875 600.840 268.045 ;
        RECT 601.460 267.875 601.630 268.045 ;
        RECT 602.250 267.875 602.420 268.045 ;
        RECT 603.040 267.875 603.210 268.045 ;
        RECT 608.490 268.145 608.660 268.315 ;
        RECT 682.945 269.420 683.115 269.590 ;
        RECT 643.730 268.735 643.900 268.905 ;
        RECT 623.090 268.140 623.260 268.310 ;
        RECT 680.145 268.340 680.315 268.510 ;
        RECT 603.830 267.875 604.000 268.045 ;
        RECT 627.450 268.005 627.620 268.175 ;
        RECT 628.240 268.005 628.410 268.175 ;
        RECT 629.030 268.005 629.200 268.175 ;
        RECT 629.820 268.005 629.990 268.175 ;
        RECT 630.610 268.005 630.780 268.175 ;
        RECT 639.300 267.715 639.470 267.885 ;
        RECT 643.350 267.765 643.520 267.935 ;
        RECT 681.075 268.155 681.245 268.325 ;
        RECT 591.750 267.270 591.920 267.440 ;
        RECT 606.370 267.135 606.540 267.305 ;
        RECT 607.160 267.135 607.330 267.305 ;
        RECT 607.950 267.135 608.120 267.305 ;
        RECT 608.740 267.135 608.910 267.305 ;
        RECT 609.530 267.135 609.700 267.305 ;
        RECT 610.120 267.185 610.290 267.355 ;
        RECT 610.910 267.185 611.080 267.355 ;
        RECT 611.700 267.185 611.870 267.355 ;
        RECT 612.490 267.185 612.660 267.355 ;
        RECT 613.280 267.185 613.450 267.355 ;
        RECT 613.950 267.135 614.120 267.305 ;
        RECT 615.530 267.135 615.700 267.305 ;
        RECT 617.110 267.135 617.280 267.305 ;
        RECT 617.710 267.155 617.880 267.325 ;
        RECT 618.500 267.155 618.670 267.325 ;
        RECT 619.290 267.155 619.460 267.325 ;
        RECT 620.080 267.155 620.250 267.325 ;
        RECT 620.870 267.155 621.040 267.325 ;
        RECT 621.460 267.135 621.630 267.305 ;
        RECT 622.250 267.135 622.420 267.305 ;
        RECT 623.040 267.135 623.210 267.305 ;
        RECT 623.830 267.135 624.000 267.305 ;
        RECT 685.830 268.430 686.000 268.600 ;
        RECT 688.645 268.630 688.815 268.800 ;
        RECT 686.775 268.235 686.945 268.405 ;
        RECT 686.775 267.875 686.945 268.045 ;
        RECT 691.590 268.140 691.760 268.310 ;
        RECT 700.175 269.440 700.345 269.610 ;
        RECT 692.530 268.410 692.700 268.580 ;
        RECT 693.950 268.575 694.120 268.745 ;
        RECT 698.305 268.175 698.475 268.345 ;
        RECT 703.060 268.450 703.230 268.620 ;
        RECT 705.875 268.650 706.045 268.820 ;
        RECT 704.005 268.255 704.175 268.425 ;
        RECT 704.005 267.895 704.175 268.065 ;
        RECT 708.820 268.160 708.990 268.330 ;
        RECT 717.745 269.540 717.915 269.710 ;
        RECT 709.760 268.430 709.930 268.600 ;
        RECT 711.180 268.595 711.350 268.765 ;
        RECT 715.875 268.275 716.045 268.445 ;
        RECT 720.630 268.550 720.800 268.720 ;
        RECT 723.445 268.750 723.615 268.920 ;
        RECT 721.575 268.355 721.745 268.525 ;
        RECT 721.575 267.995 721.745 268.165 ;
        RECT 726.390 268.260 726.560 268.430 ;
        RECT 734.915 269.570 735.085 269.740 ;
        RECT 727.330 268.530 727.500 268.700 ;
        RECT 728.750 268.695 728.920 268.865 ;
        RECT 733.045 268.305 733.215 268.475 ;
        RECT 737.800 268.580 737.970 268.750 ;
        RECT 740.615 268.780 740.785 268.950 ;
        RECT 738.745 268.385 738.915 268.555 ;
        RECT 738.745 268.025 738.915 268.195 ;
        RECT 743.560 268.290 743.730 268.460 ;
        RECT 752.725 269.630 752.895 269.800 ;
        RECT 744.500 268.560 744.670 268.730 ;
        RECT 745.920 268.725 746.090 268.895 ;
        RECT 750.855 268.365 751.025 268.535 ;
        RECT 755.610 268.640 755.780 268.810 ;
        RECT 758.425 268.840 758.595 269.010 ;
        RECT 761.370 268.350 761.540 268.520 ;
        RECT 844.890 270.785 845.060 270.955 ;
        RECT 852.000 272.845 852.530 273.735 ;
        RECT 857.100 272.265 857.270 272.435 ;
        RECT 845.850 270.100 846.020 270.270 ;
        RECT 762.310 268.620 762.480 268.790 ;
        RECT 763.730 268.785 763.900 268.955 ;
        RECT 624.620 267.135 624.790 267.305 ;
        RECT 601.525 266.235 601.695 266.405 ;
        RECT 601.885 266.235 602.055 266.405 ;
        RECT 602.245 266.235 602.415 266.405 ;
        RECT 385.740 263.965 385.910 264.135 ;
        RECT 591.750 265.915 591.920 266.085 ;
        RECT 591.750 265.555 591.920 265.725 ;
        RECT 591.750 265.195 591.920 265.365 ;
        RECT 591.750 264.835 591.920 265.005 ;
        RECT 591.750 264.475 591.920 264.645 ;
        RECT 783.045 265.800 783.215 265.970 ;
        RECT 784.475 264.860 784.645 265.030 ;
        RECT 785.445 265.800 785.615 265.970 ;
        RECT 795.945 266.870 796.115 267.040 ;
        RECT 790.725 265.800 790.895 265.970 ;
        RECT 795.945 266.510 796.115 266.680 ;
        RECT 801.575 265.860 801.745 266.030 ;
        RECT 803.000 264.895 803.170 265.065 ;
        RECT 803.975 265.860 804.145 266.030 ;
        RECT 809.255 265.860 809.425 266.030 ;
        RECT 838.645 267.410 838.815 267.580 ;
        RECT 841.460 267.875 841.630 268.045 ;
        RECT 814.480 266.615 814.650 266.785 ;
        RECT 839.580 266.800 839.750 266.970 ;
        RECT 841.460 267.515 841.630 267.685 ;
        RECT 852.615 270.895 852.785 271.065 ;
        RECT 852.615 270.535 852.785 270.705 ;
        RECT 862.850 269.215 863.020 269.385 ;
        RECT 865.450 268.990 866.700 269.880 ;
        RECT 859.035 267.440 859.205 267.610 ;
        RECT 853.750 265.660 853.920 265.830 ;
        RECT 591.750 264.115 591.920 264.285 ;
        RECT 385.740 263.605 385.910 263.775 ;
        RECT 385.740 260.495 385.910 260.665 ;
        RECT 385.740 260.135 385.910 260.305 ;
        RECT 632.515 260.245 633.405 260.775 ;
        RECT 602.990 258.625 603.160 258.795 ;
        RECT 604.570 258.625 604.740 258.795 ;
        RECT 607.510 258.635 607.680 258.805 ;
        RECT 609.090 258.635 609.260 258.805 ;
        RECT 612.030 258.635 612.200 258.805 ;
        RECT 613.610 258.635 613.780 258.805 ;
        RECT 616.460 258.615 616.630 258.785 ;
        RECT 618.040 258.615 618.210 258.785 ;
        RECT 620.840 258.625 621.010 258.795 ;
        RECT 622.420 258.625 622.590 258.795 ;
        RECT 625.160 258.615 625.330 258.785 ;
        RECT 626.740 258.615 626.910 258.785 ;
        RECT 680.055 258.545 680.225 258.715 ;
        RECT 385.740 257.025 385.910 257.195 ;
        RECT 602.990 257.155 603.160 257.325 ;
        RECT 604.570 257.155 604.740 257.325 ;
        RECT 607.510 257.165 607.680 257.335 ;
        RECT 609.090 257.165 609.260 257.335 ;
        RECT 612.030 257.165 612.200 257.335 ;
        RECT 613.610 257.165 613.780 257.335 ;
        RECT 616.460 257.145 616.630 257.315 ;
        RECT 379.160 256.665 379.330 256.835 ;
        RECT 618.040 257.145 618.210 257.315 ;
        RECT 620.840 257.155 621.010 257.325 ;
        RECT 622.420 257.155 622.590 257.325 ;
        RECT 625.160 257.145 625.330 257.315 ;
        RECT 626.740 257.145 626.910 257.315 ;
        RECT 385.740 256.665 385.910 256.835 ;
        RECT 613.220 256.215 613.390 256.385 ;
        RECT 616.050 256.130 616.220 256.300 ;
        RECT 620.435 256.295 620.605 256.465 ;
        RECT 386.920 254.380 388.170 254.910 ;
        RECT 639.070 255.350 639.240 255.520 ;
        RECT 700.150 258.205 700.320 258.375 ;
        RECT 683.330 257.720 683.500 257.890 ;
        RECT 717.915 258.200 718.085 258.370 ;
        RECT 700.590 257.685 700.760 257.855 ;
        RECT 735.155 258.230 735.325 258.400 ;
        RECT 718.390 257.695 718.560 257.865 ;
        RECT 752.635 258.190 752.805 258.360 ;
        RECT 735.630 257.705 735.800 257.875 ;
        RECT 753.095 257.675 753.265 257.845 ;
        RECT 594.115 254.805 594.285 254.975 ;
        RECT 594.475 254.805 594.645 254.975 ;
        RECT 596.770 254.470 597.300 255.000 ;
        RECT 633.680 254.065 634.210 254.595 ;
        RECT 631.380 253.655 631.550 253.825 ;
        RECT 631.740 253.655 631.910 253.825 ;
        RECT 609.970 252.395 610.140 252.565 ;
        RECT 610.760 252.395 610.930 252.565 ;
        RECT 611.550 252.395 611.720 252.565 ;
        RECT 612.340 252.395 612.510 252.565 ;
        RECT 613.130 252.395 613.300 252.565 ;
        RECT 617.560 252.365 617.730 252.535 ;
        RECT 618.350 252.365 618.520 252.535 ;
        RECT 619.140 252.365 619.310 252.535 ;
        RECT 619.930 252.365 620.100 252.535 ;
        RECT 620.720 252.365 620.890 252.535 ;
        RECT 600.520 251.615 600.690 251.785 ;
        RECT 601.310 251.615 601.480 251.785 ;
        RECT 602.100 251.615 602.270 251.785 ;
        RECT 602.890 251.615 603.060 251.785 ;
        RECT 603.680 251.615 603.850 251.785 ;
        RECT 615.210 251.875 615.380 252.045 ;
        RECT 627.300 251.745 627.470 251.915 ;
        RECT 628.090 251.745 628.260 251.915 ;
        RECT 628.880 251.745 629.050 251.915 ;
        RECT 629.670 251.745 629.840 251.915 ;
        RECT 630.460 251.745 630.630 251.915 ;
        RECT 641.555 254.725 641.725 254.895 ;
        RECT 645.100 255.170 645.270 255.340 ;
        RECT 683.235 252.600 683.405 252.770 ;
        RECT 683.865 252.870 684.035 253.040 ;
        RECT 689.175 252.880 689.345 253.050 ;
        RECT 690.515 252.590 690.685 252.760 ;
        RECT 691.085 252.560 691.255 252.730 ;
        RECT 700.465 252.620 700.635 252.790 ;
        RECT 701.095 252.890 701.265 253.060 ;
        RECT 706.405 252.900 706.575 253.070 ;
        RECT 707.745 252.610 707.915 252.780 ;
        RECT 708.315 252.580 708.485 252.750 ;
        RECT 718.035 252.720 718.205 252.890 ;
        RECT 718.665 252.990 718.835 253.160 ;
        RECT 723.975 253.000 724.145 253.170 ;
        RECT 725.315 252.710 725.485 252.880 ;
        RECT 725.885 252.680 726.055 252.850 ;
        RECT 735.205 252.750 735.375 252.920 ;
        RECT 735.835 253.020 736.005 253.190 ;
        RECT 741.145 253.030 741.315 253.200 ;
        RECT 742.485 252.740 742.655 252.910 ;
        RECT 743.055 252.710 743.225 252.880 ;
        RECT 753.015 252.810 753.185 252.980 ;
        RECT 753.645 253.080 753.815 253.250 ;
        RECT 758.955 253.090 759.125 253.260 ;
        RECT 760.865 252.770 761.035 252.940 ;
        RECT 609.970 250.925 610.140 251.095 ;
        RECT 610.760 250.925 610.930 251.095 ;
        RECT 611.550 250.925 611.720 251.095 ;
        RECT 612.340 250.925 612.510 251.095 ;
        RECT 613.130 250.925 613.300 251.095 ;
        RECT 613.800 250.875 613.970 251.045 ;
        RECT 615.380 250.875 615.550 251.045 ;
        RECT 616.960 250.875 617.130 251.045 ;
        RECT 617.560 250.895 617.730 251.065 ;
        RECT 618.350 250.895 618.520 251.065 ;
        RECT 619.140 250.895 619.310 251.065 ;
        RECT 619.930 250.895 620.100 251.065 ;
        RECT 620.720 250.895 620.890 251.065 ;
        RECT 639.545 250.955 639.715 251.125 ;
        RECT 591.520 250.270 591.690 250.440 ;
        RECT 591.520 249.910 591.690 250.080 ;
        RECT 600.520 250.145 600.690 250.315 ;
        RECT 601.310 250.145 601.480 250.315 ;
        RECT 602.100 250.145 602.270 250.315 ;
        RECT 602.890 250.145 603.060 250.315 ;
        RECT 608.340 250.415 608.510 250.585 ;
        RECT 857.195 265.675 857.365 265.845 ;
        RECT 856.120 256.775 856.290 256.945 ;
        RECT 858.890 256.710 859.060 256.880 ;
        RECT 857.070 256.325 857.240 256.495 ;
        RECT 854.760 253.870 855.290 254.400 ;
        RECT 862.805 254.375 862.975 254.545 ;
        RECT 866.365 253.050 867.255 253.580 ;
        RECT 643.580 251.005 643.750 251.175 ;
        RECT 622.940 250.410 623.110 250.580 ;
        RECT 603.680 250.145 603.850 250.315 ;
        RECT 627.300 250.275 627.470 250.445 ;
        RECT 628.090 250.275 628.260 250.445 ;
        RECT 628.880 250.275 629.050 250.445 ;
        RECT 629.670 250.275 629.840 250.445 ;
        RECT 630.460 250.275 630.630 250.445 ;
        RECT 857.130 250.650 857.300 250.820 ;
        RECT 639.150 249.985 639.320 250.155 ;
        RECT 643.200 250.035 643.370 250.205 ;
        RECT 591.520 249.550 591.690 249.720 ;
        RECT 591.520 249.190 591.690 249.360 ;
        RECT 606.220 249.405 606.390 249.575 ;
        RECT 607.010 249.405 607.180 249.575 ;
        RECT 607.800 249.405 607.970 249.575 ;
        RECT 608.590 249.405 608.760 249.575 ;
        RECT 609.380 249.405 609.550 249.575 ;
        RECT 609.970 249.455 610.140 249.625 ;
        RECT 610.760 249.455 610.930 249.625 ;
        RECT 611.550 249.455 611.720 249.625 ;
        RECT 612.340 249.455 612.510 249.625 ;
        RECT 613.130 249.455 613.300 249.625 ;
        RECT 613.800 249.405 613.970 249.575 ;
        RECT 615.380 249.405 615.550 249.575 ;
        RECT 616.960 249.405 617.130 249.575 ;
        RECT 617.560 249.425 617.730 249.595 ;
        RECT 618.350 249.425 618.520 249.595 ;
        RECT 619.140 249.425 619.310 249.595 ;
        RECT 619.930 249.425 620.100 249.595 ;
        RECT 620.720 249.425 620.890 249.595 ;
        RECT 621.310 249.405 621.480 249.575 ;
        RECT 622.100 249.405 622.270 249.575 ;
        RECT 622.890 249.405 623.060 249.575 ;
        RECT 623.680 249.405 623.850 249.575 ;
        RECT 624.470 249.405 624.640 249.575 ;
        RECT 591.520 248.830 591.690 249.000 ;
        RECT 591.520 248.470 591.690 248.640 ;
        RECT 682.925 247.890 683.095 248.060 ;
        RECT 681.055 246.625 681.225 246.795 ;
        RECT 685.810 246.900 685.980 247.070 ;
        RECT 688.625 247.100 688.795 247.270 ;
        RECT 686.755 246.705 686.925 246.875 ;
        RECT 686.755 246.345 686.925 246.515 ;
        RECT 691.570 246.610 691.740 246.780 ;
        RECT 700.155 247.910 700.325 248.080 ;
        RECT 692.510 246.880 692.680 247.050 ;
        RECT 693.930 247.045 694.100 247.215 ;
        RECT 698.285 246.645 698.455 246.815 ;
        RECT 703.040 246.920 703.210 247.090 ;
        RECT 705.855 247.120 706.025 247.290 ;
        RECT 703.985 246.725 704.155 246.895 ;
        RECT 703.985 246.365 704.155 246.535 ;
        RECT 708.800 246.630 708.970 246.800 ;
        RECT 717.725 248.010 717.895 248.180 ;
        RECT 709.740 246.900 709.910 247.070 ;
        RECT 711.160 247.065 711.330 247.235 ;
        RECT 715.855 246.745 716.025 246.915 ;
        RECT 720.610 247.020 720.780 247.190 ;
        RECT 723.425 247.220 723.595 247.390 ;
        RECT 721.555 246.825 721.725 246.995 ;
        RECT 721.555 246.465 721.725 246.635 ;
        RECT 726.370 246.730 726.540 246.900 ;
        RECT 734.895 248.040 735.065 248.210 ;
        RECT 727.310 247.000 727.480 247.170 ;
        RECT 728.730 247.165 728.900 247.335 ;
        RECT 733.025 246.775 733.195 246.945 ;
        RECT 737.780 247.050 737.950 247.220 ;
        RECT 740.595 247.250 740.765 247.420 ;
        RECT 738.725 246.855 738.895 247.025 ;
        RECT 738.725 246.495 738.895 246.665 ;
        RECT 743.540 246.760 743.710 246.930 ;
        RECT 752.705 248.100 752.875 248.270 ;
        RECT 744.480 247.030 744.650 247.200 ;
        RECT 745.900 247.195 746.070 247.365 ;
        RECT 750.835 246.835 751.005 247.005 ;
        RECT 755.590 247.110 755.760 247.280 ;
        RECT 758.405 247.310 758.575 247.480 ;
        RECT 761.350 246.820 761.520 246.990 ;
        RECT 762.290 247.090 762.460 247.260 ;
        RECT 763.710 247.255 763.880 247.425 ;
        RECT 378.800 241.305 381.850 243.275 ;
        RECT 331.035 231.305 333.365 232.555 ;
        RECT 339.330 217.580 339.500 217.750 ;
        RECT 339.690 217.580 339.860 217.750 ;
        RECT 340.050 217.580 340.220 217.750 ;
        RECT 331.510 215.215 331.680 215.385 ;
        RECT 331.510 214.855 331.680 215.025 ;
        RECT 338.090 215.215 338.260 215.385 ;
        RECT 338.090 214.855 338.260 215.025 ;
        RECT 331.510 211.745 331.680 211.915 ;
        RECT 331.510 211.385 331.680 211.555 ;
        RECT 331.510 208.275 331.680 208.445 ;
        RECT 331.510 207.915 331.680 208.085 ;
        RECT 331.510 204.805 331.680 204.975 ;
        RECT 331.510 204.445 331.680 204.615 ;
        RECT 331.510 201.335 331.680 201.505 ;
        RECT 344.670 215.215 344.840 215.385 ;
        RECT 344.670 214.855 344.840 215.025 ;
        RECT 338.090 211.745 338.260 211.915 ;
        RECT 338.090 211.385 338.260 211.555 ;
        RECT 338.090 208.275 338.260 208.445 ;
        RECT 338.090 207.915 338.260 208.085 ;
        RECT 338.090 204.805 338.260 204.975 ;
        RECT 338.090 204.445 338.260 204.615 ;
        RECT 331.510 200.975 331.680 201.145 ;
        RECT 338.090 201.335 338.260 201.505 ;
        RECT 344.670 211.745 344.840 211.915 ;
        RECT 344.670 211.385 344.840 211.555 ;
        RECT 344.670 208.275 344.840 208.445 ;
        RECT 344.670 207.915 344.840 208.085 ;
        RECT 344.670 204.805 344.840 204.975 ;
        RECT 344.670 204.445 344.840 204.615 ;
        RECT 338.090 200.975 338.260 201.145 ;
        RECT 344.670 201.335 344.840 201.505 ;
        RECT 344.670 200.975 344.840 201.145 ;
        RECT 404.675 197.330 404.845 197.500 ;
        RECT 405.035 197.330 405.205 197.500 ;
        RECT 402.480 195.105 402.650 195.275 ;
        RECT 409.060 195.105 409.230 195.275 ;
        RECT 402.480 194.745 402.650 194.915 ;
        RECT 402.480 191.635 402.650 191.805 ;
        RECT 402.480 191.275 402.650 191.445 ;
        RECT 402.480 188.165 402.650 188.335 ;
        RECT 402.480 187.805 402.650 187.975 ;
        RECT 402.480 184.695 402.650 184.865 ;
        RECT 402.480 184.335 402.650 184.505 ;
        RECT 402.480 181.225 402.650 181.395 ;
        RECT 402.480 180.865 402.650 181.035 ;
        RECT 402.480 177.755 402.650 177.925 ;
        RECT 415.640 195.105 415.810 195.275 ;
        RECT 409.060 194.745 409.230 194.915 ;
        RECT 409.060 191.635 409.230 191.805 ;
        RECT 409.060 191.275 409.230 191.445 ;
        RECT 409.060 188.165 409.230 188.335 ;
        RECT 409.060 187.805 409.230 187.975 ;
        RECT 409.060 184.695 409.230 184.865 ;
        RECT 409.060 184.335 409.230 184.505 ;
        RECT 409.060 181.225 409.230 181.395 ;
        RECT 409.060 180.865 409.230 181.035 ;
        RECT 409.060 177.755 409.230 177.925 ;
        RECT 415.640 194.745 415.810 194.915 ;
        RECT 415.640 191.635 415.810 191.805 ;
        RECT 415.640 191.275 415.810 191.445 ;
        RECT 415.640 188.165 415.810 188.335 ;
        RECT 415.640 187.805 415.810 187.975 ;
        RECT 415.640 184.695 415.810 184.865 ;
        RECT 415.640 184.335 415.810 184.505 ;
        RECT 415.640 181.225 415.810 181.395 ;
        RECT 415.640 180.865 415.810 181.035 ;
        RECT 415.640 177.755 415.810 177.925 ;
        RECT 402.480 177.395 402.650 177.565 ;
        RECT 409.060 177.395 409.230 177.565 ;
        RECT 415.640 177.395 415.810 177.565 ;
      LAYER met1 ;
        RECT 379.270 369.180 379.500 370.160 ;
        RECT 385.850 369.520 386.080 370.160 ;
        RECT 385.520 367.560 386.150 369.520 ;
        RECT 385.510 367.400 386.150 367.560 ;
        RECT 385.510 367.230 386.010 367.400 ;
        RECT 379.130 364.610 379.360 365.590 ;
        RECT 385.520 365.260 386.010 367.230 ;
        RECT 385.650 365.250 386.010 365.260 ;
        RECT 385.710 364.610 385.940 365.250 ;
        RECT 379.130 361.140 379.360 362.120 ;
        RECT 385.710 361.140 385.940 362.120 ;
        RECT 379.130 357.670 379.360 358.650 ;
        RECT 385.710 357.670 385.940 358.650 ;
        RECT 379.130 354.200 379.360 355.180 ;
        RECT 385.710 354.200 385.940 355.180 ;
        RECT 838.950 353.130 839.420 353.660 ;
        RECT 662.925 352.955 663.215 353.000 ;
        RECT 668.205 352.955 668.495 353.000 ;
        RECT 670.605 352.955 670.895 353.000 ;
        RECT 662.925 352.815 670.895 352.955 ;
        RECT 672.010 352.930 672.370 352.990 ;
        RECT 652.870 352.730 653.450 352.790 ;
        RECT 662.925 352.770 663.215 352.815 ;
        RECT 668.205 352.770 668.495 352.815 ;
        RECT 670.605 352.770 670.895 352.815 ;
        RECT 652.850 352.150 653.470 352.730 ;
        RECT 671.940 352.380 672.420 352.930 ;
        RECT 680.975 352.915 681.265 352.960 ;
        RECT 686.255 352.915 686.545 352.960 ;
        RECT 688.655 352.915 688.945 352.960 ;
        RECT 680.975 352.775 688.945 352.915 ;
        RECT 698.565 352.935 698.855 352.980 ;
        RECT 703.845 352.935 704.135 352.980 ;
        RECT 706.245 352.935 706.535 352.980 ;
        RECT 690.100 352.830 690.390 352.840 ;
        RECT 680.975 352.730 681.265 352.775 ;
        RECT 686.255 352.730 686.545 352.775 ;
        RECT 688.655 352.730 688.945 352.775 ;
        RECT 672.010 352.350 672.370 352.380 ;
        RECT 690.050 352.340 690.440 352.830 ;
        RECT 698.565 352.795 706.535 352.935 ;
        RECT 698.565 352.750 698.855 352.795 ;
        RECT 703.845 352.750 704.135 352.795 ;
        RECT 706.245 352.750 706.535 352.795 ;
        RECT 707.630 352.450 708.030 353.010 ;
        RECT 716.415 352.935 716.705 352.980 ;
        RECT 721.695 352.935 721.985 352.980 ;
        RECT 724.095 352.935 724.385 352.980 ;
        RECT 716.415 352.795 724.385 352.935 ;
        RECT 725.510 352.890 725.850 352.950 ;
        RECT 734.675 352.935 734.965 352.980 ;
        RECT 739.955 352.935 740.245 352.980 ;
        RECT 742.355 352.935 742.645 352.980 ;
        RECT 716.415 352.750 716.705 352.795 ;
        RECT 721.695 352.750 721.985 352.795 ;
        RECT 724.095 352.750 724.385 352.795 ;
        RECT 725.490 352.380 725.870 352.890 ;
        RECT 734.675 352.795 742.645 352.935 ;
        RECT 743.770 352.920 744.130 352.980 ;
        RECT 734.675 352.750 734.965 352.795 ;
        RECT 739.955 352.750 740.245 352.795 ;
        RECT 742.355 352.750 742.645 352.795 ;
        RECT 743.750 352.460 744.150 352.920 ;
        RECT 752.445 352.905 752.735 352.950 ;
        RECT 757.725 352.905 758.015 352.950 ;
        RECT 760.125 352.905 760.415 352.950 ;
        RECT 752.445 352.765 760.415 352.905 ;
        RECT 752.445 352.720 752.735 352.765 ;
        RECT 757.725 352.720 758.015 352.765 ;
        RECT 760.125 352.720 760.415 352.765 ;
        RECT 743.770 352.400 744.130 352.460 ;
        RECT 761.470 352.430 761.970 352.930 ;
        RECT 770.485 352.825 770.775 352.870 ;
        RECT 775.765 352.825 776.055 352.870 ;
        RECT 778.165 352.825 778.455 352.870 ;
        RECT 788.645 352.865 788.935 352.910 ;
        RECT 793.925 352.865 794.215 352.910 ;
        RECT 796.325 352.865 796.615 352.910 ;
        RECT 770.485 352.685 778.455 352.825 ;
        RECT 779.550 352.800 779.900 352.860 ;
        RECT 770.485 352.640 770.775 352.685 ;
        RECT 775.765 352.640 776.055 352.685 ;
        RECT 778.165 352.640 778.455 352.685 ;
        RECT 779.530 352.430 779.920 352.800 ;
        RECT 788.645 352.725 796.615 352.865 ;
        RECT 797.700 352.860 798.080 352.920 ;
        RECT 807.025 352.875 807.315 352.920 ;
        RECT 812.305 352.875 812.595 352.920 ;
        RECT 814.705 352.875 814.995 352.920 ;
        RECT 788.645 352.680 788.935 352.725 ;
        RECT 793.925 352.680 794.215 352.725 ;
        RECT 796.325 352.680 796.615 352.725 ;
        RECT 797.680 352.490 798.100 352.860 ;
        RECT 807.025 352.735 814.995 352.875 ;
        RECT 816.100 352.860 816.440 352.920 ;
        RECT 807.025 352.690 807.315 352.735 ;
        RECT 812.305 352.690 812.595 352.735 ;
        RECT 814.705 352.690 814.995 352.735 ;
        RECT 816.080 352.540 816.460 352.860 ;
        RECT 825.825 352.855 826.115 352.900 ;
        RECT 831.105 352.855 831.395 352.900 ;
        RECT 833.505 352.855 833.795 352.900 ;
        RECT 825.825 352.715 833.795 352.855 ;
        RECT 825.825 352.670 826.115 352.715 ;
        RECT 831.105 352.670 831.395 352.715 ;
        RECT 833.505 352.670 833.795 352.715 ;
        RECT 834.940 352.790 835.240 352.900 ;
        RECT 836.230 352.790 836.500 352.800 ;
        RECT 834.940 352.580 836.520 352.790 ;
        RECT 797.700 352.430 798.080 352.490 ;
        RECT 816.100 352.480 816.440 352.540 ;
        RECT 834.940 352.520 835.240 352.580 ;
        RECT 725.510 352.320 725.850 352.380 ;
        RECT 779.550 352.370 779.900 352.430 ;
        RECT 652.870 352.090 653.450 352.150 ;
        RECT 669.170 352.040 669.460 352.220 ;
        RECT 675.750 352.040 676.040 352.140 ;
        RECT 669.170 351.790 676.040 352.040 ;
        RECT 669.170 351.720 669.460 351.790 ;
        RECT 379.130 350.730 379.360 351.710 ;
        RECT 385.710 351.080 385.940 351.710 ;
        RECT 675.750 351.640 676.040 351.790 ;
        RECT 687.270 352.060 687.560 352.220 ;
        RECT 693.360 352.060 693.650 352.220 ;
        RECT 687.270 351.830 693.650 352.060 ;
        RECT 687.270 351.720 687.560 351.830 ;
        RECT 693.360 351.720 693.650 351.830 ;
        RECT 704.800 352.060 705.120 352.240 ;
        RECT 711.160 352.060 711.480 352.170 ;
        RECT 704.800 351.820 711.480 352.060 ;
        RECT 704.800 351.760 705.120 351.820 ;
        RECT 711.160 351.690 711.480 351.820 ;
        RECT 722.680 351.990 723.000 352.160 ;
        RECT 729.430 351.990 729.750 352.140 ;
        RECT 722.680 351.780 729.750 351.990 ;
        RECT 722.680 351.680 723.000 351.780 ;
        RECT 729.430 351.660 729.750 351.780 ;
        RECT 740.910 352.040 741.260 352.250 ;
        RECT 747.180 352.040 747.530 352.160 ;
        RECT 740.910 351.770 747.530 352.040 ;
        RECT 740.910 351.730 741.260 351.770 ;
        RECT 747.180 351.640 747.530 351.770 ;
        RECT 758.630 351.850 759.080 351.870 ;
        RECT 758.630 351.840 759.790 351.850 ;
        RECT 765.210 351.840 765.560 352.040 ;
        RECT 758.630 351.630 765.560 351.840 ;
        RECT 776.730 351.870 777.030 352.130 ;
        RECT 783.410 351.870 783.710 352.010 ;
        RECT 776.730 351.660 783.710 351.870 ;
        RECT 776.730 351.650 777.030 351.660 ;
        RECT 758.630 351.580 759.080 351.630 ;
        RECT 765.210 351.520 765.560 351.630 ;
        RECT 783.410 351.530 783.710 351.660 ;
        RECT 794.880 351.850 795.180 352.020 ;
        RECT 801.790 351.850 802.090 352.030 ;
        RECT 794.880 351.680 802.090 351.850 ;
        RECT 794.880 351.540 795.180 351.680 ;
        RECT 801.790 351.550 802.090 351.680 ;
        RECT 813.270 351.890 813.590 352.050 ;
        RECT 818.480 351.890 819.590 352.370 ;
        RECT 820.590 351.890 820.910 351.970 ;
        RECT 813.270 351.690 820.910 351.890 ;
        RECT 813.270 351.600 813.590 351.690 ;
        RECT 818.480 351.580 819.590 351.690 ;
        RECT 820.590 351.520 820.910 351.690 ;
        RECT 828.850 351.660 829.440 352.030 ;
        RECT 836.230 351.900 836.500 352.580 ;
        RECT 836.050 351.260 836.830 351.900 ;
        RECT 379.110 345.730 379.340 346.710 ;
        RECT 385.630 346.350 386.050 351.080 ;
        RECT 656.030 350.290 656.720 350.350 ;
        RECT 656.010 349.530 656.740 350.290 ;
        RECT 656.030 349.470 656.720 349.530 ;
        RECT 784.360 348.860 785.070 349.280 ;
        RECT 832.050 348.000 834.190 349.500 ;
        RECT 837.260 347.110 839.140 348.580 ;
        RECT 845.660 347.760 847.180 348.420 ;
        RECT 870.570 347.760 871.970 348.010 ;
        RECT 845.660 347.080 871.970 347.760 ;
        RECT 845.660 346.990 847.180 347.080 ;
        RECT 385.690 345.730 385.920 346.350 ;
        RECT 870.570 345.630 871.970 347.080 ;
        RECT 787.730 345.580 792.710 345.610 ;
        RECT 787.650 345.560 813.510 345.580 ;
        RECT 787.650 345.290 813.740 345.560 ;
        RECT 787.650 345.270 792.710 345.290 ;
        RECT 780.090 344.730 781.030 344.790 ;
        RECT 780.070 343.390 781.050 344.730 ;
        RECT 785.740 343.960 786.110 344.040 ;
        RECT 787.650 343.960 787.950 345.270 ;
        RECT 813.260 345.200 813.740 345.290 ;
        RECT 799.225 344.785 799.515 344.830 ;
        RECT 804.505 344.785 804.795 344.830 ;
        RECT 806.905 344.785 807.195 344.830 ;
        RECT 799.225 344.645 807.195 344.785 ;
        RECT 799.225 344.600 799.515 344.645 ;
        RECT 804.505 344.600 804.795 344.645 ;
        RECT 806.905 344.600 807.195 344.645 ;
        RECT 818.585 344.695 818.875 344.740 ;
        RECT 823.865 344.695 824.155 344.740 ;
        RECT 826.265 344.695 826.555 344.740 ;
        RECT 818.585 344.555 826.555 344.695 ;
        RECT 818.585 344.510 818.875 344.555 ;
        RECT 823.865 344.510 824.155 344.555 ;
        RECT 826.265 344.510 826.555 344.555 ;
        RECT 785.740 343.700 787.950 343.960 ;
        RECT 805.440 343.920 805.780 344.110 ;
        RECT 813.350 343.920 813.690 344.000 ;
        RECT 785.740 343.540 786.110 343.700 ;
        RECT 805.440 343.680 813.690 343.920 ;
        RECT 805.600 343.660 813.690 343.680 ;
        RECT 813.350 343.570 813.690 343.660 ;
        RECT 824.800 343.480 825.220 344.020 ;
        RECT 824.830 343.470 825.160 343.480 ;
        RECT 780.090 343.330 781.030 343.390 ;
        RECT 379.110 342.260 379.340 343.240 ;
        RECT 385.690 342.260 385.920 343.240 ;
        RECT 379.110 338.790 379.340 339.770 ;
        RECT 385.690 338.790 385.920 339.770 ;
        RECT 853.410 339.160 854.490 339.280 ;
        RECT 855.580 339.160 856.530 339.450 ;
        RECT 831.180 336.930 834.990 338.990 ;
        RECT 853.410 338.830 856.530 339.160 ;
        RECT 853.410 338.540 854.490 338.830 ;
        RECT 855.580 338.680 856.530 338.830 ;
        RECT 852.560 338.190 855.470 338.260 ;
        RECT 851.220 337.940 851.840 338.090 ;
        RECT 852.550 338.080 855.470 338.190 ;
        RECT 852.550 337.940 852.800 338.080 ;
        RECT 851.220 337.920 852.800 337.940 ;
        RECT 855.140 337.920 855.370 338.080 ;
        RECT 851.220 337.740 852.820 337.920 ;
        RECT 851.220 337.550 852.830 337.740 ;
        RECT 855.140 337.710 855.400 337.920 ;
        RECT 851.220 337.470 851.840 337.550 ;
        RECT 379.110 335.320 379.340 336.300 ;
        RECT 385.690 335.320 385.920 336.300 ;
        RECT 632.020 333.330 633.420 334.450 ;
        RECT 660.440 333.180 680.860 333.670 ;
        RECT 379.110 331.850 379.340 332.830 ;
        RECT 385.690 332.280 385.920 332.830 ;
        RECT 194.190 325.630 199.920 329.410 ;
        RECT 379.110 326.880 379.340 327.860 ;
        RECT 385.510 327.290 386.130 332.280 ;
        RECT 603.390 332.070 603.620 332.450 ;
        RECT 604.970 332.070 605.200 332.450 ;
        RECT 607.910 332.080 608.140 332.460 ;
        RECT 609.490 332.080 609.720 332.460 ;
        RECT 612.430 332.080 612.660 332.460 ;
        RECT 614.010 332.080 614.240 332.460 ;
        RECT 603.410 330.980 603.590 332.070 ;
        RECT 604.980 330.980 605.160 332.070 ;
        RECT 607.930 330.990 608.110 332.080 ;
        RECT 609.500 330.990 609.680 332.080 ;
        RECT 612.450 330.990 612.630 332.080 ;
        RECT 614.020 330.990 614.200 332.080 ;
        RECT 616.860 332.060 617.090 332.440 ;
        RECT 618.440 332.060 618.670 332.440 ;
        RECT 621.240 332.070 621.470 332.450 ;
        RECT 622.820 332.070 623.050 332.450 ;
        RECT 603.390 330.820 603.620 330.980 ;
        RECT 603.340 330.460 603.620 330.820 ;
        RECT 604.970 330.600 605.200 330.980 ;
        RECT 607.910 330.610 608.140 330.990 ;
        RECT 609.490 330.610 609.720 330.990 ;
        RECT 612.430 330.610 612.660 330.990 ;
        RECT 614.010 330.610 614.240 330.990 ;
        RECT 616.880 330.970 617.060 332.060 ;
        RECT 618.450 330.970 618.630 332.060 ;
        RECT 621.260 330.980 621.440 332.070 ;
        RECT 622.830 330.980 623.010 332.070 ;
        RECT 625.560 332.060 625.790 332.440 ;
        RECT 627.140 332.060 627.370 332.440 ;
        RECT 605.000 330.460 605.180 330.600 ;
        RECT 607.930 330.470 608.130 330.610 ;
        RECT 609.520 330.470 609.700 330.610 ;
        RECT 612.450 330.470 612.630 330.610 ;
        RECT 614.040 330.470 614.220 330.610 ;
        RECT 616.860 330.590 617.090 330.970 ;
        RECT 618.440 330.590 618.670 330.970 ;
        RECT 621.240 330.600 621.470 330.980 ;
        RECT 622.820 330.600 623.050 330.980 ;
        RECT 625.580 330.970 625.760 332.060 ;
        RECT 627.150 330.970 627.330 332.060 ;
        RECT 603.340 330.300 605.210 330.460 ;
        RECT 607.890 330.450 609.730 330.470 ;
        RECT 612.410 330.450 614.250 330.470 ;
        RECT 616.880 330.450 617.060 330.590 ;
        RECT 618.470 330.450 618.650 330.590 ;
        RECT 621.260 330.460 621.440 330.600 ;
        RECT 622.850 330.460 623.030 330.600 ;
        RECT 625.560 330.590 625.790 330.970 ;
        RECT 627.140 330.590 627.370 330.970 ;
        RECT 621.220 330.450 623.060 330.460 ;
        RECT 625.580 330.450 625.760 330.590 ;
        RECT 627.170 330.450 627.350 330.590 ;
        RECT 607.890 330.380 615.570 330.450 ;
        RECT 607.890 330.310 615.580 330.380 ;
        RECT 603.340 328.940 603.620 330.300 ;
        RECT 607.960 329.290 608.130 330.310 ;
        RECT 613.930 330.290 615.580 330.310 ;
        RECT 616.840 330.310 623.060 330.450 ;
        RECT 616.840 330.290 618.680 330.310 ;
        RECT 621.220 330.300 623.060 330.310 ;
        RECT 613.510 329.630 613.980 330.010 ;
        RECT 615.370 329.840 615.580 330.290 ;
        RECT 616.350 329.840 616.780 329.910 ;
        RECT 615.370 329.660 616.780 329.840 ;
        RECT 608.550 329.290 609.220 329.600 ;
        RECT 607.950 329.010 609.220 329.290 ;
        RECT 597.120 328.710 597.810 328.770 ;
        RECT 594.410 328.210 595.210 328.670 ;
        RECT 385.690 326.880 385.920 327.290 ;
        RECT 594.550 326.690 594.830 328.210 ;
        RECT 597.100 327.860 597.830 328.710 ;
        RECT 597.120 327.800 597.810 327.860 ;
        RECT 594.310 326.420 595.040 326.690 ;
        RECT 603.330 326.670 603.640 328.940 ;
        RECT 607.960 328.640 608.130 329.010 ;
        RECT 608.550 328.750 609.220 329.010 ;
        RECT 613.600 329.110 613.840 329.630 ;
        RECT 616.350 329.590 616.780 329.660 ;
        RECT 617.160 329.110 617.340 330.290 ;
        RECT 620.760 329.890 621.170 330.160 ;
        RECT 620.710 329.730 621.170 329.890 ;
        RECT 620.710 329.590 621.130 329.730 ;
        RECT 613.600 328.950 617.350 329.110 ;
        RECT 607.220 328.000 608.130 328.640 ;
        RECT 615.640 328.220 615.860 328.280 ;
        RECT 620.710 328.220 620.980 329.590 ;
        RECT 603.930 326.670 604.890 326.840 ;
        RECT 603.270 326.390 604.890 326.670 ;
        RECT 603.330 325.770 603.640 326.390 ;
        RECT 603.930 326.280 604.890 326.390 ;
        RECT 196.430 321.460 197.360 325.630 ;
        RECT 600.940 325.610 604.320 325.770 ;
        RECT 600.950 325.440 601.120 325.610 ;
        RECT 602.520 325.440 602.690 325.610 ;
        RECT 604.120 325.440 604.290 325.610 ;
        RECT 600.920 325.060 601.150 325.440 ;
        RECT 601.710 325.060 601.940 325.440 ;
        RECT 602.500 325.060 602.730 325.440 ;
        RECT 603.290 325.060 603.520 325.440 ;
        RECT 604.080 325.060 604.310 325.440 ;
        RECT 379.110 323.410 379.340 324.390 ;
        RECT 385.690 323.410 385.920 324.390 ;
        RECT 600.950 323.970 601.130 325.060 ;
        RECT 601.730 323.970 601.910 325.060 ;
        RECT 602.520 323.970 602.700 325.060 ;
        RECT 603.300 323.970 603.480 325.060 ;
        RECT 604.090 323.970 604.270 325.060 ;
        RECT 600.920 323.590 601.150 323.970 ;
        RECT 601.710 323.590 601.940 323.970 ;
        RECT 602.500 323.590 602.730 323.970 ;
        RECT 603.290 323.590 603.520 323.970 ;
        RECT 604.080 323.590 604.310 323.970 ;
        RECT 601.730 323.450 601.910 323.590 ;
        RECT 603.320 323.450 603.500 323.590 ;
        RECT 607.960 323.540 608.130 328.000 ;
        RECT 608.530 327.740 609.170 328.160 ;
        RECT 615.640 327.990 620.980 328.220 ;
        RECT 621.210 328.030 621.720 328.080 ;
        RECT 621.880 328.070 622.090 330.300 ;
        RECT 625.540 330.290 627.380 330.450 ;
        RECT 623.080 329.030 623.930 329.470 ;
        RECT 626.540 329.090 626.760 330.290 ;
        RECT 639.370 329.210 639.800 329.270 ;
        RECT 629.630 329.090 629.860 329.110 ;
        RECT 622.260 328.070 622.950 328.160 ;
        RECT 621.880 328.030 622.950 328.070 ;
        RECT 608.700 324.190 608.960 327.740 ;
        RECT 609.500 326.570 610.150 326.790 ;
        RECT 609.500 326.540 610.650 326.570 ;
        RECT 609.500 326.390 613.780 326.540 ;
        RECT 609.500 326.220 610.650 326.390 ;
        RECT 611.950 326.220 612.170 326.390 ;
        RECT 613.550 326.220 613.770 326.390 ;
        RECT 610.370 326.060 610.610 326.220 ;
        RECT 610.370 325.840 610.600 326.060 ;
        RECT 611.160 325.840 611.390 326.220 ;
        RECT 611.950 325.840 612.180 326.220 ;
        RECT 612.740 325.840 612.970 326.220 ;
        RECT 613.530 326.050 613.770 326.220 ;
        RECT 613.530 325.840 613.760 326.050 ;
        RECT 610.380 324.750 610.560 325.840 ;
        RECT 611.180 324.750 611.360 325.840 ;
        RECT 611.980 324.750 612.160 325.840 ;
        RECT 612.760 324.750 612.940 325.840 ;
        RECT 613.540 324.750 613.720 325.840 ;
        RECT 615.640 325.730 615.860 327.990 ;
        RECT 621.210 327.890 622.950 328.030 ;
        RECT 621.210 327.790 621.720 327.890 ;
        RECT 621.880 327.780 622.950 327.890 ;
        RECT 621.190 326.510 621.670 326.580 ;
        RECT 617.960 326.360 621.670 326.510 ;
        RECT 617.980 326.190 618.200 326.360 ;
        RECT 619.540 326.190 619.760 326.360 ;
        RECT 621.140 326.300 621.670 326.360 ;
        RECT 621.140 326.190 621.360 326.300 ;
        RECT 617.960 326.030 618.200 326.190 ;
        RECT 617.960 325.810 618.190 326.030 ;
        RECT 618.750 325.810 618.980 326.190 ;
        RECT 619.540 325.810 619.770 326.190 ;
        RECT 620.330 325.810 620.560 326.190 ;
        RECT 621.120 326.020 621.360 326.190 ;
        RECT 621.120 325.810 621.350 326.020 ;
        RECT 615.510 325.310 615.990 325.730 ;
        RECT 614.200 324.860 617.620 325.000 ;
        RECT 610.370 324.370 610.600 324.750 ;
        RECT 611.160 324.370 611.390 324.750 ;
        RECT 611.950 324.370 612.180 324.750 ;
        RECT 612.740 324.370 612.970 324.750 ;
        RECT 613.530 324.370 613.760 324.750 ;
        RECT 614.230 324.700 614.420 324.860 ;
        RECT 615.790 324.700 615.980 324.860 ;
        RECT 617.400 324.700 617.590 324.860 ;
        RECT 617.970 324.720 618.150 325.810 ;
        RECT 618.770 324.720 618.950 325.810 ;
        RECT 619.570 324.720 619.750 325.810 ;
        RECT 620.350 324.720 620.530 325.810 ;
        RECT 621.130 324.720 621.310 325.810 ;
        RECT 608.520 323.880 609.190 324.190 ;
        RECT 609.790 323.540 609.940 323.550 ;
        RECT 601.690 323.290 603.530 323.450 ;
        RECT 606.600 323.400 610.030 323.540 ;
        RECT 603.370 322.640 603.520 323.290 ;
        RECT 606.640 323.230 606.790 323.400 ;
        RECT 608.230 323.230 608.380 323.400 ;
        RECT 609.790 323.230 609.940 323.400 ;
        RECT 610.380 323.280 610.560 324.370 ;
        RECT 611.180 323.280 611.360 324.370 ;
        RECT 611.980 323.280 612.160 324.370 ;
        RECT 612.760 323.280 612.940 324.370 ;
        RECT 613.540 323.280 613.720 324.370 ;
        RECT 614.200 324.320 614.430 324.700 ;
        RECT 615.780 324.320 616.010 324.700 ;
        RECT 617.360 324.320 617.590 324.700 ;
        RECT 617.960 324.340 618.190 324.720 ;
        RECT 618.750 324.340 618.980 324.720 ;
        RECT 619.540 324.340 619.770 324.720 ;
        RECT 620.330 324.340 620.560 324.720 ;
        RECT 621.120 324.340 621.350 324.720 ;
        RECT 606.620 322.850 606.850 323.230 ;
        RECT 607.410 322.850 607.640 323.230 ;
        RECT 608.200 322.850 608.430 323.230 ;
        RECT 608.990 322.850 609.220 323.230 ;
        RECT 609.780 322.850 610.010 323.230 ;
        RECT 610.370 322.900 610.600 323.280 ;
        RECT 611.160 323.110 611.390 323.280 ;
        RECT 611.150 322.900 611.390 323.110 ;
        RECT 611.950 322.900 612.180 323.280 ;
        RECT 612.740 322.900 612.970 323.280 ;
        RECT 613.530 322.900 613.760 323.280 ;
        RECT 614.220 323.230 614.380 324.320 ;
        RECT 615.800 323.230 615.960 324.320 ;
        RECT 617.380 323.230 617.540 324.320 ;
        RECT 617.970 323.250 618.150 324.340 ;
        RECT 618.770 323.250 618.950 324.340 ;
        RECT 619.570 323.250 619.750 324.340 ;
        RECT 620.350 323.250 620.530 324.340 ;
        RECT 621.130 323.250 621.310 324.340 ;
        RECT 621.880 323.540 622.090 327.780 ;
        RECT 622.260 327.700 622.950 327.780 ;
        RECT 623.310 324.320 623.540 329.030 ;
        RECT 626.540 328.940 629.870 329.090 ;
        RECT 629.630 326.630 629.860 328.940 ;
        RECT 639.350 328.760 639.820 329.210 ;
        RECT 645.430 328.980 645.800 329.040 ;
        RECT 639.370 328.700 639.800 328.760 ;
        RECT 645.410 328.630 645.820 328.980 ;
        RECT 645.430 328.570 645.800 328.630 ;
        RECT 631.640 327.530 632.470 327.630 ;
        RECT 631.630 326.990 632.470 327.530 ;
        RECT 633.960 327.510 634.790 328.250 ;
        RECT 641.820 328.170 642.320 328.550 ;
        RECT 657.670 327.620 658.170 327.990 ;
        RECT 631.640 326.950 632.470 326.990 ;
        RECT 629.260 326.280 629.860 326.630 ;
        RECT 629.630 325.900 629.860 326.280 ;
        RECT 639.260 326.110 639.960 326.470 ;
        RECT 627.720 325.740 631.100 325.900 ;
        RECT 627.730 325.570 627.900 325.740 ;
        RECT 629.300 325.570 629.470 325.740 ;
        RECT 629.630 325.730 629.860 325.740 ;
        RECT 630.900 325.570 631.070 325.740 ;
        RECT 627.700 325.190 627.930 325.570 ;
        RECT 628.490 325.190 628.720 325.570 ;
        RECT 629.280 325.190 629.510 325.570 ;
        RECT 630.070 325.190 630.300 325.570 ;
        RECT 630.860 325.190 631.090 325.570 ;
        RECT 623.110 323.770 623.800 324.320 ;
        RECT 627.730 324.100 627.910 325.190 ;
        RECT 628.510 324.100 628.690 325.190 ;
        RECT 629.300 324.100 629.480 325.190 ;
        RECT 630.080 324.100 630.260 325.190 ;
        RECT 630.870 324.100 631.050 325.190 ;
        RECT 627.700 323.720 627.930 324.100 ;
        RECT 628.490 323.720 628.720 324.100 ;
        RECT 629.280 323.720 629.510 324.100 ;
        RECT 630.070 323.720 630.300 324.100 ;
        RECT 630.860 323.720 631.090 324.100 ;
        RECT 639.520 323.810 639.700 326.110 ;
        RECT 643.360 325.990 643.930 326.670 ;
        RECT 639.840 324.210 640.290 324.900 ;
        RECT 643.590 323.860 643.730 325.990 ;
        RECT 643.900 324.750 644.320 324.950 ;
        RECT 645.330 324.750 646.310 325.060 ;
        RECT 643.900 324.540 646.310 324.750 ;
        RECT 643.900 324.270 644.320 324.540 ;
        RECT 645.330 324.280 646.310 324.540 ;
        RECT 657.860 324.330 658.050 327.620 ;
        RECT 628.510 323.580 628.690 323.720 ;
        RECT 630.100 323.580 630.280 323.720 ;
        RECT 639.520 323.700 639.780 323.810 ;
        RECT 624.880 323.540 625.030 323.550 ;
        RECT 621.690 323.400 625.120 323.540 ;
        RECT 628.470 323.420 630.310 323.580 ;
        RECT 639.550 323.430 639.780 323.700 ;
        RECT 643.590 323.690 643.830 323.860 ;
        RECT 643.600 323.480 643.830 323.690 ;
        RECT 657.550 323.500 658.320 324.330 ;
        RECT 660.440 324.100 660.950 333.180 ;
        RECT 666.170 331.150 666.510 331.220 ;
        RECT 673.410 331.150 673.580 331.170 ;
        RECT 666.170 330.940 673.580 331.150 ;
        RECT 666.170 330.790 666.510 330.940 ;
        RECT 663.330 330.100 663.670 330.160 ;
        RECT 668.880 330.130 669.220 330.190 ;
        RECT 673.410 330.170 673.580 330.940 ;
        RECT 680.650 330.850 680.860 333.180 ;
        RECT 682.220 330.850 682.810 330.910 ;
        RECT 680.650 330.630 682.810 330.850 ;
        RECT 682.220 330.620 682.810 330.630 ;
        RECT 686.880 330.480 687.140 330.530 ;
        RECT 677.580 330.340 687.140 330.480 ;
        RECT 677.580 330.220 688.680 330.340 ;
        RECT 673.410 330.140 676.360 330.170 ;
        RECT 663.310 329.740 663.690 330.100 ;
        RECT 664.270 329.780 664.640 329.840 ;
        RECT 663.330 329.680 663.670 329.740 ;
        RECT 664.250 329.440 664.660 329.780 ;
        RECT 668.860 329.720 669.240 330.130 ;
        RECT 673.410 330.030 676.440 330.140 ;
        RECT 669.890 329.890 670.250 329.950 ;
        RECT 668.880 329.660 669.220 329.720 ;
        RECT 669.870 329.440 670.270 329.890 ;
        RECT 676.100 329.710 676.440 330.030 ;
        RECT 677.580 329.990 677.860 330.220 ;
        RECT 686.880 330.130 688.680 330.220 ;
        RECT 686.880 330.030 688.890 330.130 ;
        RECT 682.210 329.970 682.580 330.030 ;
        RECT 686.880 330.010 687.140 330.030 ;
        RECT 682.190 329.520 682.600 329.970 ;
        RECT 683.100 329.770 683.580 329.830 ;
        RECT 682.210 329.460 682.580 329.520 ;
        RECT 664.270 329.380 664.640 329.440 ;
        RECT 669.890 329.380 670.250 329.440 ;
        RECT 683.080 329.320 683.600 329.770 ;
        RECT 688.540 329.670 688.890 330.030 ;
        RECT 832.380 329.960 833.290 336.930 ;
        RECT 832.340 329.320 833.290 329.960 ;
        RECT 683.100 329.260 683.580 329.320 ;
        RECT 778.390 328.170 780.000 328.380 ;
        RECT 832.340 328.170 833.270 329.320 ;
        RECT 662.510 327.500 675.640 327.510 ;
        RECT 662.450 327.370 675.670 327.500 ;
        RECT 662.450 324.270 662.650 327.370 ;
        RECT 663.320 327.020 663.780 327.370 ;
        RECT 664.320 327.070 664.880 327.160 ;
        RECT 664.320 327.040 667.500 327.070 ;
        RECT 664.320 326.800 675.290 327.040 ;
        RECT 664.570 326.780 675.290 326.800 ;
        RECT 664.570 326.760 667.500 326.780 ;
        RECT 667.180 324.270 667.340 326.760 ;
        RECT 660.220 323.510 660.970 324.100 ;
        RECT 662.280 323.600 663.220 324.270 ;
        RECT 665.480 324.110 666.020 324.140 ;
        RECT 607.450 322.700 607.600 322.850 ;
        RECT 609.030 322.700 609.180 322.850 ;
        RECT 610.410 322.700 610.590 322.900 ;
        RECT 208.860 321.460 210.530 321.860 ;
        RECT 196.430 320.810 210.530 321.460 ;
        RECT 591.880 321.280 592.130 322.445 ;
        RECT 602.290 322.230 603.070 322.260 ;
        RECT 602.280 321.890 603.070 322.230 ;
        RECT 603.290 322.200 603.740 322.640 ;
        RECT 607.400 322.550 610.590 322.700 ;
        RECT 611.150 322.740 611.320 322.900 ;
        RECT 612.750 322.740 612.920 322.900 ;
        RECT 614.200 322.850 614.430 323.230 ;
        RECT 615.780 322.850 616.010 323.230 ;
        RECT 617.360 322.850 617.590 323.230 ;
        RECT 617.960 322.870 618.190 323.250 ;
        RECT 618.750 323.080 618.980 323.250 ;
        RECT 618.740 322.870 618.980 323.080 ;
        RECT 619.540 322.870 619.770 323.250 ;
        RECT 620.330 322.870 620.560 323.250 ;
        RECT 621.120 323.070 621.350 323.250 ;
        RECT 621.730 323.230 621.880 323.400 ;
        RECT 623.320 323.230 623.470 323.400 ;
        RECT 624.880 323.230 625.030 323.400 ;
        RECT 621.120 322.870 621.360 323.070 ;
        RECT 614.200 322.740 614.400 322.850 ;
        RECT 611.150 322.630 614.400 322.740 ;
        RECT 609.170 322.520 610.590 322.550 ;
        RECT 611.090 322.600 614.400 322.630 ;
        RECT 611.090 322.590 612.990 322.600 ;
        RECT 611.090 322.290 611.500 322.590 ;
        RECT 614.200 322.230 614.400 322.600 ;
        RECT 617.370 322.700 617.590 322.850 ;
        RECT 618.740 322.710 618.910 322.870 ;
        RECT 620.340 322.710 620.510 322.870 ;
        RECT 618.740 322.700 620.580 322.710 ;
        RECT 617.370 322.620 620.580 322.700 ;
        RECT 621.160 322.660 621.360 322.870 ;
        RECT 621.710 322.850 621.940 323.230 ;
        RECT 622.500 322.850 622.730 323.230 ;
        RECT 623.290 322.850 623.520 323.230 ;
        RECT 624.080 322.850 624.310 323.230 ;
        RECT 624.870 322.850 625.100 323.230 ;
        RECT 622.540 322.700 622.690 322.850 ;
        RECT 624.120 322.700 624.270 322.850 ;
        RECT 622.490 322.660 624.310 322.700 ;
        RECT 617.370 322.560 620.620 322.620 ;
        RECT 617.370 322.530 619.130 322.560 ;
        RECT 620.220 322.260 620.620 322.560 ;
        RECT 621.160 322.550 624.310 322.660 ;
        RECT 621.160 322.500 622.650 322.550 ;
        RECT 629.210 322.070 629.420 323.420 ;
        RECT 602.280 321.870 602.960 321.890 ;
        RECT 629.040 321.720 629.660 322.070 ;
        RECT 208.860 320.380 210.530 320.810 ;
        RECT 379.110 319.940 379.340 320.920 ;
        RECT 385.690 319.940 385.920 320.920 ;
        RECT 591.290 319.970 592.660 321.280 ;
        RECT 211.890 319.290 212.870 319.520 ;
        RECT 215.360 319.290 216.340 319.520 ;
        RECT 218.830 319.290 219.810 319.520 ;
        RECT 222.300 319.290 223.280 319.520 ;
        RECT 225.770 319.290 226.750 319.520 ;
        RECT 231.930 319.280 232.910 319.510 ;
        RECT 235.400 319.280 236.380 319.510 ;
        RECT 238.870 319.280 239.850 319.510 ;
        RECT 242.340 319.280 243.320 319.510 ;
        RECT 245.810 319.280 246.790 319.510 ;
        RECT 251.990 319.280 252.970 319.510 ;
        RECT 255.460 319.280 256.440 319.510 ;
        RECT 258.930 319.280 259.910 319.510 ;
        RECT 262.400 319.280 263.380 319.510 ;
        RECT 265.870 319.280 266.850 319.510 ;
        RECT 272.040 319.280 273.020 319.510 ;
        RECT 275.510 319.280 276.490 319.510 ;
        RECT 278.980 319.280 279.960 319.510 ;
        RECT 282.450 319.280 283.430 319.510 ;
        RECT 285.920 319.280 286.900 319.510 ;
        RECT 660.360 318.760 660.710 323.510 ;
        RECT 665.420 323.390 666.070 324.110 ;
        RECT 667.010 323.700 667.960 324.270 ;
        RECT 669.960 324.220 670.600 324.280 ;
        RECT 665.480 323.360 666.020 323.390 ;
        RECT 669.210 323.370 669.660 323.920 ;
        RECT 669.940 323.620 670.620 324.220 ;
        RECT 671.670 324.120 672.200 324.180 ;
        RECT 669.960 323.560 670.600 323.620 ;
        RECT 671.650 323.560 672.220 324.120 ;
        RECT 675.150 323.740 675.290 326.780 ;
        RECT 675.530 324.640 675.670 327.370 ;
        RECT 778.020 326.980 833.270 328.170 ;
        RECT 778.020 326.920 833.050 326.980 ;
        RECT 679.610 325.050 679.930 325.180 ;
        RECT 686.230 325.050 686.470 325.080 ;
        RECT 679.610 324.890 686.470 325.050 ;
        RECT 677.390 324.640 677.660 324.690 ;
        RECT 675.530 324.430 677.660 324.640 ;
        RECT 679.610 324.590 679.930 324.890 ;
        RECT 677.390 324.350 677.660 324.430 ;
        RECT 675.150 323.730 676.450 323.740 ;
        RECT 676.840 323.730 677.110 323.830 ;
        RECT 671.670 323.500 672.200 323.560 ;
        RECT 664.770 319.190 665.100 319.250 ;
        RECT 662.010 318.760 662.440 318.820 ;
        RECT 660.360 318.480 662.440 318.760 ;
        RECT 664.750 318.680 665.120 319.190 ;
        RECT 664.770 318.620 665.100 318.680 ;
        RECT 660.360 318.470 662.170 318.480 ;
        RECT 665.630 318.190 665.860 323.360 ;
        RECT 669.310 323.300 669.580 323.370 ;
        RECT 673.720 323.360 674.170 323.710 ;
        RECT 675.150 323.570 677.110 323.730 ;
        RECT 675.680 323.560 677.110 323.570 ;
        RECT 676.840 323.490 677.110 323.560 ;
        RECT 678.090 323.020 678.540 323.430 ;
        RECT 682.020 323.420 682.630 324.120 ;
        RECT 683.020 323.180 683.530 323.740 ;
        RECT 686.230 323.350 686.470 324.890 ;
        RECT 688.570 323.350 688.880 323.490 ;
        RECT 683.080 323.020 683.440 323.180 ;
        RECT 686.230 323.090 688.880 323.350 ;
        RECT 678.160 322.980 678.430 323.020 ;
        RECT 688.570 322.990 688.880 323.090 ;
        RECT 670.170 319.330 670.510 319.420 ;
        RECT 670.170 319.130 677.200 319.330 ;
        RECT 670.170 318.980 670.510 319.130 ;
        RECT 662.080 317.960 665.860 318.190 ;
        RECT 667.360 318.410 667.700 318.450 ;
        RECT 671.290 318.410 671.800 318.550 ;
        RECT 667.360 318.220 673.130 318.410 ;
        RECT 667.360 318.000 667.700 318.220 ;
        RECT 671.290 318.070 671.800 318.220 ;
        RECT 672.790 317.960 673.130 318.220 ;
        RECT 677.040 318.070 677.200 319.130 ;
        RECT 691.840 318.110 692.190 318.260 ;
        RECT 692.530 318.110 692.740 318.670 ;
        RECT 694.160 318.110 694.450 318.290 ;
        RECT 677.040 318.050 679.610 318.070 ;
        RECT 673.740 317.990 674.060 318.020 ;
        RECT 661.940 317.920 665.860 317.960 ;
        RECT 661.940 317.890 665.790 317.920 ;
        RECT 661.940 317.620 662.370 317.890 ;
        RECT 668.250 317.540 668.650 317.960 ;
        RECT 673.720 317.600 674.100 317.990 ;
        RECT 677.040 317.950 679.850 318.050 ;
        RECT 677.090 317.930 679.850 317.950 ;
        RECT 679.490 317.760 679.850 317.930 ;
        RECT 691.840 317.910 694.450 318.110 ;
        RECT 691.840 317.890 694.330 317.910 ;
        RECT 691.840 317.790 693.080 317.890 ;
        RECT 684.410 317.620 684.730 317.680 ;
        RECT 673.740 317.590 674.060 317.600 ;
        RECT 379.110 316.470 379.340 317.450 ;
        RECT 385.690 316.470 385.920 317.450 ;
        RECT 662.800 317.120 663.350 317.540 ;
        RECT 684.390 317.180 684.750 317.620 ;
        RECT 692.270 317.400 693.080 317.790 ;
        RECT 684.410 317.120 684.730 317.180 ;
        RECT 632.390 315.440 633.540 316.340 ;
        RECT 379.110 313.000 379.340 313.980 ;
        RECT 385.690 313.780 385.920 313.980 ;
        RECT 603.240 313.900 603.470 314.280 ;
        RECT 604.820 313.900 605.050 314.280 ;
        RECT 607.760 313.910 607.990 314.290 ;
        RECT 609.340 313.910 609.570 314.290 ;
        RECT 612.280 313.910 612.510 314.290 ;
        RECT 613.860 313.910 614.090 314.290 ;
        RECT 211.890 312.710 212.870 312.940 ;
        RECT 215.360 312.710 216.340 312.940 ;
        RECT 218.830 312.710 219.810 312.940 ;
        RECT 222.300 312.710 223.280 312.940 ;
        RECT 225.770 312.710 226.750 312.940 ;
        RECT 231.930 312.700 232.910 312.930 ;
        RECT 235.400 312.700 236.380 312.930 ;
        RECT 238.870 312.700 239.850 312.930 ;
        RECT 242.340 312.700 243.320 312.930 ;
        RECT 245.810 312.700 246.790 312.930 ;
        RECT 251.990 312.700 252.970 312.930 ;
        RECT 255.460 312.700 256.440 312.930 ;
        RECT 258.930 312.700 259.910 312.930 ;
        RECT 262.400 312.700 263.380 312.930 ;
        RECT 265.870 312.700 266.850 312.930 ;
        RECT 272.040 312.700 273.020 312.930 ;
        RECT 275.510 312.700 276.490 312.930 ;
        RECT 278.980 312.700 279.960 312.930 ;
        RECT 282.450 312.700 283.430 312.930 ;
        RECT 285.920 312.700 286.900 312.930 ;
        RECT 379.110 308.060 379.340 309.040 ;
        RECT 385.620 308.440 386.000 313.780 ;
        RECT 603.260 312.810 603.440 313.900 ;
        RECT 604.830 312.810 605.010 313.900 ;
        RECT 607.780 312.820 607.960 313.910 ;
        RECT 609.350 312.820 609.530 313.910 ;
        RECT 612.300 312.820 612.480 313.910 ;
        RECT 613.870 312.820 614.050 313.910 ;
        RECT 616.710 313.890 616.940 314.270 ;
        RECT 618.290 313.890 618.520 314.270 ;
        RECT 621.090 313.900 621.320 314.280 ;
        RECT 622.670 313.900 622.900 314.280 ;
        RECT 603.240 312.650 603.470 312.810 ;
        RECT 603.190 312.290 603.470 312.650 ;
        RECT 604.820 312.430 605.050 312.810 ;
        RECT 607.760 312.440 607.990 312.820 ;
        RECT 609.340 312.440 609.570 312.820 ;
        RECT 612.280 312.440 612.510 312.820 ;
        RECT 613.860 312.440 614.090 312.820 ;
        RECT 616.730 312.800 616.910 313.890 ;
        RECT 618.300 312.800 618.480 313.890 ;
        RECT 621.110 312.810 621.290 313.900 ;
        RECT 622.680 312.810 622.860 313.900 ;
        RECT 625.410 313.890 625.640 314.270 ;
        RECT 626.990 313.890 627.220 314.270 ;
        RECT 604.850 312.290 605.030 312.430 ;
        RECT 607.780 312.300 607.980 312.440 ;
        RECT 609.370 312.300 609.550 312.440 ;
        RECT 612.300 312.300 612.480 312.440 ;
        RECT 613.890 312.300 614.070 312.440 ;
        RECT 616.710 312.420 616.940 312.800 ;
        RECT 618.290 312.420 618.520 312.800 ;
        RECT 621.090 312.430 621.320 312.810 ;
        RECT 622.670 312.430 622.900 312.810 ;
        RECT 625.430 312.800 625.610 313.890 ;
        RECT 627.000 312.800 627.180 313.890 ;
        RECT 778.390 313.390 780.000 326.920 ;
        RECT 852.580 314.130 852.830 337.550 ;
        RECT 855.150 314.200 855.400 337.710 ;
        RECT 869.670 333.110 870.520 333.810 ;
        RECT 865.520 330.490 866.770 331.110 ;
        RECT 869.890 330.750 870.160 333.110 ;
        RECT 870.740 331.110 871.790 332.200 ;
        RECT 872.470 330.750 872.710 330.760 ;
        RECT 869.790 330.560 872.800 330.750 ;
        RECT 864.660 330.160 867.480 330.190 ;
        RECT 864.660 330.140 867.520 330.160 ;
        RECT 864.570 330.000 867.520 330.140 ;
        RECT 869.840 330.140 870.160 330.560 ;
        RECT 871.190 330.170 871.420 330.400 ;
        RECT 872.470 330.180 872.710 330.560 ;
        RECT 869.840 330.000 870.130 330.140 ;
        RECT 864.570 329.850 864.920 330.000 ;
        RECT 864.570 329.710 864.940 329.850 ;
        RECT 864.570 329.610 864.960 329.710 ;
        RECT 864.680 329.590 864.960 329.610 ;
        RECT 864.690 328.370 864.960 329.590 ;
        RECT 864.610 327.910 864.960 328.370 ;
        RECT 859.430 327.610 859.660 327.820 ;
        RECT 852.590 314.020 852.820 314.130 ;
        RECT 855.170 314.020 855.400 314.200 ;
        RECT 859.410 314.210 859.660 327.610 ;
        RECT 862.010 327.570 862.240 327.820 ;
        RECT 861.980 327.440 862.240 327.570 ;
        RECT 861.980 327.090 862.230 327.440 ;
        RECT 864.690 327.340 864.960 327.910 ;
        RECT 866.000 329.630 866.230 329.850 ;
        RECT 867.280 329.750 867.520 330.000 ;
        RECT 861.890 326.530 862.430 327.090 ;
        RECT 861.980 326.350 862.230 326.530 ;
        RECT 864.280 326.370 865.220 327.340 ;
        RECT 861.980 325.970 862.240 326.350 ;
        RECT 861.980 324.880 862.230 325.970 ;
        RECT 861.980 324.500 862.240 324.880 ;
        RECT 861.980 323.410 862.230 324.500 ;
        RECT 864.690 323.750 864.960 326.370 ;
        RECT 866.000 323.910 866.270 329.630 ;
        RECT 867.280 329.590 867.570 329.750 ;
        RECT 867.290 329.470 867.570 329.590 ;
        RECT 867.300 328.380 867.570 329.470 ;
        RECT 867.290 328.000 867.570 328.380 ;
        RECT 867.300 326.910 867.570 328.000 ;
        RECT 867.290 326.530 867.570 326.910 ;
        RECT 867.300 325.440 867.570 326.530 ;
        RECT 867.290 325.060 867.570 325.440 ;
        RECT 867.300 323.970 867.570 325.060 ;
        RECT 869.880 324.270 870.130 330.000 ;
        RECT 871.180 324.280 871.430 330.170 ;
        RECT 872.470 330.050 872.740 330.180 ;
        RECT 872.480 330.020 872.740 330.050 ;
        RECT 872.490 329.780 872.740 330.020 ;
        RECT 872.490 329.470 872.970 329.780 ;
        RECT 872.490 328.930 872.740 329.470 ;
        RECT 872.480 328.550 872.740 328.930 ;
        RECT 872.490 327.460 872.740 328.550 ;
        RECT 872.480 327.080 872.740 327.460 ;
        RECT 872.490 325.990 872.740 327.080 ;
        RECT 872.480 325.610 872.740 325.990 ;
        RECT 872.490 324.520 872.740 325.610 ;
        RECT 872.480 324.290 872.740 324.520 ;
        RECT 869.900 324.140 870.130 324.270 ;
        RECT 871.190 324.140 871.420 324.280 ;
        RECT 872.480 324.140 872.710 324.290 ;
        RECT 865.990 323.780 866.270 323.910 ;
        RECT 867.290 323.790 867.570 323.970 ;
        RECT 864.710 323.590 864.940 323.750 ;
        RECT 861.980 323.030 862.240 323.410 ;
        RECT 865.990 323.270 866.260 323.780 ;
        RECT 867.290 323.590 867.520 323.790 ;
        RECT 871.190 323.760 871.400 324.140 ;
        RECT 885.340 323.770 888.860 324.520 ;
        RECT 876.070 323.760 888.860 323.770 ;
        RECT 871.190 323.430 888.860 323.760 ;
        RECT 871.900 323.270 872.180 323.430 ;
        RECT 876.070 323.300 888.860 323.430 ;
        RECT 861.980 321.940 862.230 323.030 ;
        RECT 865.990 323.000 872.220 323.270 ;
        RECT 871.900 322.960 872.180 323.000 ;
        RECT 885.340 322.740 888.860 323.300 ;
        RECT 861.980 321.560 862.240 321.940 ;
        RECT 872.810 321.790 873.270 322.040 ;
        RECT 874.010 321.790 875.020 321.930 ;
        RECT 872.810 321.560 875.020 321.790 ;
        RECT 861.980 320.470 862.230 321.560 ;
        RECT 872.810 321.470 873.270 321.560 ;
        RECT 874.010 321.430 875.020 321.560 ;
        RECT 874.490 321.130 874.640 321.430 ;
        RECT 875.760 321.130 876.000 321.140 ;
        RECT 873.080 320.940 876.090 321.130 ;
        RECT 869.940 320.620 870.170 320.840 ;
        RECT 861.980 320.090 862.240 320.470 ;
        RECT 861.980 319.000 862.230 320.090 ;
        RECT 861.980 318.620 862.240 319.000 ;
        RECT 861.980 317.530 862.230 318.620 ;
        RECT 861.980 317.150 862.240 317.530 ;
        RECT 861.980 316.060 862.230 317.150 ;
        RECT 861.980 315.680 862.240 316.060 ;
        RECT 861.980 314.590 862.230 315.680 ;
        RECT 869.940 315.100 870.210 320.620 ;
        RECT 873.130 320.550 873.440 320.940 ;
        RECT 875.760 320.560 876.000 320.940 ;
        RECT 873.130 320.380 873.420 320.550 ;
        RECT 875.760 320.430 876.030 320.560 ;
        RECT 875.770 320.400 876.030 320.430 ;
        RECT 861.980 314.290 862.240 314.590 ;
        RECT 859.410 314.070 859.620 314.210 ;
        RECT 862.010 314.070 862.240 314.290 ;
        RECT 859.410 314.060 862.240 314.070 ;
        RECT 869.830 314.340 870.340 315.100 ;
        RECT 873.170 314.870 873.420 320.380 ;
        RECT 875.780 319.310 876.030 320.400 ;
        RECT 875.770 318.930 876.030 319.310 ;
        RECT 875.780 317.840 876.030 318.930 ;
        RECT 875.770 317.460 876.030 317.840 ;
        RECT 875.780 316.370 876.030 317.460 ;
        RECT 875.770 315.990 876.030 316.370 ;
        RECT 875.780 314.900 876.030 315.990 ;
        RECT 873.030 314.340 873.480 314.870 ;
        RECT 875.770 314.670 876.030 314.900 ;
        RECT 875.770 314.520 876.000 314.670 ;
        RECT 859.410 313.950 862.230 314.060 ;
        RECT 869.830 313.960 873.480 314.340 ;
        RECT 873.030 313.950 873.480 313.960 ;
        RECT 859.410 313.910 862.220 313.950 ;
        RECT 603.190 312.130 605.060 312.290 ;
        RECT 607.740 312.280 609.580 312.300 ;
        RECT 612.260 312.280 614.100 312.300 ;
        RECT 616.730 312.280 616.910 312.420 ;
        RECT 618.320 312.280 618.500 312.420 ;
        RECT 621.110 312.290 621.290 312.430 ;
        RECT 622.700 312.290 622.880 312.430 ;
        RECT 625.410 312.420 625.640 312.800 ;
        RECT 626.990 312.420 627.220 312.800 ;
        RECT 621.070 312.280 622.910 312.290 ;
        RECT 625.430 312.280 625.610 312.420 ;
        RECT 627.020 312.280 627.200 312.420 ;
        RECT 607.740 312.210 615.420 312.280 ;
        RECT 607.740 312.140 615.430 312.210 ;
        RECT 603.190 310.770 603.470 312.130 ;
        RECT 607.810 311.120 607.980 312.140 ;
        RECT 613.780 312.120 615.430 312.140 ;
        RECT 616.690 312.140 622.910 312.280 ;
        RECT 616.690 312.120 618.530 312.140 ;
        RECT 621.070 312.130 622.910 312.140 ;
        RECT 613.360 311.460 613.830 311.840 ;
        RECT 615.220 311.670 615.430 312.120 ;
        RECT 616.200 311.670 616.630 311.740 ;
        RECT 615.220 311.490 616.630 311.670 ;
        RECT 608.400 311.120 609.070 311.430 ;
        RECT 607.800 310.840 609.070 311.120 ;
        RECT 596.970 310.540 597.660 310.600 ;
        RECT 594.260 310.040 595.060 310.500 ;
        RECT 594.400 308.520 594.680 310.040 ;
        RECT 596.950 309.690 597.680 310.540 ;
        RECT 596.970 309.630 597.660 309.690 ;
        RECT 385.690 308.060 385.920 308.440 ;
        RECT 594.160 308.250 594.890 308.520 ;
        RECT 603.180 308.500 603.490 310.770 ;
        RECT 607.810 310.470 607.980 310.840 ;
        RECT 608.400 310.580 609.070 310.840 ;
        RECT 613.450 310.940 613.690 311.460 ;
        RECT 616.200 311.420 616.630 311.490 ;
        RECT 617.010 310.940 617.190 312.120 ;
        RECT 620.610 311.720 621.020 311.990 ;
        RECT 620.560 311.560 621.020 311.720 ;
        RECT 620.560 311.420 620.980 311.560 ;
        RECT 613.450 310.780 617.200 310.940 ;
        RECT 607.070 309.830 607.980 310.470 ;
        RECT 615.490 310.050 615.710 310.110 ;
        RECT 620.560 310.050 620.830 311.420 ;
        RECT 603.780 308.500 604.740 308.670 ;
        RECT 603.120 308.220 604.740 308.500 ;
        RECT 603.180 307.600 603.490 308.220 ;
        RECT 603.780 308.110 604.740 308.220 ;
        RECT 600.790 307.440 604.170 307.600 ;
        RECT 600.800 307.270 600.970 307.440 ;
        RECT 602.370 307.270 602.540 307.440 ;
        RECT 603.970 307.270 604.140 307.440 ;
        RECT 211.890 306.130 212.870 306.360 ;
        RECT 215.360 306.130 216.340 306.360 ;
        RECT 218.830 306.130 219.810 306.360 ;
        RECT 222.300 306.130 223.280 306.360 ;
        RECT 225.770 306.130 226.750 306.360 ;
        RECT 231.930 306.120 232.910 306.350 ;
        RECT 235.400 306.120 236.380 306.350 ;
        RECT 238.870 306.120 239.850 306.350 ;
        RECT 242.340 306.120 243.320 306.350 ;
        RECT 245.810 306.120 246.790 306.350 ;
        RECT 251.990 306.120 252.970 306.350 ;
        RECT 255.460 306.120 256.440 306.350 ;
        RECT 258.930 306.120 259.910 306.350 ;
        RECT 262.400 306.120 263.380 306.350 ;
        RECT 265.870 306.120 266.850 306.350 ;
        RECT 272.040 306.120 273.020 306.350 ;
        RECT 275.510 306.120 276.490 306.350 ;
        RECT 278.980 306.120 279.960 306.350 ;
        RECT 282.450 306.120 283.430 306.350 ;
        RECT 285.920 306.120 286.900 306.350 ;
        RECT 288.530 304.740 290.200 306.490 ;
        RECT 591.500 305.990 592.700 307.160 ;
        RECT 600.770 306.890 601.000 307.270 ;
        RECT 601.560 306.890 601.790 307.270 ;
        RECT 602.350 306.890 602.580 307.270 ;
        RECT 603.140 306.890 603.370 307.270 ;
        RECT 603.930 306.890 604.160 307.270 ;
        RECT 299.530 304.740 301.590 304.860 ;
        RECT 288.530 303.820 301.590 304.740 ;
        RECT 379.110 304.590 379.340 305.570 ;
        RECT 385.690 304.590 385.920 305.570 ;
        RECT 591.900 304.235 592.150 305.990 ;
        RECT 600.800 305.800 600.980 306.890 ;
        RECT 601.580 305.800 601.760 306.890 ;
        RECT 602.370 305.800 602.550 306.890 ;
        RECT 603.150 305.800 603.330 306.890 ;
        RECT 603.940 305.800 604.120 306.890 ;
        RECT 600.770 305.420 601.000 305.800 ;
        RECT 601.560 305.420 601.790 305.800 ;
        RECT 602.350 305.420 602.580 305.800 ;
        RECT 603.140 305.420 603.370 305.800 ;
        RECT 603.930 305.420 604.160 305.800 ;
        RECT 601.580 305.280 601.760 305.420 ;
        RECT 603.170 305.280 603.350 305.420 ;
        RECT 607.810 305.370 607.980 309.830 ;
        RECT 608.380 309.570 609.020 309.990 ;
        RECT 615.490 309.820 620.830 310.050 ;
        RECT 621.060 309.860 621.570 309.910 ;
        RECT 621.730 309.900 621.940 312.130 ;
        RECT 625.390 312.120 627.230 312.280 ;
        RECT 622.930 310.860 623.780 311.300 ;
        RECT 626.390 310.920 626.610 312.120 ;
        RECT 778.390 311.440 780.640 313.390 ;
        RECT 639.220 311.040 639.650 311.100 ;
        RECT 629.480 310.920 629.710 310.940 ;
        RECT 622.110 309.900 622.800 309.990 ;
        RECT 621.730 309.860 622.800 309.900 ;
        RECT 608.550 306.020 608.810 309.570 ;
        RECT 609.350 308.400 610.000 308.620 ;
        RECT 609.350 308.370 610.500 308.400 ;
        RECT 609.350 308.220 613.630 308.370 ;
        RECT 609.350 308.050 610.500 308.220 ;
        RECT 611.800 308.050 612.020 308.220 ;
        RECT 613.400 308.050 613.620 308.220 ;
        RECT 610.220 307.890 610.460 308.050 ;
        RECT 610.220 307.670 610.450 307.890 ;
        RECT 611.010 307.670 611.240 308.050 ;
        RECT 611.800 307.670 612.030 308.050 ;
        RECT 612.590 307.670 612.820 308.050 ;
        RECT 613.380 307.880 613.620 308.050 ;
        RECT 613.380 307.670 613.610 307.880 ;
        RECT 610.230 306.580 610.410 307.670 ;
        RECT 611.030 306.580 611.210 307.670 ;
        RECT 611.830 306.580 612.010 307.670 ;
        RECT 612.610 306.580 612.790 307.670 ;
        RECT 613.390 306.580 613.570 307.670 ;
        RECT 615.490 307.560 615.710 309.820 ;
        RECT 621.060 309.720 622.800 309.860 ;
        RECT 621.060 309.620 621.570 309.720 ;
        RECT 621.730 309.610 622.800 309.720 ;
        RECT 621.040 308.340 621.520 308.410 ;
        RECT 617.810 308.190 621.520 308.340 ;
        RECT 617.830 308.020 618.050 308.190 ;
        RECT 619.390 308.020 619.610 308.190 ;
        RECT 620.990 308.130 621.520 308.190 ;
        RECT 620.990 308.020 621.210 308.130 ;
        RECT 617.810 307.860 618.050 308.020 ;
        RECT 617.810 307.640 618.040 307.860 ;
        RECT 618.600 307.640 618.830 308.020 ;
        RECT 619.390 307.640 619.620 308.020 ;
        RECT 620.180 307.640 620.410 308.020 ;
        RECT 620.970 307.850 621.210 308.020 ;
        RECT 620.970 307.640 621.200 307.850 ;
        RECT 615.360 307.140 615.840 307.560 ;
        RECT 614.050 306.690 617.470 306.830 ;
        RECT 610.220 306.200 610.450 306.580 ;
        RECT 611.010 306.200 611.240 306.580 ;
        RECT 611.800 306.200 612.030 306.580 ;
        RECT 612.590 306.200 612.820 306.580 ;
        RECT 613.380 306.200 613.610 306.580 ;
        RECT 614.080 306.530 614.270 306.690 ;
        RECT 615.640 306.530 615.830 306.690 ;
        RECT 617.250 306.530 617.440 306.690 ;
        RECT 617.820 306.550 618.000 307.640 ;
        RECT 618.620 306.550 618.800 307.640 ;
        RECT 619.420 306.550 619.600 307.640 ;
        RECT 620.200 306.550 620.380 307.640 ;
        RECT 620.980 306.550 621.160 307.640 ;
        RECT 608.370 305.710 609.040 306.020 ;
        RECT 609.640 305.370 609.790 305.380 ;
        RECT 601.540 305.120 603.380 305.280 ;
        RECT 606.450 305.230 609.880 305.370 ;
        RECT 603.220 304.470 603.370 305.120 ;
        RECT 606.490 305.060 606.640 305.230 ;
        RECT 608.080 305.060 608.230 305.230 ;
        RECT 609.640 305.060 609.790 305.230 ;
        RECT 610.230 305.110 610.410 306.200 ;
        RECT 611.030 305.110 611.210 306.200 ;
        RECT 611.830 305.110 612.010 306.200 ;
        RECT 612.610 305.110 612.790 306.200 ;
        RECT 613.390 305.110 613.570 306.200 ;
        RECT 614.050 306.150 614.280 306.530 ;
        RECT 615.630 306.150 615.860 306.530 ;
        RECT 617.210 306.150 617.440 306.530 ;
        RECT 617.810 306.170 618.040 306.550 ;
        RECT 618.600 306.170 618.830 306.550 ;
        RECT 619.390 306.170 619.620 306.550 ;
        RECT 620.180 306.170 620.410 306.550 ;
        RECT 620.970 306.170 621.200 306.550 ;
        RECT 606.470 304.680 606.700 305.060 ;
        RECT 607.260 304.680 607.490 305.060 ;
        RECT 608.050 304.680 608.280 305.060 ;
        RECT 608.840 304.680 609.070 305.060 ;
        RECT 609.630 304.680 609.860 305.060 ;
        RECT 610.220 304.730 610.450 305.110 ;
        RECT 611.010 304.940 611.240 305.110 ;
        RECT 611.000 304.730 611.240 304.940 ;
        RECT 611.800 304.730 612.030 305.110 ;
        RECT 612.590 304.730 612.820 305.110 ;
        RECT 613.380 304.730 613.610 305.110 ;
        RECT 614.070 305.060 614.230 306.150 ;
        RECT 615.650 305.060 615.810 306.150 ;
        RECT 617.230 305.060 617.390 306.150 ;
        RECT 617.820 305.080 618.000 306.170 ;
        RECT 618.620 305.080 618.800 306.170 ;
        RECT 619.420 305.080 619.600 306.170 ;
        RECT 620.200 305.080 620.380 306.170 ;
        RECT 620.980 305.080 621.160 306.170 ;
        RECT 621.730 305.370 621.940 309.610 ;
        RECT 622.110 309.530 622.800 309.610 ;
        RECT 623.160 306.150 623.390 310.860 ;
        RECT 626.390 310.770 629.720 310.920 ;
        RECT 629.480 308.460 629.710 310.770 ;
        RECT 639.200 310.590 639.670 311.040 ;
        RECT 645.280 310.810 645.650 310.870 ;
        RECT 639.220 310.530 639.650 310.590 ;
        RECT 645.260 310.460 645.670 310.810 ;
        RECT 645.280 310.400 645.650 310.460 ;
        RECT 631.570 308.560 632.520 309.450 ;
        RECT 633.810 309.340 634.640 310.080 ;
        RECT 641.670 310.000 642.170 310.380 ;
        RECT 666.200 309.280 667.570 309.340 ;
        RECT 629.110 308.110 629.710 308.460 ;
        RECT 629.480 307.730 629.710 308.110 ;
        RECT 639.110 307.940 639.810 308.300 ;
        RECT 627.570 307.570 630.950 307.730 ;
        RECT 627.580 307.400 627.750 307.570 ;
        RECT 629.150 307.400 629.320 307.570 ;
        RECT 629.480 307.560 629.710 307.570 ;
        RECT 630.750 307.400 630.920 307.570 ;
        RECT 627.550 307.020 627.780 307.400 ;
        RECT 628.340 307.020 628.570 307.400 ;
        RECT 629.130 307.020 629.360 307.400 ;
        RECT 629.920 307.020 630.150 307.400 ;
        RECT 630.710 307.020 630.940 307.400 ;
        RECT 622.960 305.600 623.650 306.150 ;
        RECT 627.580 305.930 627.760 307.020 ;
        RECT 628.360 305.930 628.540 307.020 ;
        RECT 629.150 305.930 629.330 307.020 ;
        RECT 629.930 305.930 630.110 307.020 ;
        RECT 630.720 305.930 630.900 307.020 ;
        RECT 627.550 305.550 627.780 305.930 ;
        RECT 628.340 305.550 628.570 305.930 ;
        RECT 629.130 305.550 629.360 305.930 ;
        RECT 629.920 305.550 630.150 305.930 ;
        RECT 630.710 305.550 630.940 305.930 ;
        RECT 639.370 305.640 639.550 307.940 ;
        RECT 643.210 307.820 643.780 308.500 ;
        RECT 666.180 307.830 667.590 309.280 ;
        RECT 639.690 306.040 640.140 306.730 ;
        RECT 643.440 305.690 643.580 307.820 ;
        RECT 666.200 307.770 667.570 307.830 ;
        RECT 643.750 306.580 644.170 306.780 ;
        RECT 645.180 306.580 646.160 306.890 ;
        RECT 643.750 306.370 646.160 306.580 ;
        RECT 643.750 306.100 644.170 306.370 ;
        RECT 645.180 306.110 646.160 306.370 ;
        RECT 628.360 305.410 628.540 305.550 ;
        RECT 629.950 305.410 630.130 305.550 ;
        RECT 639.370 305.530 639.630 305.640 ;
        RECT 624.730 305.370 624.880 305.380 ;
        RECT 621.540 305.230 624.970 305.370 ;
        RECT 628.320 305.250 630.160 305.410 ;
        RECT 639.400 305.260 639.630 305.530 ;
        RECT 643.440 305.520 643.680 305.690 ;
        RECT 643.450 305.310 643.680 305.520 ;
        RECT 607.300 304.530 607.450 304.680 ;
        RECT 608.880 304.530 609.030 304.680 ;
        RECT 610.260 304.530 610.440 304.730 ;
        RECT 288.530 301.980 290.200 303.820 ;
        RECT 211.850 298.300 212.830 298.530 ;
        RECT 215.320 298.300 216.300 298.530 ;
        RECT 218.790 298.300 219.770 298.530 ;
        RECT 222.260 298.300 223.240 298.530 ;
        RECT 225.730 298.300 226.710 298.530 ;
        RECT 231.820 298.300 232.800 298.530 ;
        RECT 235.290 298.300 236.270 298.530 ;
        RECT 238.760 298.300 239.740 298.530 ;
        RECT 242.230 298.300 243.210 298.530 ;
        RECT 245.700 298.300 246.680 298.530 ;
        RECT 251.930 298.300 252.910 298.530 ;
        RECT 255.400 298.300 256.380 298.530 ;
        RECT 258.870 298.300 259.850 298.530 ;
        RECT 262.340 298.300 263.320 298.530 ;
        RECT 265.810 298.300 266.790 298.530 ;
        RECT 272.040 298.300 273.020 298.530 ;
        RECT 275.510 298.300 276.490 298.530 ;
        RECT 278.980 298.300 279.960 298.530 ;
        RECT 282.450 298.300 283.430 298.530 ;
        RECT 285.920 298.300 286.900 298.530 ;
        RECT 4.630 296.310 5.610 296.540 ;
        RECT 8.100 296.310 9.080 296.540 ;
        RECT 11.570 296.310 12.550 296.540 ;
        RECT 17.970 296.290 18.950 296.520 ;
        RECT 21.440 296.290 22.420 296.520 ;
        RECT 24.910 296.290 25.890 296.520 ;
        RECT 31.340 296.320 32.320 296.550 ;
        RECT 34.810 296.320 35.790 296.550 ;
        RECT 38.280 296.320 39.260 296.550 ;
        RECT 44.570 296.320 45.550 296.550 ;
        RECT 48.040 296.320 49.020 296.550 ;
        RECT 51.510 296.320 52.490 296.550 ;
        RECT 57.840 296.290 58.820 296.520 ;
        RECT 61.310 296.290 62.290 296.520 ;
        RECT 64.780 296.290 65.760 296.520 ;
        RECT 71.110 296.320 72.090 296.550 ;
        RECT 74.580 296.320 75.560 296.550 ;
        RECT 78.050 296.320 79.030 296.550 ;
        RECT 84.240 296.340 85.220 296.570 ;
        RECT 87.710 296.340 88.690 296.570 ;
        RECT 91.180 296.340 92.160 296.570 ;
        RECT 97.660 296.560 98.640 296.790 ;
        RECT 101.130 296.560 102.110 296.790 ;
        RECT 211.850 291.720 212.830 291.950 ;
        RECT 215.320 291.720 216.300 291.950 ;
        RECT 218.790 291.720 219.770 291.950 ;
        RECT 222.260 291.720 223.240 291.950 ;
        RECT 225.730 291.720 226.710 291.950 ;
        RECT 231.820 291.720 232.800 291.950 ;
        RECT 235.290 291.720 236.270 291.950 ;
        RECT 238.760 291.720 239.740 291.950 ;
        RECT 242.230 291.720 243.210 291.950 ;
        RECT 245.700 291.720 246.680 291.950 ;
        RECT 251.930 291.720 252.910 291.950 ;
        RECT 255.400 291.720 256.380 291.950 ;
        RECT 258.870 291.720 259.850 291.950 ;
        RECT 262.340 291.720 263.320 291.950 ;
        RECT 265.810 291.720 266.790 291.950 ;
        RECT 272.040 291.720 273.020 291.950 ;
        RECT 275.510 291.720 276.490 291.950 ;
        RECT 278.980 291.720 279.960 291.950 ;
        RECT 282.450 291.720 283.430 291.950 ;
        RECT 285.920 291.720 286.900 291.950 ;
        RECT 4.630 289.730 5.610 289.960 ;
        RECT 8.100 289.730 9.080 289.960 ;
        RECT 11.570 289.730 12.550 289.960 ;
        RECT 17.970 289.710 18.950 289.940 ;
        RECT 21.440 289.710 22.420 289.940 ;
        RECT 24.910 289.710 25.890 289.940 ;
        RECT 31.340 289.740 32.320 289.970 ;
        RECT 34.810 289.740 35.790 289.970 ;
        RECT 38.280 289.740 39.260 289.970 ;
        RECT 44.570 289.740 45.550 289.970 ;
        RECT 48.040 289.740 49.020 289.970 ;
        RECT 51.510 289.740 52.490 289.970 ;
        RECT 57.840 289.710 58.820 289.940 ;
        RECT 61.310 289.710 62.290 289.940 ;
        RECT 64.780 289.710 65.760 289.940 ;
        RECT 71.110 289.740 72.090 289.970 ;
        RECT 74.580 289.740 75.560 289.970 ;
        RECT 78.050 289.740 79.030 289.970 ;
        RECT 84.240 289.760 85.220 289.990 ;
        RECT 87.710 289.760 88.690 289.990 ;
        RECT 91.180 289.760 92.160 289.990 ;
        RECT 97.660 289.980 98.640 290.210 ;
        RECT 101.130 289.980 102.110 290.210 ;
        RECT 294.310 285.390 295.950 286.500 ;
        RECT 296.130 285.390 297.600 286.310 ;
        RECT 211.850 285.140 212.830 285.370 ;
        RECT 215.320 285.140 216.300 285.370 ;
        RECT 218.790 285.140 219.770 285.370 ;
        RECT 222.260 285.140 223.240 285.370 ;
        RECT 225.730 285.140 226.710 285.370 ;
        RECT 231.820 285.140 232.800 285.370 ;
        RECT 235.290 285.140 236.270 285.370 ;
        RECT 238.760 285.140 239.740 285.370 ;
        RECT 242.230 285.140 243.210 285.370 ;
        RECT 245.700 285.140 246.680 285.370 ;
        RECT 251.930 285.140 252.910 285.370 ;
        RECT 255.400 285.140 256.380 285.370 ;
        RECT 258.870 285.140 259.850 285.370 ;
        RECT 262.340 285.140 263.320 285.370 ;
        RECT 265.810 285.140 266.790 285.370 ;
        RECT 272.040 285.140 273.020 285.370 ;
        RECT 275.510 285.140 276.490 285.370 ;
        RECT 278.980 285.140 279.960 285.370 ;
        RECT 282.450 285.140 283.430 285.370 ;
        RECT 285.920 285.140 286.900 285.370 ;
        RECT 294.310 284.690 297.600 285.390 ;
        RECT 294.310 284.140 295.950 284.690 ;
        RECT 296.130 284.250 297.600 284.690 ;
        RECT 4.630 283.150 5.610 283.380 ;
        RECT 8.100 283.150 9.080 283.380 ;
        RECT 11.570 283.150 12.550 283.380 ;
        RECT 17.970 283.130 18.950 283.360 ;
        RECT 21.440 283.130 22.420 283.360 ;
        RECT 24.910 283.130 25.890 283.360 ;
        RECT 31.340 283.160 32.320 283.390 ;
        RECT 34.810 283.160 35.790 283.390 ;
        RECT 38.280 283.160 39.260 283.390 ;
        RECT 44.570 283.160 45.550 283.390 ;
        RECT 48.040 283.160 49.020 283.390 ;
        RECT 51.510 283.160 52.490 283.390 ;
        RECT 57.840 283.130 58.820 283.360 ;
        RECT 61.310 283.130 62.290 283.360 ;
        RECT 64.780 283.130 65.760 283.360 ;
        RECT 71.110 283.160 72.090 283.390 ;
        RECT 74.580 283.160 75.560 283.390 ;
        RECT 78.050 283.160 79.030 283.390 ;
        RECT 84.240 283.180 85.220 283.410 ;
        RECT 87.710 283.180 88.690 283.410 ;
        RECT 91.180 283.180 92.160 283.410 ;
        RECT 97.660 283.400 98.640 283.630 ;
        RECT 101.130 283.400 102.110 283.630 ;
        RECT 154.850 278.010 156.390 278.690 ;
        RECT 149.840 277.980 156.390 278.010 ;
        RECT 118.140 277.750 119.120 277.980 ;
        RECT 121.610 277.750 122.590 277.980 ;
        RECT 125.080 277.750 126.060 277.980 ;
        RECT 128.550 277.750 129.530 277.980 ;
        RECT 132.020 277.750 133.000 277.980 ;
        RECT 135.490 277.750 136.470 277.980 ;
        RECT 138.960 277.750 139.940 277.980 ;
        RECT 142.430 277.750 143.410 277.980 ;
        RECT 145.900 277.750 146.880 277.980 ;
        RECT 149.370 277.750 156.390 277.980 ;
        RECT 149.840 277.690 156.390 277.750 ;
        RECT 154.850 277.150 156.390 277.690 ;
        RECT 4.630 276.570 5.610 276.800 ;
        RECT 8.100 276.570 9.080 276.800 ;
        RECT 11.570 276.570 12.550 276.800 ;
        RECT 17.970 276.550 18.950 276.780 ;
        RECT 21.440 276.550 22.420 276.780 ;
        RECT 24.910 276.550 25.890 276.780 ;
        RECT 31.340 276.580 32.320 276.810 ;
        RECT 34.810 276.580 35.790 276.810 ;
        RECT 38.280 276.580 39.260 276.810 ;
        RECT 44.570 276.580 45.550 276.810 ;
        RECT 48.040 276.580 49.020 276.810 ;
        RECT 51.510 276.580 52.490 276.810 ;
        RECT 57.840 276.550 58.820 276.780 ;
        RECT 61.310 276.550 62.290 276.780 ;
        RECT 64.780 276.550 65.760 276.780 ;
        RECT 71.110 276.580 72.090 276.810 ;
        RECT 74.580 276.580 75.560 276.810 ;
        RECT 78.050 276.580 79.030 276.810 ;
        RECT 84.240 276.600 85.220 276.830 ;
        RECT 87.710 276.600 88.690 276.830 ;
        RECT 91.180 276.600 92.160 276.830 ;
        RECT 97.660 276.820 98.640 277.050 ;
        RECT 101.130 276.820 102.110 277.050 ;
        RECT 118.140 271.170 119.120 271.400 ;
        RECT 121.610 271.170 122.590 271.400 ;
        RECT 125.080 271.170 126.060 271.400 ;
        RECT 128.550 271.170 129.530 271.400 ;
        RECT 132.020 271.170 133.000 271.400 ;
        RECT 135.490 271.170 136.470 271.400 ;
        RECT 138.960 271.170 139.940 271.400 ;
        RECT 142.430 271.170 143.410 271.400 ;
        RECT 145.900 271.170 146.880 271.400 ;
        RECT 149.370 271.170 150.350 271.400 ;
        RECT 4.630 269.990 5.610 270.220 ;
        RECT 8.100 269.990 9.080 270.220 ;
        RECT 11.570 269.990 12.550 270.220 ;
        RECT 17.970 269.970 18.950 270.200 ;
        RECT 21.440 269.970 22.420 270.200 ;
        RECT 24.910 269.970 25.890 270.200 ;
        RECT 31.340 270.000 32.320 270.230 ;
        RECT 34.810 270.000 35.790 270.230 ;
        RECT 38.280 270.000 39.260 270.230 ;
        RECT 44.570 270.000 45.550 270.230 ;
        RECT 48.040 270.000 49.020 270.230 ;
        RECT 51.510 270.000 52.490 270.230 ;
        RECT 57.840 269.970 58.820 270.200 ;
        RECT 61.310 269.970 62.290 270.200 ;
        RECT 64.780 269.970 65.760 270.200 ;
        RECT 71.110 270.000 72.090 270.230 ;
        RECT 74.580 270.000 75.560 270.230 ;
        RECT 78.050 270.000 79.030 270.230 ;
        RECT 84.240 270.020 85.220 270.250 ;
        RECT 87.710 270.020 88.690 270.250 ;
        RECT 91.180 270.020 92.160 270.250 ;
        RECT 97.660 270.240 98.640 270.470 ;
        RECT 101.130 270.240 102.110 270.470 ;
        RECT 299.530 252.160 301.590 303.820 ;
        RECT 602.070 303.750 602.850 304.190 ;
        RECT 603.140 304.030 603.590 304.470 ;
        RECT 607.250 304.380 610.440 304.530 ;
        RECT 611.000 304.570 611.170 304.730 ;
        RECT 612.600 304.570 612.770 304.730 ;
        RECT 614.050 304.680 614.280 305.060 ;
        RECT 615.630 304.680 615.860 305.060 ;
        RECT 617.210 304.680 617.440 305.060 ;
        RECT 617.810 304.700 618.040 305.080 ;
        RECT 618.600 304.910 618.830 305.080 ;
        RECT 618.590 304.700 618.830 304.910 ;
        RECT 619.390 304.700 619.620 305.080 ;
        RECT 620.180 304.700 620.410 305.080 ;
        RECT 620.970 304.900 621.200 305.080 ;
        RECT 621.580 305.060 621.730 305.230 ;
        RECT 623.170 305.060 623.320 305.230 ;
        RECT 624.730 305.060 624.880 305.230 ;
        RECT 620.970 304.700 621.210 304.900 ;
        RECT 614.050 304.570 614.250 304.680 ;
        RECT 611.000 304.460 614.250 304.570 ;
        RECT 609.020 304.350 610.440 304.380 ;
        RECT 610.940 304.430 614.250 304.460 ;
        RECT 610.940 304.420 612.840 304.430 ;
        RECT 610.940 304.120 611.350 304.420 ;
        RECT 614.050 304.060 614.250 304.430 ;
        RECT 617.220 304.530 617.440 304.680 ;
        RECT 618.590 304.540 618.760 304.700 ;
        RECT 620.190 304.540 620.360 304.700 ;
        RECT 618.590 304.530 620.430 304.540 ;
        RECT 617.220 304.450 620.430 304.530 ;
        RECT 621.010 304.490 621.210 304.700 ;
        RECT 621.560 304.680 621.790 305.060 ;
        RECT 622.350 304.680 622.580 305.060 ;
        RECT 623.140 304.680 623.370 305.060 ;
        RECT 623.930 304.680 624.160 305.060 ;
        RECT 624.720 304.680 624.950 305.060 ;
        RECT 622.390 304.530 622.540 304.680 ;
        RECT 623.970 304.530 624.120 304.680 ;
        RECT 622.340 304.490 624.160 304.530 ;
        RECT 617.220 304.390 620.470 304.450 ;
        RECT 617.220 304.360 618.980 304.390 ;
        RECT 620.070 304.090 620.470 304.390 ;
        RECT 621.010 304.380 624.160 304.490 ;
        RECT 621.010 304.330 622.500 304.380 ;
        RECT 629.060 303.900 629.270 305.250 ;
        RECT 628.890 303.550 629.510 303.900 ;
        RECT 379.110 301.120 379.340 302.100 ;
        RECT 385.690 301.120 385.920 302.100 ;
        RECT 591.900 301.750 592.150 303.185 ;
        RECT 696.370 302.210 697.530 302.270 ;
        RECT 591.540 300.580 592.740 301.750 ;
        RECT 696.350 300.840 697.550 302.210 ;
        RECT 696.370 300.780 697.530 300.840 ;
        RECT 379.110 297.650 379.340 298.630 ;
        RECT 385.690 297.650 385.920 298.630 ;
        RECT 747.780 297.850 748.100 297.910 ;
        RECT 712.440 297.790 712.830 297.850 ;
        RECT 694.980 297.410 695.320 297.470 ;
        RECT 632.300 296.050 633.790 297.100 ;
        RECT 682.075 297.075 682.365 297.120 ;
        RECT 684.475 297.075 684.765 297.120 ;
        RECT 689.755 297.075 690.045 297.120 ;
        RECT 682.075 296.935 690.045 297.075 ;
        RECT 694.960 297.030 695.340 297.410 ;
        RECT 699.565 297.035 699.855 297.080 ;
        RECT 701.965 297.035 702.255 297.080 ;
        RECT 707.245 297.035 707.535 297.080 ;
        RECT 694.980 296.970 695.320 297.030 ;
        RECT 682.075 296.890 682.365 296.935 ;
        RECT 684.475 296.890 684.765 296.935 ;
        RECT 689.755 296.890 690.045 296.935 ;
        RECT 699.565 296.895 707.535 297.035 ;
        RECT 712.420 297.020 712.850 297.790 ;
        RECT 730.050 297.750 730.400 297.810 ;
        RECT 717.175 297.095 717.465 297.140 ;
        RECT 719.575 297.095 719.865 297.140 ;
        RECT 724.855 297.095 725.145 297.140 ;
        RECT 712.440 296.960 712.830 297.020 ;
        RECT 717.175 296.955 725.145 297.095 ;
        RECT 730.030 297.000 730.420 297.750 ;
        RECT 747.760 297.110 748.120 297.850 ;
        RECT 765.480 297.710 765.860 297.770 ;
        RECT 765.460 297.110 765.880 297.710 ;
        RECT 734.875 297.045 735.165 297.090 ;
        RECT 737.275 297.045 737.565 297.090 ;
        RECT 742.555 297.045 742.845 297.090 ;
        RECT 747.780 297.050 748.100 297.110 ;
        RECT 717.175 296.910 717.465 296.955 ;
        RECT 719.575 296.910 719.865 296.955 ;
        RECT 724.855 296.910 725.145 296.955 ;
        RECT 730.050 296.940 730.400 297.000 ;
        RECT 699.565 296.850 699.855 296.895 ;
        RECT 701.965 296.850 702.255 296.895 ;
        RECT 707.245 296.850 707.535 296.895 ;
        RECT 734.875 296.905 742.845 297.045 ;
        RECT 734.875 296.860 735.165 296.905 ;
        RECT 737.275 296.860 737.565 296.905 ;
        RECT 742.555 296.860 742.845 296.905 ;
        RECT 752.615 297.035 752.905 297.080 ;
        RECT 755.015 297.035 755.305 297.080 ;
        RECT 760.295 297.035 760.585 297.080 ;
        RECT 765.480 297.050 765.860 297.110 ;
        RECT 752.615 296.895 760.585 297.035 ;
        RECT 752.615 296.850 752.905 296.895 ;
        RECT 755.015 296.850 755.305 296.895 ;
        RECT 760.295 296.850 760.585 296.895 ;
        RECT 778.390 296.820 780.000 311.440 ;
        RECT 834.110 306.970 834.460 307.030 ;
        RECT 811.510 306.940 834.460 306.970 ;
        RECT 811.400 306.710 834.460 306.940 ;
        RECT 811.400 306.660 811.770 306.710 ;
        RECT 834.110 306.570 834.460 306.710 ;
        RECT 794.420 305.550 795.990 306.260 ;
        RECT 813.070 306.220 813.550 306.380 ;
        RECT 814.780 306.220 815.190 306.230 ;
        RECT 798.495 306.135 798.785 306.180 ;
        RECT 800.895 306.135 801.185 306.180 ;
        RECT 806.175 306.135 806.465 306.180 ;
        RECT 798.495 305.995 806.465 306.135 ;
        RECT 798.495 305.950 798.785 305.995 ;
        RECT 800.895 305.950 801.185 305.995 ;
        RECT 806.175 305.950 806.465 305.995 ;
        RECT 813.070 306.080 815.190 306.220 ;
        RECT 813.070 305.990 813.550 306.080 ;
        RECT 814.780 305.970 815.190 306.080 ;
        RECT 816.255 306.135 816.545 306.180 ;
        RECT 818.655 306.135 818.945 306.180 ;
        RECT 823.935 306.135 824.225 306.180 ;
        RECT 816.255 305.995 824.225 306.135 ;
        RECT 816.255 305.950 816.545 305.995 ;
        RECT 818.655 305.950 818.945 305.995 ;
        RECT 823.935 305.950 824.225 305.995 ;
        RECT 829.140 306.140 829.460 306.160 ;
        RECT 837.520 306.140 837.840 306.220 ;
        RECT 829.140 305.940 837.840 306.140 ;
        RECT 811.400 305.800 811.780 305.890 ;
        RECT 811.400 305.700 817.880 305.800 ;
        RECT 829.140 305.760 829.460 305.940 ;
        RECT 837.520 305.820 837.840 305.940 ;
        RECT 811.400 305.640 818.000 305.700 ;
        RECT 797.050 305.550 797.360 305.620 ;
        RECT 811.400 305.600 811.780 305.640 ;
        RECT 794.420 305.320 797.360 305.550 ;
        RECT 817.620 305.410 818.000 305.640 ;
        RECT 834.120 305.650 834.590 305.730 ;
        RECT 838.870 305.650 839.160 305.910 ;
        RECT 834.120 305.540 839.160 305.650 ;
        RECT 839.430 305.730 839.710 305.810 ;
        RECT 842.860 305.730 843.140 305.980 ;
        RECT 839.430 305.580 843.140 305.730 ;
        RECT 839.430 305.570 843.020 305.580 ;
        RECT 834.120 305.470 839.060 305.540 ;
        RECT 834.120 305.430 834.590 305.470 ;
        RECT 839.430 305.410 839.710 305.570 ;
        RECT 832.800 305.380 833.110 305.390 ;
        RECT 794.420 305.030 795.990 305.320 ;
        RECT 797.050 305.230 797.360 305.320 ;
        RECT 799.850 304.890 800.240 305.300 ;
        RECT 799.910 304.880 800.190 304.890 ;
        RECT 832.690 304.820 833.200 305.380 ;
        RECT 832.800 304.790 833.110 304.820 ;
        RECT 832.380 296.910 833.290 296.990 ;
        RECT 832.380 296.820 833.380 296.910 ;
        RECT 680.560 296.470 681.010 296.660 ;
        RECT 698.090 296.470 698.540 296.610 ;
        RECT 715.660 296.470 716.110 296.660 ;
        RECT 733.380 296.470 733.830 296.630 ;
        RECT 751.110 296.590 751.560 296.610 ;
        RECT 770.550 296.590 833.380 296.820 ;
        RECT 751.110 296.470 833.380 296.590 ;
        RECT 680.560 296.430 833.380 296.470 ;
        RECT 678.560 296.370 833.380 296.430 ;
        RECT 678.560 296.290 751.560 296.370 ;
        RECT 678.560 296.270 680.920 296.290 ;
        RECT 698.090 296.270 698.540 296.290 ;
        RECT 751.110 296.270 751.560 296.290 ;
        RECT 770.550 296.260 833.380 296.370 ;
        RECT 683.420 295.790 683.850 296.060 ;
        RECT 700.900 295.810 701.350 296.130 ;
        RECT 778.390 296.050 780.000 296.260 ;
        RECT 832.380 296.130 833.380 296.260 ;
        RECT 683.460 295.780 683.820 295.790 ;
        RECT 379.110 294.180 379.340 295.160 ;
        RECT 385.690 294.930 385.920 295.160 ;
        RECT 379.110 289.180 379.340 290.160 ;
        RECT 385.620 289.590 386.000 294.930 ;
        RECT 603.190 294.720 603.420 295.100 ;
        RECT 604.770 294.720 605.000 295.100 ;
        RECT 607.710 294.730 607.940 295.110 ;
        RECT 609.290 294.730 609.520 295.110 ;
        RECT 612.230 294.730 612.460 295.110 ;
        RECT 613.810 294.730 614.040 295.110 ;
        RECT 603.210 293.630 603.390 294.720 ;
        RECT 604.780 293.630 604.960 294.720 ;
        RECT 607.730 293.640 607.910 294.730 ;
        RECT 609.300 293.640 609.480 294.730 ;
        RECT 612.250 293.640 612.430 294.730 ;
        RECT 613.820 293.640 614.000 294.730 ;
        RECT 616.660 294.710 616.890 295.090 ;
        RECT 618.240 294.710 618.470 295.090 ;
        RECT 621.040 294.720 621.270 295.100 ;
        RECT 622.620 294.720 622.850 295.100 ;
        RECT 603.190 293.470 603.420 293.630 ;
        RECT 603.140 293.110 603.420 293.470 ;
        RECT 604.770 293.250 605.000 293.630 ;
        RECT 607.710 293.260 607.940 293.640 ;
        RECT 609.290 293.260 609.520 293.640 ;
        RECT 612.230 293.260 612.460 293.640 ;
        RECT 613.810 293.260 614.040 293.640 ;
        RECT 616.680 293.620 616.860 294.710 ;
        RECT 618.250 293.620 618.430 294.710 ;
        RECT 621.060 293.630 621.240 294.720 ;
        RECT 622.630 293.630 622.810 294.720 ;
        RECT 625.360 294.710 625.590 295.090 ;
        RECT 626.940 294.710 627.170 295.090 ;
        RECT 604.800 293.110 604.980 293.250 ;
        RECT 607.730 293.120 607.930 293.260 ;
        RECT 609.320 293.120 609.500 293.260 ;
        RECT 612.250 293.120 612.430 293.260 ;
        RECT 613.840 293.120 614.020 293.260 ;
        RECT 616.660 293.240 616.890 293.620 ;
        RECT 618.240 293.240 618.470 293.620 ;
        RECT 621.040 293.250 621.270 293.630 ;
        RECT 622.620 293.250 622.850 293.630 ;
        RECT 625.380 293.620 625.560 294.710 ;
        RECT 626.950 293.620 627.130 294.710 ;
        RECT 673.630 294.250 674.140 294.280 ;
        RECT 700.770 294.250 701.630 294.460 ;
        RECT 673.600 293.800 701.630 294.250 ;
        RECT 603.140 292.950 605.010 293.110 ;
        RECT 607.690 293.100 609.530 293.120 ;
        RECT 612.210 293.100 614.050 293.120 ;
        RECT 616.680 293.100 616.860 293.240 ;
        RECT 618.270 293.100 618.450 293.240 ;
        RECT 621.060 293.110 621.240 293.250 ;
        RECT 622.650 293.110 622.830 293.250 ;
        RECT 625.360 293.240 625.590 293.620 ;
        RECT 626.940 293.240 627.170 293.620 ;
        RECT 621.020 293.100 622.860 293.110 ;
        RECT 625.380 293.100 625.560 293.240 ;
        RECT 626.970 293.100 627.150 293.240 ;
        RECT 607.690 293.030 615.370 293.100 ;
        RECT 607.690 292.960 615.380 293.030 ;
        RECT 603.140 291.590 603.420 292.950 ;
        RECT 607.760 291.940 607.930 292.960 ;
        RECT 613.730 292.940 615.380 292.960 ;
        RECT 616.640 292.960 622.860 293.100 ;
        RECT 616.640 292.940 618.480 292.960 ;
        RECT 621.020 292.950 622.860 292.960 ;
        RECT 613.310 292.280 613.780 292.660 ;
        RECT 615.170 292.490 615.380 292.940 ;
        RECT 616.150 292.490 616.580 292.560 ;
        RECT 615.170 292.310 616.580 292.490 ;
        RECT 608.350 291.940 609.020 292.250 ;
        RECT 607.750 291.660 609.020 291.940 ;
        RECT 596.920 291.360 597.610 291.420 ;
        RECT 594.210 290.860 595.010 291.320 ;
        RECT 385.690 289.180 385.920 289.590 ;
        RECT 594.350 289.340 594.630 290.860 ;
        RECT 596.900 290.510 597.630 291.360 ;
        RECT 596.920 290.450 597.610 290.510 ;
        RECT 594.110 289.070 594.840 289.340 ;
        RECT 603.130 289.320 603.440 291.590 ;
        RECT 607.760 291.290 607.930 291.660 ;
        RECT 608.350 291.400 609.020 291.660 ;
        RECT 613.400 291.760 613.640 292.280 ;
        RECT 616.150 292.240 616.580 292.310 ;
        RECT 616.960 291.760 617.140 292.940 ;
        RECT 620.560 292.540 620.970 292.810 ;
        RECT 620.510 292.380 620.970 292.540 ;
        RECT 620.510 292.240 620.930 292.380 ;
        RECT 613.400 291.600 617.150 291.760 ;
        RECT 607.020 290.650 607.930 291.290 ;
        RECT 615.440 290.870 615.660 290.930 ;
        RECT 620.510 290.870 620.780 292.240 ;
        RECT 603.730 289.320 604.690 289.490 ;
        RECT 603.070 289.040 604.690 289.320 ;
        RECT 603.130 288.420 603.440 289.040 ;
        RECT 603.730 288.930 604.690 289.040 ;
        RECT 591.250 287.170 592.740 288.410 ;
        RECT 600.740 288.260 604.120 288.420 ;
        RECT 600.750 288.090 600.920 288.260 ;
        RECT 602.320 288.090 602.490 288.260 ;
        RECT 603.920 288.090 604.090 288.260 ;
        RECT 600.720 287.710 600.950 288.090 ;
        RECT 601.510 287.710 601.740 288.090 ;
        RECT 602.300 287.710 602.530 288.090 ;
        RECT 603.090 287.710 603.320 288.090 ;
        RECT 603.880 287.710 604.110 288.090 ;
        RECT 379.110 285.710 379.340 286.690 ;
        RECT 385.690 285.710 385.920 286.690 ;
        RECT 591.870 285.465 592.120 287.170 ;
        RECT 600.750 286.620 600.930 287.710 ;
        RECT 601.530 286.620 601.710 287.710 ;
        RECT 602.320 286.620 602.500 287.710 ;
        RECT 603.100 286.620 603.280 287.710 ;
        RECT 603.890 286.620 604.070 287.710 ;
        RECT 600.720 286.240 600.950 286.620 ;
        RECT 601.510 286.240 601.740 286.620 ;
        RECT 602.300 286.240 602.530 286.620 ;
        RECT 603.090 286.240 603.320 286.620 ;
        RECT 603.880 286.240 604.110 286.620 ;
        RECT 601.530 286.100 601.710 286.240 ;
        RECT 603.120 286.100 603.300 286.240 ;
        RECT 607.760 286.190 607.930 290.650 ;
        RECT 608.330 290.390 608.970 290.810 ;
        RECT 615.440 290.640 620.780 290.870 ;
        RECT 621.010 290.680 621.520 290.730 ;
        RECT 621.680 290.720 621.890 292.950 ;
        RECT 625.340 292.940 627.180 293.100 ;
        RECT 622.880 291.680 623.730 292.120 ;
        RECT 626.340 291.740 626.560 292.940 ;
        RECT 673.630 292.600 674.140 293.800 ;
        RECT 700.770 293.770 701.630 293.800 ;
        RECT 833.080 293.130 833.380 296.130 ;
        RECT 855.890 295.720 856.380 295.840 ;
        RECT 854.310 295.690 856.380 295.720 ;
        RECT 854.000 295.490 856.380 295.690 ;
        RECT 858.730 295.680 859.130 295.790 ;
        RECT 858.730 295.540 860.070 295.680 ;
        RECT 854.000 295.220 854.600 295.490 ;
        RECT 855.890 295.460 856.380 295.490 ;
        RECT 856.850 295.100 857.300 295.490 ;
        RECT 858.730 295.470 859.130 295.540 ;
        RECT 842.360 294.470 842.660 294.590 ;
        RECT 843.760 294.470 844.280 294.530 ;
        RECT 842.360 294.240 844.280 294.470 ;
        RECT 842.360 294.090 842.660 294.240 ;
        RECT 843.760 294.130 844.280 294.240 ;
        RECT 639.170 291.860 639.600 291.920 ;
        RECT 629.430 291.740 629.660 291.760 ;
        RECT 622.060 290.720 622.750 290.810 ;
        RECT 621.680 290.680 622.750 290.720 ;
        RECT 608.500 286.840 608.760 290.390 ;
        RECT 609.300 289.220 609.950 289.440 ;
        RECT 609.300 289.190 610.450 289.220 ;
        RECT 609.300 289.040 613.580 289.190 ;
        RECT 609.300 288.870 610.450 289.040 ;
        RECT 611.750 288.870 611.970 289.040 ;
        RECT 613.350 288.870 613.570 289.040 ;
        RECT 610.170 288.710 610.410 288.870 ;
        RECT 610.170 288.490 610.400 288.710 ;
        RECT 610.960 288.490 611.190 288.870 ;
        RECT 611.750 288.490 611.980 288.870 ;
        RECT 612.540 288.490 612.770 288.870 ;
        RECT 613.330 288.700 613.570 288.870 ;
        RECT 613.330 288.490 613.560 288.700 ;
        RECT 610.180 287.400 610.360 288.490 ;
        RECT 610.980 287.400 611.160 288.490 ;
        RECT 611.780 287.400 611.960 288.490 ;
        RECT 612.560 287.400 612.740 288.490 ;
        RECT 613.340 287.400 613.520 288.490 ;
        RECT 615.440 288.380 615.660 290.640 ;
        RECT 621.010 290.540 622.750 290.680 ;
        RECT 621.010 290.440 621.520 290.540 ;
        RECT 621.680 290.430 622.750 290.540 ;
        RECT 620.990 289.160 621.470 289.230 ;
        RECT 617.760 289.010 621.470 289.160 ;
        RECT 617.780 288.840 618.000 289.010 ;
        RECT 619.340 288.840 619.560 289.010 ;
        RECT 620.940 288.950 621.470 289.010 ;
        RECT 620.940 288.840 621.160 288.950 ;
        RECT 617.760 288.680 618.000 288.840 ;
        RECT 617.760 288.460 617.990 288.680 ;
        RECT 618.550 288.460 618.780 288.840 ;
        RECT 619.340 288.460 619.570 288.840 ;
        RECT 620.130 288.460 620.360 288.840 ;
        RECT 620.920 288.670 621.160 288.840 ;
        RECT 620.920 288.460 621.150 288.670 ;
        RECT 615.310 287.960 615.790 288.380 ;
        RECT 614.000 287.510 617.420 287.650 ;
        RECT 610.170 287.020 610.400 287.400 ;
        RECT 610.960 287.020 611.190 287.400 ;
        RECT 611.750 287.020 611.980 287.400 ;
        RECT 612.540 287.020 612.770 287.400 ;
        RECT 613.330 287.020 613.560 287.400 ;
        RECT 614.030 287.350 614.220 287.510 ;
        RECT 615.590 287.350 615.780 287.510 ;
        RECT 617.200 287.350 617.390 287.510 ;
        RECT 617.770 287.370 617.950 288.460 ;
        RECT 618.570 287.370 618.750 288.460 ;
        RECT 619.370 287.370 619.550 288.460 ;
        RECT 620.150 287.370 620.330 288.460 ;
        RECT 620.930 287.370 621.110 288.460 ;
        RECT 608.320 286.530 608.990 286.840 ;
        RECT 609.590 286.190 609.740 286.200 ;
        RECT 601.490 285.940 603.330 286.100 ;
        RECT 606.400 286.050 609.830 286.190 ;
        RECT 603.170 285.290 603.320 285.940 ;
        RECT 606.440 285.880 606.590 286.050 ;
        RECT 608.030 285.880 608.180 286.050 ;
        RECT 609.590 285.880 609.740 286.050 ;
        RECT 610.180 285.930 610.360 287.020 ;
        RECT 610.980 285.930 611.160 287.020 ;
        RECT 611.780 285.930 611.960 287.020 ;
        RECT 612.560 285.930 612.740 287.020 ;
        RECT 613.340 285.930 613.520 287.020 ;
        RECT 614.000 286.970 614.230 287.350 ;
        RECT 615.580 286.970 615.810 287.350 ;
        RECT 617.160 286.970 617.390 287.350 ;
        RECT 617.760 286.990 617.990 287.370 ;
        RECT 618.550 286.990 618.780 287.370 ;
        RECT 619.340 286.990 619.570 287.370 ;
        RECT 620.130 286.990 620.360 287.370 ;
        RECT 620.920 286.990 621.150 287.370 ;
        RECT 606.420 285.500 606.650 285.880 ;
        RECT 607.210 285.500 607.440 285.880 ;
        RECT 608.000 285.500 608.230 285.880 ;
        RECT 608.790 285.500 609.020 285.880 ;
        RECT 609.580 285.500 609.810 285.880 ;
        RECT 610.170 285.550 610.400 285.930 ;
        RECT 610.960 285.760 611.190 285.930 ;
        RECT 610.950 285.550 611.190 285.760 ;
        RECT 611.750 285.550 611.980 285.930 ;
        RECT 612.540 285.550 612.770 285.930 ;
        RECT 613.330 285.550 613.560 285.930 ;
        RECT 614.020 285.880 614.180 286.970 ;
        RECT 615.600 285.880 615.760 286.970 ;
        RECT 617.180 285.880 617.340 286.970 ;
        RECT 617.770 285.900 617.950 286.990 ;
        RECT 618.570 285.900 618.750 286.990 ;
        RECT 619.370 285.900 619.550 286.990 ;
        RECT 620.150 285.900 620.330 286.990 ;
        RECT 620.930 285.900 621.110 286.990 ;
        RECT 621.680 286.190 621.890 290.430 ;
        RECT 622.060 290.350 622.750 290.430 ;
        RECT 623.110 286.970 623.340 291.680 ;
        RECT 626.340 291.590 629.670 291.740 ;
        RECT 629.430 289.280 629.660 291.590 ;
        RECT 639.150 291.410 639.620 291.860 ;
        RECT 645.230 291.630 645.600 291.690 ;
        RECT 639.170 291.350 639.600 291.410 ;
        RECT 645.210 291.280 645.620 291.630 ;
        RECT 645.230 291.220 645.600 291.280 ;
        RECT 631.320 289.670 632.060 290.280 ;
        RECT 633.760 290.160 634.590 290.900 ;
        RECT 641.620 290.820 642.120 291.200 ;
        RECT 629.060 288.930 629.660 289.280 ;
        RECT 629.430 288.550 629.660 288.930 ;
        RECT 639.060 288.760 639.760 289.120 ;
        RECT 627.520 288.390 630.900 288.550 ;
        RECT 627.530 288.220 627.700 288.390 ;
        RECT 629.100 288.220 629.270 288.390 ;
        RECT 629.430 288.380 629.660 288.390 ;
        RECT 630.700 288.220 630.870 288.390 ;
        RECT 627.500 287.840 627.730 288.220 ;
        RECT 628.290 287.840 628.520 288.220 ;
        RECT 629.080 287.840 629.310 288.220 ;
        RECT 629.870 287.840 630.100 288.220 ;
        RECT 630.660 287.840 630.890 288.220 ;
        RECT 622.910 286.420 623.600 286.970 ;
        RECT 627.530 286.750 627.710 287.840 ;
        RECT 628.310 286.750 628.490 287.840 ;
        RECT 629.100 286.750 629.280 287.840 ;
        RECT 629.880 286.750 630.060 287.840 ;
        RECT 630.670 286.750 630.850 287.840 ;
        RECT 627.500 286.370 627.730 286.750 ;
        RECT 628.290 286.370 628.520 286.750 ;
        RECT 629.080 286.370 629.310 286.750 ;
        RECT 629.870 286.370 630.100 286.750 ;
        RECT 630.660 286.370 630.890 286.750 ;
        RECT 639.320 286.460 639.500 288.760 ;
        RECT 643.160 288.640 643.730 289.320 ;
        RECT 639.640 286.860 640.090 287.550 ;
        RECT 643.390 286.510 643.530 288.640 ;
        RECT 643.700 287.400 644.120 287.600 ;
        RECT 645.130 287.400 646.110 287.710 ;
        RECT 643.700 287.190 646.110 287.400 ;
        RECT 643.700 286.920 644.120 287.190 ;
        RECT 645.130 286.930 646.110 287.190 ;
        RECT 628.310 286.230 628.490 286.370 ;
        RECT 629.900 286.230 630.080 286.370 ;
        RECT 639.320 286.350 639.580 286.460 ;
        RECT 624.680 286.190 624.830 286.200 ;
        RECT 621.490 286.050 624.920 286.190 ;
        RECT 628.270 286.070 630.110 286.230 ;
        RECT 639.350 286.080 639.580 286.350 ;
        RECT 643.390 286.340 643.630 286.510 ;
        RECT 643.400 286.130 643.630 286.340 ;
        RECT 607.250 285.350 607.400 285.500 ;
        RECT 608.830 285.350 608.980 285.500 ;
        RECT 610.210 285.350 610.390 285.550 ;
        RECT 601.930 284.540 602.880 285.010 ;
        RECT 603.090 284.850 603.540 285.290 ;
        RECT 607.200 285.200 610.390 285.350 ;
        RECT 610.950 285.390 611.120 285.550 ;
        RECT 612.550 285.390 612.720 285.550 ;
        RECT 614.000 285.500 614.230 285.880 ;
        RECT 615.580 285.500 615.810 285.880 ;
        RECT 617.160 285.500 617.390 285.880 ;
        RECT 617.760 285.520 617.990 285.900 ;
        RECT 618.550 285.730 618.780 285.900 ;
        RECT 618.540 285.520 618.780 285.730 ;
        RECT 619.340 285.520 619.570 285.900 ;
        RECT 620.130 285.520 620.360 285.900 ;
        RECT 620.920 285.720 621.150 285.900 ;
        RECT 621.530 285.880 621.680 286.050 ;
        RECT 623.120 285.880 623.270 286.050 ;
        RECT 624.680 285.880 624.830 286.050 ;
        RECT 620.920 285.520 621.160 285.720 ;
        RECT 614.000 285.390 614.200 285.500 ;
        RECT 610.950 285.280 614.200 285.390 ;
        RECT 608.970 285.170 610.390 285.200 ;
        RECT 610.890 285.250 614.200 285.280 ;
        RECT 610.890 285.240 612.790 285.250 ;
        RECT 610.890 284.940 611.300 285.240 ;
        RECT 614.000 284.880 614.200 285.250 ;
        RECT 617.170 285.350 617.390 285.500 ;
        RECT 618.540 285.360 618.710 285.520 ;
        RECT 620.140 285.360 620.310 285.520 ;
        RECT 618.540 285.350 620.380 285.360 ;
        RECT 617.170 285.270 620.380 285.350 ;
        RECT 620.960 285.310 621.160 285.520 ;
        RECT 621.510 285.500 621.740 285.880 ;
        RECT 622.300 285.500 622.530 285.880 ;
        RECT 623.090 285.500 623.320 285.880 ;
        RECT 623.880 285.500 624.110 285.880 ;
        RECT 624.670 285.500 624.900 285.880 ;
        RECT 622.340 285.350 622.490 285.500 ;
        RECT 623.920 285.350 624.070 285.500 ;
        RECT 622.290 285.310 624.110 285.350 ;
        RECT 617.170 285.210 620.420 285.270 ;
        RECT 617.170 285.180 618.930 285.210 ;
        RECT 620.020 284.910 620.420 285.210 ;
        RECT 620.960 285.200 624.110 285.310 ;
        RECT 620.960 285.150 622.450 285.200 ;
        RECT 629.010 284.720 629.220 286.070 ;
        RECT 379.110 282.240 379.340 283.220 ;
        RECT 385.690 282.240 385.920 283.220 ;
        RECT 591.870 282.870 592.120 284.415 ;
        RECT 628.840 284.370 629.460 284.720 ;
        RECT 591.190 281.630 592.680 282.870 ;
        RECT 379.110 278.770 379.340 279.750 ;
        RECT 385.690 278.770 385.920 279.750 ;
        RECT 632.340 277.530 633.560 278.800 ;
        RECT 379.110 275.300 379.340 276.280 ;
        RECT 385.690 276.030 385.920 276.280 ;
        RECT 603.110 276.250 603.340 276.630 ;
        RECT 604.690 276.250 604.920 276.630 ;
        RECT 607.630 276.260 607.860 276.640 ;
        RECT 609.210 276.260 609.440 276.640 ;
        RECT 612.150 276.260 612.380 276.640 ;
        RECT 613.730 276.260 613.960 276.640 ;
        RECT 379.130 270.320 379.360 271.300 ;
        RECT 385.620 270.690 386.000 276.030 ;
        RECT 603.130 275.160 603.310 276.250 ;
        RECT 604.700 275.160 604.880 276.250 ;
        RECT 607.650 275.170 607.830 276.260 ;
        RECT 609.220 275.170 609.400 276.260 ;
        RECT 612.170 275.170 612.350 276.260 ;
        RECT 613.740 275.170 613.920 276.260 ;
        RECT 616.580 276.240 616.810 276.620 ;
        RECT 618.160 276.240 618.390 276.620 ;
        RECT 620.960 276.250 621.190 276.630 ;
        RECT 622.540 276.250 622.770 276.630 ;
        RECT 603.110 275.000 603.340 275.160 ;
        RECT 603.060 274.640 603.340 275.000 ;
        RECT 604.690 274.780 604.920 275.160 ;
        RECT 607.630 274.790 607.860 275.170 ;
        RECT 609.210 274.790 609.440 275.170 ;
        RECT 612.150 274.790 612.380 275.170 ;
        RECT 613.730 274.790 613.960 275.170 ;
        RECT 616.600 275.150 616.780 276.240 ;
        RECT 618.170 275.150 618.350 276.240 ;
        RECT 620.980 275.160 621.160 276.250 ;
        RECT 622.550 275.160 622.730 276.250 ;
        RECT 625.280 276.240 625.510 276.620 ;
        RECT 626.860 276.240 627.090 276.620 ;
        RECT 604.720 274.640 604.900 274.780 ;
        RECT 607.650 274.650 607.850 274.790 ;
        RECT 609.240 274.650 609.420 274.790 ;
        RECT 612.170 274.650 612.350 274.790 ;
        RECT 613.760 274.650 613.940 274.790 ;
        RECT 616.580 274.770 616.810 275.150 ;
        RECT 618.160 274.770 618.390 275.150 ;
        RECT 620.960 274.780 621.190 275.160 ;
        RECT 622.540 274.780 622.770 275.160 ;
        RECT 625.300 275.150 625.480 276.240 ;
        RECT 626.870 275.150 627.050 276.240 ;
        RECT 603.060 274.480 604.930 274.640 ;
        RECT 607.610 274.630 609.450 274.650 ;
        RECT 612.130 274.630 613.970 274.650 ;
        RECT 616.600 274.630 616.780 274.770 ;
        RECT 618.190 274.630 618.370 274.770 ;
        RECT 620.980 274.640 621.160 274.780 ;
        RECT 622.570 274.640 622.750 274.780 ;
        RECT 625.280 274.770 625.510 275.150 ;
        RECT 626.860 274.770 627.090 275.150 ;
        RECT 620.940 274.630 622.780 274.640 ;
        RECT 625.300 274.630 625.480 274.770 ;
        RECT 626.890 274.630 627.070 274.770 ;
        RECT 673.630 274.680 674.110 292.600 ;
        RECT 832.730 291.570 834.140 293.130 ;
        RECT 836.000 293.120 836.450 293.980 ;
        RECT 840.450 293.530 840.850 293.750 ;
        RECT 852.620 293.530 853.710 293.780 ;
        RECT 840.450 293.360 853.710 293.530 ;
        RECT 840.450 293.190 840.850 293.360 ;
        RECT 836.060 292.980 836.310 293.120 ;
        RECT 852.620 292.980 853.710 293.360 ;
        RECT 819.020 290.980 819.520 291.070 ;
        RECT 813.410 290.710 819.520 290.980 ;
        RECT 820.000 290.860 820.400 290.920 ;
        RECT 813.410 290.650 819.150 290.710 ;
        RECT 694.740 290.530 696.190 290.590 ;
        RECT 694.720 289.280 696.210 290.530 ;
        RECT 813.410 290.110 813.700 290.650 ;
        RECT 819.980 290.470 820.420 290.860 ;
        RECT 821.860 290.640 822.240 290.780 ;
        RECT 820.000 290.410 820.400 290.470 ;
        RECT 821.860 290.450 824.050 290.640 ;
        RECT 821.860 290.290 822.240 290.450 ;
        RECT 678.120 288.720 696.210 289.280 ;
        RECT 678.150 287.370 678.480 288.720 ;
        RECT 694.720 288.550 696.210 288.720 ;
        RECT 813.440 288.830 813.690 290.110 ;
        RECT 823.800 289.010 824.050 290.450 ;
        RECT 827.420 289.300 827.900 289.340 ;
        RECT 831.950 289.300 832.430 289.320 ;
        RECT 824.530 289.010 824.910 289.150 ;
        RECT 823.800 288.840 824.910 289.010 ;
        RECT 827.420 289.080 832.430 289.300 ;
        RECT 827.420 288.940 827.900 289.080 ;
        RECT 831.950 288.920 832.430 289.080 ;
        RECT 694.740 288.490 696.190 288.550 ;
        RECT 678.150 280.240 678.470 287.370 ;
        RECT 802.010 281.550 803.000 281.610 ;
        RECT 799.630 281.000 800.050 281.360 ;
        RECT 801.990 280.560 803.020 281.550 ;
        RECT 802.010 280.500 803.000 280.560 ;
        RECT 679.950 280.240 680.370 280.310 ;
        RECT 678.150 280.010 680.370 280.240 ;
        RECT 678.150 280.000 680.200 280.010 ;
        RECT 678.150 279.890 678.470 280.000 ;
        RECT 694.880 279.860 695.840 279.970 ;
        RECT 700.050 279.860 700.460 279.970 ;
        RECT 694.680 279.670 700.460 279.860 ;
        RECT 713.330 279.820 714.110 279.960 ;
        RECT 717.840 279.820 718.200 279.950 ;
        RECT 683.140 279.110 683.730 279.610 ;
        RECT 694.680 279.540 700.170 279.670 ;
        RECT 694.880 279.220 695.840 279.540 ;
        RECT 700.640 279.530 701.150 279.720 ;
        RECT 712.990 279.680 718.200 279.820 ;
        RECT 727.130 279.820 727.920 279.860 ;
        RECT 735.080 279.840 735.440 279.980 ;
        RECT 729.950 279.820 735.440 279.840 ;
        RECT 727.130 279.710 735.440 279.820 ;
        RECT 747.410 279.800 748.180 279.920 ;
        RECT 752.560 279.800 752.920 279.940 ;
        RECT 712.990 279.610 717.980 279.680 ;
        RECT 700.530 279.070 701.150 279.530 ;
        RECT 713.330 279.220 714.110 279.610 ;
        RECT 727.130 279.570 735.240 279.710 ;
        RECT 747.410 279.670 752.920 279.800 ;
        RECT 727.130 279.530 730.110 279.570 ;
        RECT 747.410 279.550 752.800 279.670 ;
        RECT 700.640 279.020 701.150 279.070 ;
        RECT 718.220 279.050 718.760 279.500 ;
        RECT 727.130 279.200 727.920 279.530 ;
        RECT 735.540 279.490 735.930 279.550 ;
        RECT 735.520 279.150 735.950 279.490 ;
        RECT 747.410 279.180 748.180 279.550 ;
        RECT 735.540 279.090 735.930 279.150 ;
        RECT 752.950 279.100 753.450 279.480 ;
        RECT 813.440 277.860 813.700 288.830 ;
        RECT 824.530 288.660 824.910 288.840 ;
        RECT 833.220 288.650 833.800 289.020 ;
        RECT 833.990 288.670 834.320 288.860 ;
        RECT 836.070 288.670 836.300 292.980 ;
        RECT 843.740 292.380 844.360 292.820 ;
        RECT 846.580 292.380 847.000 292.400 ;
        RECT 843.740 292.240 847.000 292.380 ;
        RECT 846.580 292.100 847.000 292.240 ;
        RECT 848.980 291.750 849.930 292.560 ;
        RECT 859.900 292.190 860.050 295.540 ;
        RECT 859.900 292.170 863.020 292.190 ;
        RECT 859.900 292.010 863.080 292.170 ;
        RECT 862.710 291.730 863.080 292.010 ;
        RECT 865.070 292.150 866.400 292.490 ;
        RECT 868.130 292.150 869.240 292.260 ;
        RECT 865.070 291.830 869.240 292.150 ;
        RECT 865.070 291.710 866.400 291.830 ;
        RECT 868.130 291.690 869.240 291.830 ;
        RECT 856.930 290.030 857.300 290.090 ;
        RECT 856.910 289.620 857.320 290.030 ;
        RECT 856.930 289.560 857.300 289.620 ;
        RECT 833.990 288.520 836.300 288.670 ;
        RECT 840.490 288.520 840.840 288.580 ;
        RECT 833.990 288.460 834.320 288.520 ;
        RECT 836.070 288.500 836.300 288.520 ;
        RECT 825.480 288.210 825.810 288.360 ;
        RECT 823.650 288.040 825.810 288.210 ;
        RECT 840.470 288.150 840.860 288.520 ;
        RECT 840.490 288.090 840.840 288.150 ;
        RECT 821.850 287.410 822.180 287.440 ;
        RECT 823.650 287.410 823.820 288.040 ;
        RECT 825.480 287.910 825.810 288.040 ;
        RECT 821.850 287.220 823.820 287.410 ;
        RECT 821.850 286.990 822.180 287.220 ;
        RECT 823.650 287.210 823.820 287.220 ;
        RECT 814.400 286.730 815.110 286.870 ;
        RECT 840.320 286.730 840.920 286.880 ;
        RECT 814.400 286.450 840.920 286.730 ;
        RECT 814.400 286.430 824.410 286.450 ;
        RECT 814.400 286.220 815.110 286.430 ;
        RECT 840.320 286.410 840.920 286.450 ;
        RECT 818.990 285.880 819.460 285.940 ;
        RECT 818.970 285.400 819.480 285.880 ;
        RECT 816.250 285.170 817.370 285.390 ;
        RECT 818.990 285.340 819.460 285.400 ;
        RECT 819.960 285.170 820.380 285.580 ;
        RECT 832.890 285.300 834.320 286.290 ;
        RECT 816.250 285.090 820.380 285.170 ;
        RECT 816.250 284.930 820.180 285.090 ;
        RECT 816.250 284.550 817.370 284.930 ;
        RECT 856.030 284.800 856.360 285.040 ;
        RECT 855.340 284.790 856.360 284.800 ;
        RECT 825.550 284.590 856.360 284.790 ;
        RECT 858.890 284.610 859.160 284.700 ;
        RECT 825.550 284.580 856.210 284.590 ;
        RECT 825.550 284.570 855.490 284.580 ;
        RECT 825.550 284.310 850.560 284.570 ;
        RECT 853.860 284.420 855.050 284.430 ;
        RECT 856.950 284.420 857.410 284.510 ;
        RECT 821.670 281.040 822.170 281.390 ;
        RECT 825.550 281.140 825.820 284.310 ;
        RECT 853.860 284.210 857.410 284.420 ;
        RECT 858.890 284.450 860.390 284.610 ;
        RECT 858.890 284.300 859.160 284.450 ;
        RECT 853.860 284.160 855.050 284.210 ;
        RECT 852.880 283.700 853.430 283.850 ;
        RECT 853.860 283.700 854.120 284.160 ;
        RECT 856.950 284.140 857.410 284.210 ;
        RECT 852.880 283.350 854.120 283.700 ;
        RECT 852.880 283.220 853.430 283.350 ;
        RECT 830.930 281.150 831.240 281.240 ;
        RECT 841.020 281.180 841.500 281.550 ;
        RECT 835.340 281.150 835.650 281.180 ;
        RECT 820.780 280.550 821.220 280.880 ;
        RECT 823.320 280.790 823.700 280.930 ;
        RECT 825.290 280.790 826.060 281.140 ;
        RECT 830.930 281.000 835.650 281.150 ;
        RECT 830.930 280.860 831.240 281.000 ;
        RECT 835.340 280.800 835.650 281.000 ;
        RECT 843.830 281.090 844.290 281.210 ;
        RECT 848.300 281.090 848.760 281.160 ;
        RECT 843.830 280.950 848.760 281.090 ;
        RECT 849.710 281.010 850.050 281.070 ;
        RECT 823.320 280.590 826.060 280.790 ;
        RECT 828.050 280.730 828.480 280.790 ;
        RECT 823.320 280.470 823.700 280.590 ;
        RECT 825.290 280.300 826.060 280.590 ;
        RECT 828.030 280.270 828.500 280.730 ;
        RECT 829.020 280.620 829.420 280.680 ;
        RECT 828.050 280.210 828.480 280.270 ;
        RECT 829.000 280.000 829.440 280.620 ;
        RECT 836.600 280.550 837.050 280.930 ;
        RECT 843.830 280.860 844.290 280.950 ;
        RECT 848.300 280.810 848.760 280.950 ;
        RECT 837.200 280.580 837.620 280.670 ;
        RECT 838.590 280.580 839.100 280.650 ;
        RECT 837.200 280.420 839.100 280.580 ;
        RECT 837.200 280.320 837.620 280.420 ;
        RECT 838.200 280.410 838.410 280.420 ;
        RECT 838.590 280.310 839.100 280.420 ;
        RECT 841.010 280.270 841.460 280.600 ;
        RECT 849.690 280.590 850.070 281.010 ;
        RECT 850.260 280.700 850.680 280.760 ;
        RECT 851.890 280.700 852.700 280.870 ;
        RECT 849.710 280.530 850.050 280.590 ;
        RECT 850.260 280.500 852.700 280.700 ;
        RECT 850.260 280.400 850.680 280.500 ;
        RECT 841.940 280.300 842.340 280.360 ;
        RECT 829.020 279.940 829.420 280.000 ;
        RECT 839.490 279.920 839.930 280.130 ;
        RECT 841.920 279.880 842.360 280.300 ;
        RECT 851.890 280.190 852.700 280.500 ;
        RECT 841.940 279.820 842.340 279.880 ;
        RECT 836.490 278.520 837.190 278.700 ;
        RECT 834.650 278.280 837.190 278.520 ;
        RECT 834.670 277.860 835.000 278.280 ;
        RECT 836.490 278.180 837.190 278.280 ;
        RECT 840.630 278.220 841.330 278.700 ;
        RECT 813.440 277.830 835.000 277.860 ;
        RECT 813.440 277.610 838.210 277.830 ;
        RECT 813.440 277.580 813.700 277.610 ;
        RECT 834.710 277.590 838.210 277.610 ;
        RECT 834.740 276.470 835.000 277.590 ;
        RECT 853.010 277.560 853.570 278.110 ;
        RECT 834.540 276.100 835.270 276.470 ;
        RECT 673.630 274.650 677.360 274.680 ;
        RECT 678.790 274.650 679.210 274.660 ;
        RECT 679.790 274.650 680.350 274.890 ;
        RECT 681.840 274.650 682.100 274.780 ;
        RECT 607.610 274.560 615.290 274.630 ;
        RECT 607.610 274.490 615.300 274.560 ;
        RECT 603.060 273.120 603.340 274.480 ;
        RECT 607.680 273.470 607.850 274.490 ;
        RECT 613.650 274.470 615.300 274.490 ;
        RECT 616.560 274.490 622.780 274.630 ;
        RECT 616.560 274.470 618.400 274.490 ;
        RECT 620.940 274.480 622.780 274.490 ;
        RECT 613.230 273.810 613.700 274.190 ;
        RECT 615.090 274.020 615.300 274.470 ;
        RECT 616.070 274.020 616.500 274.090 ;
        RECT 615.090 273.840 616.500 274.020 ;
        RECT 608.270 273.470 608.940 273.780 ;
        RECT 607.670 273.190 608.940 273.470 ;
        RECT 596.840 272.890 597.530 272.950 ;
        RECT 594.130 272.390 594.930 272.850 ;
        RECT 594.270 270.870 594.550 272.390 ;
        RECT 596.820 272.040 597.550 272.890 ;
        RECT 596.840 271.980 597.530 272.040 ;
        RECT 385.710 270.320 385.940 270.690 ;
        RECT 594.030 270.600 594.760 270.870 ;
        RECT 603.050 270.850 603.360 273.120 ;
        RECT 607.680 272.820 607.850 273.190 ;
        RECT 608.270 272.930 608.940 273.190 ;
        RECT 613.320 273.290 613.560 273.810 ;
        RECT 616.070 273.770 616.500 273.840 ;
        RECT 616.880 273.290 617.060 274.470 ;
        RECT 620.480 274.070 620.890 274.340 ;
        RECT 620.430 273.910 620.890 274.070 ;
        RECT 620.430 273.770 620.850 273.910 ;
        RECT 613.320 273.130 617.070 273.290 ;
        RECT 606.940 272.180 607.850 272.820 ;
        RECT 615.360 272.400 615.580 272.460 ;
        RECT 620.430 272.400 620.700 273.770 ;
        RECT 603.650 270.850 604.610 271.020 ;
        RECT 602.990 270.570 604.610 270.850 ;
        RECT 591.250 268.980 592.620 270.020 ;
        RECT 603.050 269.950 603.360 270.570 ;
        RECT 603.650 270.460 604.610 270.570 ;
        RECT 600.660 269.790 604.040 269.950 ;
        RECT 600.670 269.620 600.840 269.790 ;
        RECT 602.240 269.620 602.410 269.790 ;
        RECT 603.840 269.620 604.010 269.790 ;
        RECT 600.640 269.240 600.870 269.620 ;
        RECT 601.430 269.240 601.660 269.620 ;
        RECT 602.220 269.240 602.450 269.620 ;
        RECT 603.010 269.240 603.240 269.620 ;
        RECT 603.800 269.240 604.030 269.620 ;
        RECT 379.130 266.850 379.360 267.830 ;
        RECT 385.710 266.850 385.940 267.830 ;
        RECT 591.710 267.205 591.960 268.980 ;
        RECT 600.670 268.150 600.850 269.240 ;
        RECT 601.450 268.150 601.630 269.240 ;
        RECT 602.240 268.150 602.420 269.240 ;
        RECT 603.020 268.150 603.200 269.240 ;
        RECT 603.810 268.150 603.990 269.240 ;
        RECT 600.640 267.770 600.870 268.150 ;
        RECT 601.430 267.770 601.660 268.150 ;
        RECT 602.220 267.770 602.450 268.150 ;
        RECT 603.010 267.770 603.240 268.150 ;
        RECT 603.800 267.770 604.030 268.150 ;
        RECT 601.450 267.630 601.630 267.770 ;
        RECT 603.040 267.630 603.220 267.770 ;
        RECT 607.680 267.720 607.850 272.180 ;
        RECT 608.250 271.920 608.890 272.340 ;
        RECT 615.360 272.170 620.700 272.400 ;
        RECT 620.930 272.210 621.440 272.260 ;
        RECT 621.600 272.250 621.810 274.480 ;
        RECT 625.260 274.470 627.100 274.630 ;
        RECT 673.630 274.480 682.100 274.650 ;
        RECT 683.780 274.590 684.160 274.640 ;
        RECT 685.430 274.590 685.940 274.820 ;
        RECT 689.090 274.590 689.470 274.650 ;
        RECT 622.800 273.210 623.650 273.650 ;
        RECT 626.260 273.270 626.480 274.470 ;
        RECT 673.630 274.440 679.210 274.480 ;
        RECT 673.630 274.380 679.170 274.440 ;
        RECT 679.790 274.390 680.350 274.480 ;
        RECT 681.840 274.410 682.100 274.480 ;
        RECT 673.630 274.330 677.360 274.380 ;
        RECT 680.980 274.210 681.580 274.230 ;
        RECT 683.150 274.210 683.580 274.480 ;
        RECT 683.780 274.450 689.470 274.590 ;
        RECT 701.010 274.610 701.390 274.660 ;
        RECT 702.660 274.610 703.170 274.840 ;
        RECT 718.580 274.710 718.960 274.760 ;
        RECT 720.230 274.710 720.740 274.940 ;
        RECT 723.890 274.710 724.270 274.770 ;
        RECT 706.320 274.610 706.700 274.670 ;
        RECT 683.780 274.330 684.160 274.450 ;
        RECT 679.140 274.070 683.580 274.210 ;
        RECT 685.430 274.130 685.940 274.450 ;
        RECT 689.090 274.340 689.470 274.450 ;
        RECT 686.520 274.160 687.110 274.260 ;
        RECT 690.500 274.160 690.740 274.380 ;
        RECT 680.980 273.840 681.580 274.070 ;
        RECT 683.150 273.980 683.580 274.070 ;
        RECT 686.380 274.030 690.740 274.160 ;
        RECT 691.000 274.260 691.380 274.320 ;
        RECT 692.770 274.270 693.550 274.510 ;
        RECT 692.770 274.260 693.830 274.270 ;
        RECT 691.000 274.110 693.830 274.260 ;
        RECT 698.210 274.230 698.810 274.250 ;
        RECT 700.370 274.230 700.840 274.550 ;
        RECT 701.010 274.470 706.700 274.610 ;
        RECT 718.580 274.570 724.270 274.710 ;
        RECT 735.750 274.740 736.130 274.790 ;
        RECT 737.400 274.740 737.910 274.970 ;
        RECT 753.560 274.800 753.940 274.850 ;
        RECT 755.210 274.800 755.720 275.030 ;
        RECT 758.870 274.800 759.250 274.860 ;
        RECT 741.060 274.740 741.440 274.800 ;
        RECT 701.010 274.350 701.390 274.470 ;
        RECT 691.000 274.030 691.380 274.110 ;
        RECT 692.770 274.100 693.830 274.110 ;
        RECT 686.380 273.970 690.710 274.030 ;
        RECT 639.090 273.390 639.520 273.450 ;
        RECT 686.520 273.440 687.110 273.970 ;
        RECT 692.770 273.730 693.550 274.100 ;
        RECT 696.370 274.090 700.840 274.230 ;
        RECT 702.660 274.150 703.170 274.470 ;
        RECT 706.320 274.360 706.700 274.470 ;
        RECT 703.750 274.180 704.340 274.280 ;
        RECT 707.730 274.180 707.970 274.400 ;
        RECT 698.210 273.860 698.810 274.090 ;
        RECT 700.370 274.000 700.840 274.090 ;
        RECT 703.610 274.050 707.970 274.180 ;
        RECT 708.230 274.280 708.610 274.340 ;
        RECT 710.020 274.280 711.020 274.540 ;
        RECT 715.780 274.330 716.380 274.350 ;
        RECT 717.990 274.330 718.430 274.550 ;
        RECT 718.580 274.450 718.960 274.570 ;
        RECT 708.230 274.130 711.020 274.280 ;
        RECT 713.940 274.190 718.430 274.330 ;
        RECT 720.230 274.250 720.740 274.570 ;
        RECT 723.890 274.460 724.270 274.570 ;
        RECT 721.320 274.280 721.910 274.380 ;
        RECT 725.300 274.280 725.540 274.500 ;
        RECT 708.230 274.050 708.610 274.130 ;
        RECT 703.610 273.990 707.940 274.050 ;
        RECT 703.750 273.460 704.340 273.990 ;
        RECT 710.020 273.640 711.020 274.130 ;
        RECT 715.780 273.960 716.380 274.190 ;
        RECT 717.990 274.170 718.430 274.190 ;
        RECT 718.010 274.150 718.270 274.170 ;
        RECT 721.180 274.150 725.540 274.280 ;
        RECT 725.800 274.380 726.180 274.440 ;
        RECT 727.550 274.380 728.510 274.670 ;
        RECT 735.750 274.600 741.440 274.740 ;
        RECT 735.180 274.540 735.440 274.550 ;
        RECT 725.800 274.230 728.510 274.380 ;
        RECT 732.950 274.360 733.550 274.380 ;
        RECT 735.120 274.360 735.550 274.540 ;
        RECT 735.750 274.480 736.130 274.600 ;
        RECT 725.800 274.150 726.180 274.230 ;
        RECT 721.180 274.090 725.510 274.150 ;
        RECT 721.320 273.560 721.910 274.090 ;
        RECT 727.550 273.870 728.510 274.230 ;
        RECT 731.110 274.220 735.550 274.360 ;
        RECT 737.400 274.280 737.910 274.600 ;
        RECT 741.060 274.490 741.440 274.600 ;
        RECT 738.490 274.310 739.080 274.410 ;
        RECT 742.470 274.310 742.710 274.530 ;
        RECT 732.950 273.990 733.550 274.220 ;
        RECT 735.120 274.200 735.550 274.220 ;
        RECT 735.180 274.180 735.440 274.200 ;
        RECT 738.350 274.180 742.710 274.310 ;
        RECT 742.970 274.410 743.350 274.470 ;
        RECT 744.860 274.410 746.050 274.800 ;
        RECT 753.560 274.660 759.250 274.800 ;
        RECT 752.990 274.580 753.250 274.610 ;
        RECT 750.760 274.420 751.360 274.440 ;
        RECT 752.920 274.420 753.400 274.580 ;
        RECT 753.560 274.540 753.940 274.660 ;
        RECT 742.970 274.260 746.050 274.410 ;
        RECT 748.920 274.280 753.400 274.420 ;
        RECT 755.210 274.340 755.720 274.660 ;
        RECT 758.870 274.550 759.250 274.660 ;
        RECT 760.780 274.470 761.160 274.530 ;
        RECT 762.570 274.470 763.640 274.890 ;
        RECT 851.870 274.800 852.620 275.390 ;
        RECT 742.970 274.180 743.350 274.260 ;
        RECT 738.350 274.120 742.680 274.180 ;
        RECT 738.490 273.590 739.080 274.120 ;
        RECT 744.860 273.840 746.050 274.260 ;
        RECT 750.760 274.050 751.360 274.280 ;
        RECT 752.920 274.260 753.400 274.280 ;
        RECT 760.780 274.320 763.640 274.470 ;
        RECT 752.990 274.240 753.250 274.260 ;
        RECT 760.780 274.240 761.160 274.320 ;
        RECT 762.570 273.950 763.640 274.320 ;
        RECT 795.880 274.110 796.200 274.350 ;
        RECT 797.480 274.110 798.460 274.450 ;
        RECT 795.880 273.890 798.460 274.110 ;
        RECT 814.760 274.420 815.080 274.670 ;
        RECT 815.770 274.420 816.700 274.580 ;
        RECT 814.760 274.200 816.700 274.420 ;
        RECT 814.760 273.960 815.080 274.200 ;
        RECT 795.880 273.610 796.200 273.890 ;
        RECT 797.480 273.620 798.460 273.890 ;
        RECT 815.770 273.810 816.700 274.200 ;
        RECT 833.610 274.330 833.940 274.470 ;
        RECT 834.550 274.330 835.120 274.600 ;
        RECT 833.610 274.040 835.120 274.330 ;
        RECT 833.610 273.750 833.940 274.040 ;
        RECT 834.550 274.030 835.120 274.040 ;
        RECT 782.975 273.515 783.265 273.560 ;
        RECT 785.375 273.515 785.665 273.560 ;
        RECT 790.655 273.515 790.945 273.560 ;
        RECT 629.350 273.270 629.580 273.290 ;
        RECT 621.980 272.250 622.670 272.340 ;
        RECT 621.600 272.210 622.670 272.250 ;
        RECT 608.420 268.370 608.680 271.920 ;
        RECT 609.220 270.750 609.870 270.970 ;
        RECT 609.220 270.720 610.370 270.750 ;
        RECT 609.220 270.570 613.500 270.720 ;
        RECT 609.220 270.400 610.370 270.570 ;
        RECT 611.670 270.400 611.890 270.570 ;
        RECT 613.270 270.400 613.490 270.570 ;
        RECT 610.090 270.240 610.330 270.400 ;
        RECT 610.090 270.020 610.320 270.240 ;
        RECT 610.880 270.020 611.110 270.400 ;
        RECT 611.670 270.020 611.900 270.400 ;
        RECT 612.460 270.020 612.690 270.400 ;
        RECT 613.250 270.230 613.490 270.400 ;
        RECT 613.250 270.020 613.480 270.230 ;
        RECT 610.100 268.930 610.280 270.020 ;
        RECT 610.900 268.930 611.080 270.020 ;
        RECT 611.700 268.930 611.880 270.020 ;
        RECT 612.480 268.930 612.660 270.020 ;
        RECT 613.260 268.930 613.440 270.020 ;
        RECT 615.360 269.910 615.580 272.170 ;
        RECT 620.930 272.070 622.670 272.210 ;
        RECT 620.930 271.970 621.440 272.070 ;
        RECT 621.600 271.960 622.670 272.070 ;
        RECT 620.910 270.690 621.390 270.760 ;
        RECT 617.680 270.540 621.390 270.690 ;
        RECT 617.700 270.370 617.920 270.540 ;
        RECT 619.260 270.370 619.480 270.540 ;
        RECT 620.860 270.480 621.390 270.540 ;
        RECT 620.860 270.370 621.080 270.480 ;
        RECT 617.680 270.210 617.920 270.370 ;
        RECT 617.680 269.990 617.910 270.210 ;
        RECT 618.470 269.990 618.700 270.370 ;
        RECT 619.260 269.990 619.490 270.370 ;
        RECT 620.050 269.990 620.280 270.370 ;
        RECT 620.840 270.200 621.080 270.370 ;
        RECT 620.840 269.990 621.070 270.200 ;
        RECT 615.230 269.490 615.710 269.910 ;
        RECT 613.920 269.040 617.340 269.180 ;
        RECT 610.090 268.550 610.320 268.930 ;
        RECT 610.880 268.550 611.110 268.930 ;
        RECT 611.670 268.550 611.900 268.930 ;
        RECT 612.460 268.550 612.690 268.930 ;
        RECT 613.250 268.550 613.480 268.930 ;
        RECT 613.950 268.880 614.140 269.040 ;
        RECT 615.510 268.880 615.700 269.040 ;
        RECT 617.120 268.880 617.310 269.040 ;
        RECT 617.690 268.900 617.870 269.990 ;
        RECT 618.490 268.900 618.670 269.990 ;
        RECT 619.290 268.900 619.470 269.990 ;
        RECT 620.070 268.900 620.250 269.990 ;
        RECT 620.850 268.900 621.030 269.990 ;
        RECT 608.240 268.060 608.910 268.370 ;
        RECT 609.510 267.720 609.660 267.730 ;
        RECT 601.410 267.470 603.250 267.630 ;
        RECT 606.320 267.580 609.750 267.720 ;
        RECT 603.090 266.820 603.240 267.470 ;
        RECT 606.360 267.410 606.510 267.580 ;
        RECT 607.950 267.410 608.100 267.580 ;
        RECT 609.510 267.410 609.660 267.580 ;
        RECT 610.100 267.460 610.280 268.550 ;
        RECT 610.900 267.460 611.080 268.550 ;
        RECT 611.700 267.460 611.880 268.550 ;
        RECT 612.480 267.460 612.660 268.550 ;
        RECT 613.260 267.460 613.440 268.550 ;
        RECT 613.920 268.500 614.150 268.880 ;
        RECT 615.500 268.500 615.730 268.880 ;
        RECT 617.080 268.500 617.310 268.880 ;
        RECT 617.680 268.520 617.910 268.900 ;
        RECT 618.470 268.520 618.700 268.900 ;
        RECT 619.260 268.520 619.490 268.900 ;
        RECT 620.050 268.520 620.280 268.900 ;
        RECT 620.840 268.520 621.070 268.900 ;
        RECT 606.340 267.030 606.570 267.410 ;
        RECT 607.130 267.030 607.360 267.410 ;
        RECT 607.920 267.030 608.150 267.410 ;
        RECT 608.710 267.030 608.940 267.410 ;
        RECT 609.500 267.030 609.730 267.410 ;
        RECT 610.090 267.080 610.320 267.460 ;
        RECT 610.880 267.290 611.110 267.460 ;
        RECT 610.870 267.080 611.110 267.290 ;
        RECT 611.670 267.080 611.900 267.460 ;
        RECT 612.460 267.080 612.690 267.460 ;
        RECT 613.250 267.080 613.480 267.460 ;
        RECT 613.940 267.410 614.100 268.500 ;
        RECT 615.520 267.410 615.680 268.500 ;
        RECT 617.100 267.410 617.260 268.500 ;
        RECT 617.690 267.430 617.870 268.520 ;
        RECT 618.490 267.430 618.670 268.520 ;
        RECT 619.290 267.430 619.470 268.520 ;
        RECT 620.070 267.430 620.250 268.520 ;
        RECT 620.850 267.430 621.030 268.520 ;
        RECT 621.600 267.720 621.810 271.960 ;
        RECT 621.980 271.880 622.670 271.960 ;
        RECT 623.030 268.500 623.260 273.210 ;
        RECT 626.260 273.120 629.590 273.270 ;
        RECT 629.350 270.810 629.580 273.120 ;
        RECT 639.070 272.940 639.540 273.390 ;
        RECT 782.975 273.375 790.945 273.515 ;
        RECT 782.975 273.330 783.265 273.375 ;
        RECT 785.375 273.330 785.665 273.375 ;
        RECT 790.655 273.330 790.945 273.375 ;
        RECT 801.865 273.505 802.155 273.550 ;
        RECT 804.265 273.505 804.555 273.550 ;
        RECT 809.545 273.505 809.835 273.550 ;
        RECT 801.865 273.365 809.835 273.505 ;
        RECT 801.865 273.320 802.155 273.365 ;
        RECT 804.265 273.320 804.555 273.365 ;
        RECT 809.545 273.320 809.835 273.365 ;
        RECT 820.715 273.475 821.005 273.520 ;
        RECT 823.115 273.475 823.405 273.520 ;
        RECT 828.395 273.475 828.685 273.520 ;
        RECT 820.715 273.335 828.685 273.475 ;
        RECT 820.715 273.290 821.005 273.335 ;
        RECT 823.115 273.290 823.405 273.335 ;
        RECT 828.395 273.290 828.685 273.335 ;
        RECT 645.150 273.160 645.520 273.220 ;
        RECT 639.090 272.880 639.520 272.940 ;
        RECT 645.130 272.810 645.540 273.160 ;
        RECT 645.150 272.750 645.520 272.810 ;
        RECT 631.440 271.070 632.060 271.730 ;
        RECT 633.680 271.690 634.510 272.430 ;
        RECT 641.540 272.350 642.040 272.730 ;
        RECT 803.270 272.690 803.610 272.750 ;
        RECT 784.340 272.600 784.730 272.660 ;
        RECT 784.320 272.250 784.750 272.600 ;
        RECT 784.340 272.190 784.730 272.250 ;
        RECT 803.250 272.240 803.630 272.690 ;
        RECT 822.110 272.660 822.450 272.720 ;
        RECT 822.090 272.280 822.470 272.660 ;
        RECT 834.710 272.380 834.870 274.030 ;
        RECT 836.970 273.720 837.500 274.050 ;
        RECT 839.220 273.720 839.510 273.970 ;
        RECT 852.100 273.810 852.380 274.800 ;
        RECT 836.970 273.570 839.510 273.720 ;
        RECT 836.970 273.510 839.430 273.570 ;
        RECT 836.970 273.440 837.500 273.510 ;
        RECT 841.830 273.190 842.160 273.520 ;
        RECT 843.270 273.190 843.430 273.200 ;
        RECT 836.720 273.000 837.510 273.080 ;
        RECT 839.800 273.000 840.230 273.080 ;
        RECT 836.720 272.800 840.230 273.000 ;
        RECT 841.830 273.020 843.430 273.190 ;
        RECT 841.830 272.820 842.160 273.020 ;
        RECT 836.720 272.780 840.010 272.800 ;
        RECT 836.720 272.660 837.510 272.780 ;
        RECT 834.700 272.370 837.320 272.380 ;
        RECT 838.960 272.370 839.380 272.560 ;
        RECT 803.270 272.180 803.610 272.240 ;
        RECT 822.110 272.220 822.450 272.280 ;
        RECT 834.700 272.210 839.380 272.370 ;
        RECT 834.700 272.200 839.200 272.210 ;
        RECT 834.700 272.180 837.320 272.200 ;
        RECT 628.980 270.460 629.580 270.810 ;
        RECT 629.350 270.080 629.580 270.460 ;
        RECT 638.980 270.290 639.680 270.650 ;
        RECT 627.440 269.920 630.820 270.080 ;
        RECT 627.450 269.750 627.620 269.920 ;
        RECT 629.020 269.750 629.190 269.920 ;
        RECT 629.350 269.910 629.580 269.920 ;
        RECT 630.620 269.750 630.790 269.920 ;
        RECT 627.420 269.370 627.650 269.750 ;
        RECT 628.210 269.370 628.440 269.750 ;
        RECT 629.000 269.370 629.230 269.750 ;
        RECT 629.790 269.370 630.020 269.750 ;
        RECT 630.580 269.370 630.810 269.750 ;
        RECT 622.830 267.950 623.520 268.500 ;
        RECT 627.450 268.280 627.630 269.370 ;
        RECT 628.230 268.280 628.410 269.370 ;
        RECT 629.020 268.280 629.200 269.370 ;
        RECT 629.800 268.280 629.980 269.370 ;
        RECT 630.590 268.280 630.770 269.370 ;
        RECT 627.420 267.900 627.650 268.280 ;
        RECT 628.210 267.900 628.440 268.280 ;
        RECT 629.000 267.900 629.230 268.280 ;
        RECT 629.790 267.900 630.020 268.280 ;
        RECT 630.580 267.900 630.810 268.280 ;
        RECT 639.240 267.990 639.420 270.290 ;
        RECT 643.080 270.170 643.650 270.850 ;
        RECT 822.040 270.490 822.570 270.920 ;
        RECT 843.270 270.910 843.430 273.020 ;
        RECT 851.970 272.770 852.560 273.810 ;
        RECT 853.130 272.080 853.350 277.560 ;
        RECT 853.860 272.430 854.120 283.350 ;
        RECT 860.200 283.010 860.390 284.450 ;
        RECT 861.830 283.010 862.100 283.050 ;
        RECT 860.200 282.840 862.100 283.010 ;
        RECT 861.830 282.650 862.100 282.840 ;
        RECT 862.790 282.470 863.100 282.860 ;
        RECT 865.100 282.640 865.970 283.200 ;
        RECT 860.180 282.330 860.410 282.340 ;
        RECT 862.820 282.330 863.050 282.470 ;
        RECT 860.180 282.130 863.050 282.330 ;
        RECT 865.360 282.220 865.670 282.640 ;
        RECT 865.190 282.160 866.010 282.220 ;
        RECT 858.890 280.860 859.200 280.970 ;
        RECT 860.180 280.860 860.410 282.130 ;
        RECT 862.820 282.120 863.050 282.130 ;
        RECT 865.170 281.200 866.030 282.160 ;
        RECT 865.190 281.140 866.010 281.200 ;
        RECT 858.890 280.710 860.410 280.860 ;
        RECT 858.890 280.700 860.350 280.710 ;
        RECT 858.890 280.570 859.200 280.700 ;
        RECT 857.010 279.290 857.370 279.350 ;
        RECT 856.990 278.860 857.390 279.290 ;
        RECT 857.010 278.800 857.370 278.860 ;
        RECT 856.950 272.430 857.420 272.530 ;
        RECT 853.860 272.200 857.420 272.430 ;
        RECT 852.950 271.510 853.550 272.080 ;
        RECT 844.720 270.910 845.230 271.060 ;
        RECT 843.270 270.740 845.230 270.910 ;
        RECT 844.720 270.680 845.230 270.740 ;
        RECT 852.430 270.870 852.970 271.150 ;
        RECT 853.860 270.870 854.120 272.200 ;
        RECT 856.950 272.170 857.420 272.200 ;
        RECT 852.430 270.590 854.160 270.870 ;
        RECT 639.560 268.390 640.010 269.080 ;
        RECT 643.310 268.040 643.450 270.170 ;
        RECT 717.700 269.760 717.960 269.850 ;
        RECT 724.390 269.760 725.640 269.820 ;
        RECT 682.900 269.640 683.160 269.730 ;
        RECT 689.590 269.640 690.840 269.700 ;
        RECT 682.900 269.420 690.840 269.640 ;
        RECT 682.900 269.280 683.160 269.420 ;
        RECT 689.590 269.410 690.840 269.420 ;
        RECT 700.130 269.660 700.390 269.750 ;
        RECT 706.820 269.660 708.070 269.720 ;
        RECT 700.130 269.440 708.070 269.660 ;
        RECT 717.700 269.540 725.640 269.760 ;
        RECT 643.620 268.930 644.040 269.130 ;
        RECT 645.050 268.930 646.030 269.240 ;
        RECT 643.620 268.720 646.030 268.930 ;
        RECT 688.570 268.820 688.890 268.970 ;
        RECT 643.620 268.450 644.040 268.720 ;
        RECT 645.050 268.460 646.030 268.720 ;
        RECT 685.770 268.710 686.060 268.750 ;
        RECT 679.980 268.220 680.490 268.660 ;
        RECT 680.050 268.200 680.410 268.220 ;
        RECT 628.230 267.760 628.410 267.900 ;
        RECT 629.820 267.760 630.000 267.900 ;
        RECT 639.240 267.880 639.500 267.990 ;
        RECT 624.600 267.720 624.750 267.730 ;
        RECT 621.410 267.580 624.840 267.720 ;
        RECT 628.190 267.600 630.030 267.760 ;
        RECT 639.270 267.610 639.500 267.880 ;
        RECT 643.310 267.870 643.550 268.040 ;
        RECT 680.930 267.980 681.390 268.490 ;
        RECT 685.720 268.230 686.150 268.710 ;
        RECT 688.570 268.680 689.770 268.820 ;
        RECT 690.660 268.740 690.830 269.410 ;
        RECT 700.130 269.300 700.390 269.440 ;
        RECT 706.820 269.430 708.070 269.440 ;
        RECT 694.040 268.850 695.520 268.880 ;
        RECT 686.650 268.430 687.070 268.490 ;
        RECT 688.570 268.460 688.890 268.680 ;
        RECT 643.320 267.660 643.550 267.870 ;
        RECT 686.630 267.850 687.090 268.430 ;
        RECT 689.610 268.240 689.760 268.680 ;
        RECT 690.660 268.660 692.610 268.740 ;
        RECT 690.660 268.560 692.820 268.660 ;
        RECT 691.470 268.240 691.880 268.390 ;
        RECT 692.410 268.330 692.820 268.560 ;
        RECT 693.910 268.600 695.520 268.850 ;
        RECT 705.800 268.840 706.120 268.990 ;
        RECT 703.000 268.730 703.290 268.770 ;
        RECT 693.910 268.470 694.160 268.600 ;
        RECT 689.610 268.060 691.880 268.240 ;
        RECT 689.610 268.040 691.720 268.060 ;
        RECT 698.160 268.000 698.620 268.510 ;
        RECT 702.950 268.250 703.380 268.730 ;
        RECT 705.800 268.700 707.000 268.840 ;
        RECT 707.890 268.760 708.060 269.430 ;
        RECT 711.040 268.900 711.500 269.540 ;
        RECT 717.700 269.400 717.960 269.540 ;
        RECT 724.390 269.530 725.640 269.540 ;
        RECT 734.870 269.790 735.130 269.880 ;
        RECT 752.680 269.850 752.940 269.940 ;
        RECT 759.370 269.850 760.620 269.910 ;
        RECT 741.560 269.790 742.810 269.850 ;
        RECT 734.870 269.570 742.810 269.790 ;
        RECT 723.370 268.940 723.690 269.090 ;
        RECT 703.880 268.450 704.300 268.510 ;
        RECT 705.800 268.480 706.120 268.700 ;
        RECT 703.860 267.870 704.320 268.450 ;
        RECT 706.840 268.260 706.990 268.700 ;
        RECT 707.890 268.680 709.840 268.760 ;
        RECT 711.040 268.740 712.750 268.900 ;
        RECT 720.570 268.830 720.860 268.870 ;
        RECT 707.890 268.580 710.050 268.680 ;
        RECT 708.700 268.260 709.110 268.410 ;
        RECT 709.640 268.350 710.050 268.580 ;
        RECT 711.140 268.620 712.750 268.740 ;
        RECT 711.140 268.490 711.390 268.620 ;
        RECT 706.840 268.080 709.110 268.260 ;
        RECT 715.730 268.100 716.190 268.610 ;
        RECT 720.520 268.350 720.950 268.830 ;
        RECT 723.370 268.800 724.570 268.940 ;
        RECT 725.460 268.860 725.630 269.530 ;
        RECT 734.870 269.430 735.130 269.570 ;
        RECT 741.560 269.560 742.810 269.570 ;
        RECT 728.840 268.970 730.320 269.000 ;
        RECT 721.450 268.550 721.870 268.610 ;
        RECT 723.370 268.580 723.690 268.800 ;
        RECT 706.840 268.060 708.950 268.080 ;
        RECT 721.430 267.970 721.890 268.550 ;
        RECT 724.410 268.360 724.560 268.800 ;
        RECT 725.460 268.780 727.410 268.860 ;
        RECT 728.710 268.780 730.320 268.970 ;
        RECT 740.540 268.970 740.860 269.120 ;
        RECT 737.740 268.860 738.030 268.900 ;
        RECT 725.460 268.680 727.620 268.780 ;
        RECT 726.270 268.360 726.680 268.510 ;
        RECT 727.210 268.450 727.620 268.680 ;
        RECT 728.590 268.720 730.320 268.780 ;
        RECT 724.410 268.180 726.680 268.360 ;
        RECT 724.410 268.160 726.520 268.180 ;
        RECT 721.450 267.910 721.870 267.970 ;
        RECT 728.590 267.920 729.120 268.720 ;
        RECT 732.900 268.130 733.360 268.640 ;
        RECT 737.690 268.380 738.120 268.860 ;
        RECT 740.540 268.830 741.740 268.970 ;
        RECT 742.630 268.890 742.800 269.560 ;
        RECT 745.810 269.030 746.220 269.780 ;
        RECT 752.680 269.630 760.620 269.850 ;
        RECT 752.680 269.490 752.940 269.630 ;
        RECT 759.370 269.620 760.620 269.630 ;
        RECT 758.350 269.030 758.670 269.180 ;
        RECT 738.620 268.580 739.040 268.640 ;
        RECT 740.540 268.610 740.860 268.830 ;
        RECT 738.600 268.000 739.060 268.580 ;
        RECT 741.580 268.390 741.730 268.830 ;
        RECT 742.630 268.810 744.580 268.890 ;
        RECT 745.810 268.880 747.490 269.030 ;
        RECT 755.550 268.920 755.840 268.960 ;
        RECT 742.630 268.710 744.790 268.810 ;
        RECT 743.440 268.390 743.850 268.540 ;
        RECT 744.380 268.480 744.790 268.710 ;
        RECT 745.880 268.750 747.490 268.880 ;
        RECT 745.880 268.620 746.130 268.750 ;
        RECT 741.580 268.210 743.850 268.390 ;
        RECT 741.580 268.190 743.690 268.210 ;
        RECT 750.710 268.190 751.170 268.700 ;
        RECT 755.500 268.440 755.930 268.920 ;
        RECT 758.350 268.890 759.550 269.030 ;
        RECT 760.440 268.950 760.610 269.620 ;
        RECT 763.820 269.060 765.300 269.090 ;
        RECT 758.350 268.670 758.670 268.890 ;
        RECT 759.390 268.450 759.540 268.890 ;
        RECT 760.440 268.870 762.390 268.950 ;
        RECT 763.690 268.940 765.300 269.060 ;
        RECT 760.440 268.770 762.600 268.870 ;
        RECT 761.250 268.450 761.660 268.600 ;
        RECT 762.190 268.540 762.600 268.770 ;
        RECT 763.620 268.810 765.300 268.940 ;
        RECT 759.390 268.270 761.660 268.450 ;
        RECT 763.620 268.280 764.070 268.810 ;
        RECT 759.390 268.250 761.500 268.270 ;
        RECT 822.070 268.190 822.420 270.490 ;
        RECT 852.430 270.450 852.970 270.590 ;
        RECT 845.700 270.210 846.170 270.370 ;
        RECT 843.230 270.190 846.170 270.210 ;
        RECT 843.220 270.000 846.170 270.190 ;
        RECT 843.220 269.980 845.950 270.000 ;
        RECT 822.070 268.170 830.050 268.190 ;
        RECT 738.620 267.940 739.040 268.000 ;
        RECT 822.070 267.900 830.090 268.170 ;
        RECT 686.650 267.790 687.070 267.850 ;
        RECT 703.880 267.810 704.300 267.870 ;
        RECT 607.170 266.880 607.320 267.030 ;
        RECT 608.750 266.880 608.900 267.030 ;
        RECT 610.130 266.880 610.310 267.080 ;
        RECT 591.710 264.660 591.960 266.155 ;
        RECT 601.360 266.090 602.710 266.600 ;
        RECT 603.010 266.380 603.460 266.820 ;
        RECT 607.120 266.730 610.310 266.880 ;
        RECT 610.870 266.920 611.040 267.080 ;
        RECT 612.470 266.920 612.640 267.080 ;
        RECT 613.920 267.030 614.150 267.410 ;
        RECT 615.500 267.030 615.730 267.410 ;
        RECT 617.080 267.030 617.310 267.410 ;
        RECT 617.680 267.050 617.910 267.430 ;
        RECT 618.470 267.260 618.700 267.430 ;
        RECT 618.460 267.050 618.700 267.260 ;
        RECT 619.260 267.050 619.490 267.430 ;
        RECT 620.050 267.050 620.280 267.430 ;
        RECT 620.840 267.250 621.070 267.430 ;
        RECT 621.450 267.410 621.600 267.580 ;
        RECT 623.040 267.410 623.190 267.580 ;
        RECT 624.600 267.410 624.750 267.580 ;
        RECT 620.840 267.050 621.080 267.250 ;
        RECT 613.920 266.920 614.120 267.030 ;
        RECT 610.870 266.810 614.120 266.920 ;
        RECT 608.890 266.700 610.310 266.730 ;
        RECT 610.810 266.780 614.120 266.810 ;
        RECT 610.810 266.770 612.710 266.780 ;
        RECT 610.810 266.470 611.220 266.770 ;
        RECT 613.920 266.410 614.120 266.780 ;
        RECT 617.090 266.880 617.310 267.030 ;
        RECT 618.460 266.890 618.630 267.050 ;
        RECT 620.060 266.890 620.230 267.050 ;
        RECT 618.460 266.880 620.300 266.890 ;
        RECT 617.090 266.800 620.300 266.880 ;
        RECT 620.880 266.840 621.080 267.050 ;
        RECT 621.430 267.030 621.660 267.410 ;
        RECT 622.220 267.030 622.450 267.410 ;
        RECT 623.010 267.030 623.240 267.410 ;
        RECT 623.800 267.030 624.030 267.410 ;
        RECT 624.590 267.030 624.820 267.410 ;
        RECT 622.260 266.880 622.410 267.030 ;
        RECT 623.840 266.880 623.990 267.030 ;
        RECT 622.210 266.840 624.030 266.880 ;
        RECT 617.090 266.740 620.340 266.800 ;
        RECT 617.090 266.710 618.850 266.740 ;
        RECT 619.940 266.440 620.340 266.740 ;
        RECT 620.880 266.730 624.030 266.840 ;
        RECT 620.880 266.680 622.370 266.730 ;
        RECT 628.930 266.250 629.140 267.600 ;
        RECT 795.870 266.970 796.190 267.130 ;
        RECT 797.500 266.970 798.450 267.290 ;
        RECT 795.870 266.740 798.450 266.970 ;
        RECT 795.870 266.420 796.190 266.740 ;
        RECT 797.500 266.530 798.450 266.740 ;
        RECT 814.400 266.820 814.730 267.000 ;
        RECT 816.080 266.820 817.030 267.190 ;
        RECT 814.400 266.630 817.030 266.820 ;
        RECT 814.400 266.400 814.730 266.630 ;
        RECT 816.080 266.430 817.030 266.630 ;
        RECT 628.760 265.900 629.380 266.250 ;
        RECT 801.515 266.015 801.805 266.060 ;
        RECT 803.915 266.015 804.205 266.060 ;
        RECT 809.195 266.015 809.485 266.060 ;
        RECT 782.985 265.955 783.275 266.000 ;
        RECT 785.385 265.955 785.675 266.000 ;
        RECT 790.665 265.955 790.955 266.000 ;
        RECT 782.985 265.815 790.955 265.955 ;
        RECT 801.515 265.875 809.485 266.015 ;
        RECT 801.515 265.830 801.805 265.875 ;
        RECT 803.915 265.830 804.205 265.875 ;
        RECT 809.195 265.830 809.485 265.875 ;
        RECT 782.985 265.770 783.275 265.815 ;
        RECT 785.385 265.770 785.675 265.815 ;
        RECT 790.665 265.770 790.955 265.815 ;
        RECT 784.390 265.150 784.730 265.210 ;
        RECT 802.920 265.180 803.250 265.240 ;
        RECT 784.370 264.740 784.750 265.150 ;
        RECT 802.900 264.780 803.270 265.180 ;
        RECT 379.130 263.380 379.360 264.360 ;
        RECT 385.710 263.380 385.940 264.360 ;
        RECT 591.050 263.590 592.560 264.660 ;
        RECT 692.350 264.440 693.980 264.700 ;
        RECT 784.390 264.680 784.730 264.740 ;
        RECT 802.920 264.720 803.250 264.780 ;
        RECT 678.230 263.890 693.980 264.440 ;
        RECT 379.130 259.910 379.360 260.890 ;
        RECT 385.710 259.910 385.940 260.890 ;
        RECT 632.160 259.980 633.650 260.970 ;
        RECT 602.960 258.520 603.190 258.900 ;
        RECT 604.540 258.520 604.770 258.900 ;
        RECT 607.480 258.530 607.710 258.910 ;
        RECT 609.060 258.530 609.290 258.910 ;
        RECT 612.000 258.530 612.230 258.910 ;
        RECT 613.580 258.530 613.810 258.910 ;
        RECT 602.980 257.430 603.160 258.520 ;
        RECT 604.550 257.430 604.730 258.520 ;
        RECT 607.500 257.440 607.680 258.530 ;
        RECT 609.070 257.440 609.250 258.530 ;
        RECT 612.020 257.440 612.200 258.530 ;
        RECT 613.590 257.440 613.770 258.530 ;
        RECT 616.430 258.510 616.660 258.890 ;
        RECT 618.010 258.510 618.240 258.890 ;
        RECT 620.810 258.520 621.040 258.900 ;
        RECT 622.390 258.520 622.620 258.900 ;
        RECT 379.130 256.440 379.360 257.420 ;
        RECT 385.710 256.440 385.940 257.420 ;
        RECT 602.960 257.270 603.190 257.430 ;
        RECT 602.910 256.910 603.190 257.270 ;
        RECT 604.540 257.050 604.770 257.430 ;
        RECT 607.480 257.060 607.710 257.440 ;
        RECT 609.060 257.060 609.290 257.440 ;
        RECT 612.000 257.060 612.230 257.440 ;
        RECT 613.580 257.060 613.810 257.440 ;
        RECT 616.450 257.420 616.630 258.510 ;
        RECT 618.020 257.420 618.200 258.510 ;
        RECT 620.830 257.430 621.010 258.520 ;
        RECT 622.400 257.430 622.580 258.520 ;
        RECT 625.130 258.510 625.360 258.890 ;
        RECT 626.710 258.510 626.940 258.890 ;
        RECT 678.230 258.710 678.530 263.890 ;
        RECT 692.350 263.500 693.980 263.890 ;
        RECT 829.540 260.970 830.090 267.900 ;
        RECT 841.390 267.970 841.700 268.150 ;
        RECT 843.220 267.970 843.410 269.980 ;
        RECT 836.850 267.670 837.420 267.820 ;
        RECT 841.390 267.740 843.410 267.970 ;
        RECT 836.850 267.660 838.620 267.670 ;
        RECT 836.850 267.460 838.990 267.660 ;
        RECT 836.850 267.400 837.420 267.460 ;
        RECT 838.470 267.330 838.990 267.460 ;
        RECT 841.390 267.410 841.700 267.740 ;
        RECT 843.220 267.730 843.410 267.740 ;
        RECT 839.490 267.080 839.840 267.140 ;
        RECT 839.470 266.690 839.860 267.080 ;
        RECT 850.820 267.000 851.750 267.670 ;
        RECT 839.490 266.630 839.840 266.690 ;
        RECT 851.050 262.270 851.380 267.000 ;
        RECT 852.670 262.420 852.880 270.450 ;
        RECT 862.750 269.160 863.120 269.440 ;
        RECT 862.840 268.990 863.030 269.160 ;
        RECT 860.050 268.960 863.030 268.990 ;
        RECT 860.050 268.810 863.020 268.960 ;
        RECT 865.320 268.810 866.830 270.060 ;
        RECT 858.950 267.640 859.290 267.780 ;
        RECT 860.050 267.640 860.290 268.810 ;
        RECT 858.950 267.450 860.290 267.640 ;
        RECT 858.950 267.270 859.290 267.450 ;
        RECT 860.050 267.440 860.290 267.450 ;
        RECT 853.550 265.770 854.120 265.990 ;
        RECT 857.090 265.770 857.470 266.010 ;
        RECT 853.550 265.570 857.470 265.770 ;
        RECT 853.550 265.500 854.120 265.570 ;
        RECT 857.090 265.510 857.470 265.570 ;
        RECT 853.080 264.990 853.630 265.310 ;
        RECT 853.080 264.790 853.720 264.990 ;
        RECT 850.820 261.510 851.850 262.270 ;
        RECT 852.470 261.780 853.260 262.420 ;
        RECT 853.490 261.650 853.720 264.790 ;
        RECT 853.350 261.220 853.920 261.650 ;
        RECT 866.170 260.970 866.540 268.810 ;
        RECT 829.540 260.560 866.540 260.970 ;
        RECT 846.570 258.970 847.500 259.290 ;
        RECT 853.310 258.970 853.940 259.230 ;
        RECT 679.930 258.710 680.350 258.780 ;
        RECT 604.570 256.910 604.750 257.050 ;
        RECT 607.500 256.920 607.700 257.060 ;
        RECT 609.090 256.920 609.270 257.060 ;
        RECT 612.020 256.920 612.200 257.060 ;
        RECT 613.610 256.920 613.790 257.060 ;
        RECT 616.430 257.040 616.660 257.420 ;
        RECT 618.010 257.040 618.240 257.420 ;
        RECT 620.810 257.050 621.040 257.430 ;
        RECT 622.390 257.050 622.620 257.430 ;
        RECT 625.150 257.420 625.330 258.510 ;
        RECT 626.720 257.420 626.900 258.510 ;
        RECT 678.230 258.480 680.350 258.710 ;
        RECT 846.570 258.740 853.940 258.970 ;
        RECT 846.570 258.710 853.540 258.740 ;
        RECT 678.230 258.470 680.180 258.480 ;
        RECT 694.430 258.330 695.140 258.420 ;
        RECT 700.030 258.330 700.440 258.440 ;
        RECT 694.430 258.140 700.440 258.330 ;
        RECT 712.700 258.290 713.540 258.400 ;
        RECT 717.820 258.290 718.180 258.420 ;
        RECT 683.120 257.580 683.710 258.080 ;
        RECT 694.430 258.010 700.150 258.140 ;
        RECT 694.430 257.790 695.140 258.010 ;
        RECT 700.620 258.000 701.130 258.190 ;
        RECT 700.510 257.540 701.130 258.000 ;
        RECT 712.700 258.150 718.180 258.290 ;
        RECT 729.880 258.310 730.750 258.420 ;
        RECT 735.060 258.310 735.420 258.450 ;
        RECT 729.880 258.180 735.420 258.310 ;
        RECT 747.450 258.270 748.360 258.420 ;
        RECT 752.540 258.270 752.900 258.410 ;
        RECT 712.700 258.080 717.960 258.150 ;
        RECT 712.700 257.840 713.540 258.080 ;
        RECT 729.880 258.040 735.220 258.180 ;
        RECT 747.450 258.140 752.900 258.270 ;
        RECT 846.570 258.190 847.500 258.710 ;
        RECT 700.620 257.490 701.130 257.540 ;
        RECT 718.200 257.520 718.740 257.970 ;
        RECT 729.880 257.790 730.750 258.040 ;
        RECT 747.450 258.020 752.780 258.140 ;
        RECT 735.520 257.960 735.910 258.020 ;
        RECT 735.500 257.620 735.930 257.960 ;
        RECT 747.450 257.790 748.360 258.020 ;
        RECT 735.520 257.560 735.910 257.620 ;
        RECT 752.930 257.570 753.430 257.950 ;
        RECT 602.910 256.750 604.780 256.910 ;
        RECT 607.460 256.900 609.300 256.920 ;
        RECT 611.980 256.900 613.820 256.920 ;
        RECT 616.450 256.900 616.630 257.040 ;
        RECT 618.040 256.900 618.220 257.040 ;
        RECT 620.830 256.910 621.010 257.050 ;
        RECT 622.420 256.910 622.600 257.050 ;
        RECT 625.130 257.040 625.360 257.420 ;
        RECT 626.710 257.040 626.940 257.420 ;
        RECT 620.790 256.900 622.630 256.910 ;
        RECT 625.150 256.900 625.330 257.040 ;
        RECT 626.740 256.900 626.920 257.040 ;
        RECT 607.460 256.830 615.140 256.900 ;
        RECT 607.460 256.760 615.150 256.830 ;
        RECT 602.910 255.390 603.190 256.750 ;
        RECT 607.530 255.740 607.700 256.760 ;
        RECT 613.500 256.740 615.150 256.760 ;
        RECT 616.410 256.760 622.630 256.900 ;
        RECT 616.410 256.740 618.250 256.760 ;
        RECT 620.790 256.750 622.630 256.760 ;
        RECT 613.080 256.080 613.550 256.460 ;
        RECT 614.940 256.290 615.150 256.740 ;
        RECT 615.920 256.290 616.350 256.360 ;
        RECT 614.940 256.110 616.350 256.290 ;
        RECT 608.120 255.740 608.790 256.050 ;
        RECT 607.520 255.460 608.790 255.740 ;
        RECT 386.610 255.110 388.450 255.270 ;
        RECT 596.690 255.160 597.380 255.220 ;
        RECT 386.470 253.990 388.450 255.110 ;
        RECT 593.980 254.660 594.780 255.120 ;
        RECT 299.360 249.250 340.190 252.160 ;
        RECT 299.530 249.070 301.590 249.250 ;
        RECT 334.070 232.800 336.270 233.440 ;
        RECT 332.750 232.650 336.270 232.800 ;
        RECT 330.860 231.210 336.270 232.650 ;
        RECT 332.750 230.790 336.270 231.210 ;
        RECT 334.070 229.870 336.270 230.790 ;
        RECT 339.090 218.140 340.190 249.250 ;
        RECT 378.610 241.100 382.040 243.480 ;
        RECT 379.800 238.950 380.990 241.100 ;
        RECT 386.470 240.010 388.100 253.990 ;
        RECT 594.120 253.140 594.400 254.660 ;
        RECT 596.670 254.310 597.400 255.160 ;
        RECT 596.690 254.250 597.380 254.310 ;
        RECT 593.880 252.870 594.610 253.140 ;
        RECT 602.900 253.120 603.210 255.390 ;
        RECT 607.530 255.090 607.700 255.460 ;
        RECT 608.120 255.200 608.790 255.460 ;
        RECT 613.170 255.560 613.410 256.080 ;
        RECT 615.920 256.040 616.350 256.110 ;
        RECT 616.730 255.560 616.910 256.740 ;
        RECT 620.330 256.340 620.740 256.610 ;
        RECT 620.280 256.180 620.740 256.340 ;
        RECT 620.280 256.040 620.700 256.180 ;
        RECT 613.170 255.400 616.920 255.560 ;
        RECT 606.790 254.450 607.700 255.090 ;
        RECT 615.210 254.670 615.430 254.730 ;
        RECT 620.280 254.670 620.550 256.040 ;
        RECT 603.500 253.120 604.460 253.290 ;
        RECT 602.840 252.840 604.460 253.120 ;
        RECT 602.900 252.220 603.210 252.840 ;
        RECT 603.500 252.730 604.460 252.840 ;
        RECT 600.510 252.060 603.890 252.220 ;
        RECT 600.520 251.890 600.690 252.060 ;
        RECT 602.090 251.890 602.260 252.060 ;
        RECT 603.690 251.890 603.860 252.060 ;
        RECT 591.190 250.160 592.240 251.600 ;
        RECT 600.490 251.510 600.720 251.890 ;
        RECT 601.280 251.510 601.510 251.890 ;
        RECT 602.070 251.510 602.300 251.890 ;
        RECT 602.860 251.510 603.090 251.890 ;
        RECT 603.650 251.510 603.880 251.890 ;
        RECT 600.520 250.420 600.700 251.510 ;
        RECT 601.300 250.420 601.480 251.510 ;
        RECT 602.090 250.420 602.270 251.510 ;
        RECT 602.870 250.420 603.050 251.510 ;
        RECT 603.660 250.420 603.840 251.510 ;
        RECT 591.480 248.405 591.730 250.160 ;
        RECT 600.490 250.040 600.720 250.420 ;
        RECT 601.280 250.040 601.510 250.420 ;
        RECT 602.070 250.040 602.300 250.420 ;
        RECT 602.860 250.040 603.090 250.420 ;
        RECT 603.650 250.040 603.880 250.420 ;
        RECT 601.300 249.900 601.480 250.040 ;
        RECT 602.890 249.900 603.070 250.040 ;
        RECT 607.530 249.990 607.700 254.450 ;
        RECT 608.100 254.190 608.740 254.610 ;
        RECT 615.210 254.440 620.550 254.670 ;
        RECT 620.780 254.480 621.290 254.530 ;
        RECT 621.450 254.520 621.660 256.750 ;
        RECT 625.110 256.740 626.950 256.900 ;
        RECT 622.650 255.480 623.500 255.920 ;
        RECT 626.110 255.540 626.330 256.740 ;
        RECT 855.980 256.680 856.430 257.040 ;
        RECT 858.820 256.840 859.130 257.110 ;
        RECT 858.820 256.830 860.270 256.840 ;
        RECT 751.620 256.260 752.300 256.320 ;
        RECT 850.920 256.260 851.720 256.640 ;
        RECT 856.950 256.460 857.360 256.670 ;
        RECT 858.820 256.660 860.450 256.830 ;
        RECT 858.820 256.480 859.130 256.660 ;
        RECT 751.620 255.920 851.720 256.260 ;
        RECT 852.910 256.220 857.360 256.460 ;
        RECT 751.620 255.720 752.300 255.920 ;
        RECT 850.920 255.760 851.720 255.920 ;
        RECT 638.940 255.660 639.370 255.720 ;
        RECT 629.200 255.540 629.430 255.560 ;
        RECT 621.830 254.520 622.520 254.610 ;
        RECT 621.450 254.480 622.520 254.520 ;
        RECT 608.270 250.640 608.530 254.190 ;
        RECT 609.070 253.020 609.720 253.240 ;
        RECT 609.070 252.990 610.220 253.020 ;
        RECT 609.070 252.840 613.350 252.990 ;
        RECT 609.070 252.670 610.220 252.840 ;
        RECT 611.520 252.670 611.740 252.840 ;
        RECT 613.120 252.670 613.340 252.840 ;
        RECT 609.940 252.510 610.180 252.670 ;
        RECT 609.940 252.290 610.170 252.510 ;
        RECT 610.730 252.290 610.960 252.670 ;
        RECT 611.520 252.290 611.750 252.670 ;
        RECT 612.310 252.290 612.540 252.670 ;
        RECT 613.100 252.500 613.340 252.670 ;
        RECT 613.100 252.290 613.330 252.500 ;
        RECT 609.950 251.200 610.130 252.290 ;
        RECT 610.750 251.200 610.930 252.290 ;
        RECT 611.550 251.200 611.730 252.290 ;
        RECT 612.330 251.200 612.510 252.290 ;
        RECT 613.110 251.200 613.290 252.290 ;
        RECT 615.210 252.180 615.430 254.440 ;
        RECT 620.780 254.340 622.520 254.480 ;
        RECT 620.780 254.240 621.290 254.340 ;
        RECT 621.450 254.230 622.520 254.340 ;
        RECT 620.760 252.960 621.240 253.030 ;
        RECT 617.530 252.810 621.240 252.960 ;
        RECT 617.550 252.640 617.770 252.810 ;
        RECT 619.110 252.640 619.330 252.810 ;
        RECT 620.710 252.750 621.240 252.810 ;
        RECT 620.710 252.640 620.930 252.750 ;
        RECT 617.530 252.480 617.770 252.640 ;
        RECT 617.530 252.260 617.760 252.480 ;
        RECT 618.320 252.260 618.550 252.640 ;
        RECT 619.110 252.260 619.340 252.640 ;
        RECT 619.900 252.260 620.130 252.640 ;
        RECT 620.690 252.470 620.930 252.640 ;
        RECT 620.690 252.260 620.920 252.470 ;
        RECT 615.080 251.760 615.560 252.180 ;
        RECT 613.770 251.310 617.190 251.450 ;
        RECT 609.940 250.820 610.170 251.200 ;
        RECT 610.730 250.820 610.960 251.200 ;
        RECT 611.520 250.820 611.750 251.200 ;
        RECT 612.310 250.820 612.540 251.200 ;
        RECT 613.100 250.820 613.330 251.200 ;
        RECT 613.800 251.150 613.990 251.310 ;
        RECT 615.360 251.150 615.550 251.310 ;
        RECT 616.970 251.150 617.160 251.310 ;
        RECT 617.540 251.170 617.720 252.260 ;
        RECT 618.340 251.170 618.520 252.260 ;
        RECT 619.140 251.170 619.320 252.260 ;
        RECT 619.920 251.170 620.100 252.260 ;
        RECT 620.700 251.170 620.880 252.260 ;
        RECT 608.090 250.330 608.760 250.640 ;
        RECT 609.360 249.990 609.510 250.000 ;
        RECT 601.260 249.740 603.100 249.900 ;
        RECT 606.170 249.850 609.600 249.990 ;
        RECT 602.940 249.090 603.090 249.740 ;
        RECT 606.210 249.680 606.360 249.850 ;
        RECT 607.800 249.680 607.950 249.850 ;
        RECT 609.360 249.680 609.510 249.850 ;
        RECT 609.950 249.730 610.130 250.820 ;
        RECT 610.750 249.730 610.930 250.820 ;
        RECT 611.550 249.730 611.730 250.820 ;
        RECT 612.330 249.730 612.510 250.820 ;
        RECT 613.110 249.730 613.290 250.820 ;
        RECT 613.770 250.770 614.000 251.150 ;
        RECT 615.350 250.770 615.580 251.150 ;
        RECT 616.930 250.770 617.160 251.150 ;
        RECT 617.530 250.790 617.760 251.170 ;
        RECT 618.320 250.790 618.550 251.170 ;
        RECT 619.110 250.790 619.340 251.170 ;
        RECT 619.900 250.790 620.130 251.170 ;
        RECT 620.690 250.790 620.920 251.170 ;
        RECT 606.190 249.300 606.420 249.680 ;
        RECT 606.980 249.300 607.210 249.680 ;
        RECT 607.770 249.300 608.000 249.680 ;
        RECT 608.560 249.300 608.790 249.680 ;
        RECT 609.350 249.300 609.580 249.680 ;
        RECT 609.940 249.350 610.170 249.730 ;
        RECT 610.730 249.560 610.960 249.730 ;
        RECT 610.720 249.350 610.960 249.560 ;
        RECT 611.520 249.350 611.750 249.730 ;
        RECT 612.310 249.350 612.540 249.730 ;
        RECT 613.100 249.350 613.330 249.730 ;
        RECT 613.790 249.680 613.950 250.770 ;
        RECT 615.370 249.680 615.530 250.770 ;
        RECT 616.950 249.680 617.110 250.770 ;
        RECT 617.540 249.700 617.720 250.790 ;
        RECT 618.340 249.700 618.520 250.790 ;
        RECT 619.140 249.700 619.320 250.790 ;
        RECT 619.920 249.700 620.100 250.790 ;
        RECT 620.700 249.700 620.880 250.790 ;
        RECT 621.450 249.990 621.660 254.230 ;
        RECT 621.830 254.150 622.520 254.230 ;
        RECT 622.880 250.770 623.110 255.480 ;
        RECT 626.110 255.390 629.440 255.540 ;
        RECT 629.200 253.080 629.430 255.390 ;
        RECT 638.920 255.210 639.390 255.660 ;
        RECT 645.000 255.430 645.370 255.490 ;
        RECT 852.930 255.440 853.160 256.220 ;
        RECT 856.950 256.150 857.360 256.220 ;
        RECT 638.940 255.150 639.370 255.210 ;
        RECT 644.980 255.080 645.390 255.430 ;
        RECT 645.000 255.020 645.370 255.080 ;
        RECT 631.290 253.410 631.990 254.040 ;
        RECT 633.530 253.960 634.360 254.700 ;
        RECT 641.390 254.620 641.890 255.000 ;
        RECT 852.680 254.630 853.510 255.440 ;
        RECT 860.190 254.720 860.450 256.660 ;
        RECT 860.190 254.640 862.900 254.720 ;
        RECT 860.190 254.510 863.120 254.640 ;
        RECT 854.570 254.250 855.480 254.480 ;
        RECT 862.660 254.280 863.120 254.510 ;
        RECT 853.590 254.220 855.480 254.250 ;
        RECT 728.180 254.000 855.480 254.220 ;
        RECT 628.830 252.730 629.430 253.080 ;
        RECT 629.200 252.350 629.430 252.730 ;
        RECT 638.830 252.560 639.530 252.920 ;
        RECT 627.290 252.190 630.670 252.350 ;
        RECT 627.300 252.020 627.470 252.190 ;
        RECT 628.870 252.020 629.040 252.190 ;
        RECT 629.200 252.180 629.430 252.190 ;
        RECT 630.470 252.020 630.640 252.190 ;
        RECT 627.270 251.640 627.500 252.020 ;
        RECT 628.060 251.640 628.290 252.020 ;
        RECT 628.850 251.640 629.080 252.020 ;
        RECT 629.640 251.640 629.870 252.020 ;
        RECT 630.430 251.640 630.660 252.020 ;
        RECT 622.680 250.220 623.370 250.770 ;
        RECT 627.300 250.550 627.480 251.640 ;
        RECT 628.080 250.550 628.260 251.640 ;
        RECT 628.870 250.550 629.050 251.640 ;
        RECT 629.650 250.550 629.830 251.640 ;
        RECT 630.440 250.550 630.620 251.640 ;
        RECT 627.270 250.170 627.500 250.550 ;
        RECT 628.060 250.170 628.290 250.550 ;
        RECT 628.850 250.170 629.080 250.550 ;
        RECT 629.640 250.170 629.870 250.550 ;
        RECT 630.430 250.170 630.660 250.550 ;
        RECT 639.090 250.260 639.270 252.560 ;
        RECT 642.930 252.440 643.500 253.120 ;
        RECT 683.760 253.060 684.140 253.110 ;
        RECT 685.410 253.060 685.920 253.290 ;
        RECT 689.070 253.060 689.450 253.120 ;
        RECT 680.960 252.680 681.560 252.700 ;
        RECT 683.130 252.680 683.560 252.950 ;
        RECT 683.760 252.920 689.450 253.060 ;
        RECT 683.760 252.800 684.140 252.920 ;
        RECT 679.120 252.540 683.560 252.680 ;
        RECT 685.410 252.600 685.920 252.920 ;
        RECT 689.070 252.810 689.450 252.920 ;
        RECT 686.500 252.630 687.090 252.730 ;
        RECT 690.480 252.630 690.720 252.850 ;
        RECT 639.410 250.660 639.860 251.350 ;
        RECT 643.160 250.310 643.300 252.440 ;
        RECT 680.960 252.310 681.560 252.540 ;
        RECT 683.130 252.450 683.560 252.540 ;
        RECT 686.360 252.500 690.720 252.630 ;
        RECT 690.980 252.730 691.360 252.790 ;
        RECT 693.240 252.740 694.100 253.140 ;
        RECT 700.990 253.080 701.370 253.130 ;
        RECT 702.640 253.080 703.150 253.310 ;
        RECT 718.560 253.180 718.940 253.230 ;
        RECT 720.210 253.180 720.720 253.410 ;
        RECT 723.870 253.180 724.250 253.240 ;
        RECT 706.300 253.080 706.680 253.140 ;
        RECT 693.100 252.730 694.100 252.740 ;
        RECT 690.980 252.580 694.100 252.730 ;
        RECT 698.190 252.700 698.790 252.720 ;
        RECT 700.350 252.700 700.820 253.020 ;
        RECT 700.990 252.940 706.680 253.080 ;
        RECT 718.560 253.040 724.250 253.180 ;
        RECT 700.990 252.820 701.370 252.940 ;
        RECT 690.980 252.500 691.360 252.580 ;
        RECT 693.100 252.570 694.100 252.580 ;
        RECT 686.360 252.440 690.690 252.500 ;
        RECT 686.500 251.910 687.090 252.440 ;
        RECT 693.240 252.120 694.100 252.570 ;
        RECT 696.350 252.560 700.820 252.700 ;
        RECT 702.640 252.620 703.150 252.940 ;
        RECT 706.300 252.830 706.680 252.940 ;
        RECT 703.730 252.650 704.320 252.750 ;
        RECT 707.710 252.650 707.950 252.870 ;
        RECT 698.190 252.330 698.790 252.560 ;
        RECT 700.350 252.470 700.820 252.560 ;
        RECT 703.590 252.520 707.950 252.650 ;
        RECT 708.210 252.750 708.590 252.810 ;
        RECT 710.280 252.750 711.240 252.900 ;
        RECT 715.760 252.800 716.360 252.820 ;
        RECT 717.970 252.800 718.410 253.020 ;
        RECT 718.560 252.920 718.940 253.040 ;
        RECT 708.210 252.600 711.240 252.750 ;
        RECT 713.920 252.660 718.410 252.800 ;
        RECT 720.210 252.720 720.720 253.040 ;
        RECT 723.870 252.930 724.250 253.040 ;
        RECT 721.300 252.750 721.890 252.850 ;
        RECT 725.280 252.750 725.520 252.970 ;
        RECT 708.210 252.520 708.590 252.600 ;
        RECT 703.590 252.460 707.920 252.520 ;
        RECT 703.730 251.930 704.320 252.460 ;
        RECT 710.280 252.170 711.240 252.600 ;
        RECT 715.760 252.430 716.360 252.660 ;
        RECT 717.970 252.640 718.410 252.660 ;
        RECT 717.990 252.620 718.250 252.640 ;
        RECT 721.160 252.620 725.520 252.750 ;
        RECT 725.780 252.850 726.160 252.910 ;
        RECT 728.190 252.870 728.420 254.000 ;
        RECT 853.590 253.960 855.480 254.000 ;
        RECT 854.570 253.790 855.480 253.960 ;
        RECT 735.730 253.210 736.110 253.260 ;
        RECT 737.380 253.210 737.890 253.440 ;
        RECT 753.540 253.270 753.920 253.320 ;
        RECT 755.190 253.270 755.700 253.500 ;
        RECT 758.850 253.270 759.230 253.330 ;
        RECT 741.040 253.210 741.420 253.270 ;
        RECT 735.730 253.070 741.420 253.210 ;
        RECT 753.540 253.130 759.230 253.270 ;
        RECT 735.160 253.010 735.420 253.020 ;
        RECT 727.790 252.850 728.420 252.870 ;
        RECT 725.780 252.700 728.420 252.850 ;
        RECT 732.930 252.830 733.530 252.850 ;
        RECT 735.100 252.830 735.530 253.010 ;
        RECT 735.730 252.950 736.110 253.070 ;
        RECT 725.780 252.620 726.160 252.700 ;
        RECT 727.790 252.690 728.420 252.700 ;
        RECT 731.090 252.690 735.530 252.830 ;
        RECT 737.380 252.750 737.890 253.070 ;
        RECT 741.040 252.960 741.420 253.070 ;
        RECT 738.470 252.780 739.060 252.880 ;
        RECT 742.450 252.780 742.690 253.000 ;
        RECT 728.190 252.680 728.420 252.690 ;
        RECT 721.160 252.560 725.490 252.620 ;
        RECT 721.300 252.030 721.890 252.560 ;
        RECT 732.930 252.460 733.530 252.690 ;
        RECT 735.100 252.670 735.530 252.690 ;
        RECT 735.160 252.650 735.420 252.670 ;
        RECT 738.330 252.650 742.690 252.780 ;
        RECT 742.950 252.880 743.330 252.940 ;
        RECT 745.270 252.900 745.960 253.070 ;
        RECT 752.970 253.050 753.230 253.080 ;
        RECT 745.090 252.880 745.960 252.900 ;
        RECT 750.740 252.890 751.340 252.910 ;
        RECT 752.900 252.890 753.380 253.050 ;
        RECT 753.540 253.010 753.920 253.130 ;
        RECT 742.950 252.730 745.960 252.880 ;
        RECT 748.900 252.750 753.380 252.890 ;
        RECT 755.190 252.810 755.700 253.130 ;
        RECT 758.850 253.020 759.230 253.130 ;
        RECT 760.760 252.940 761.140 253.000 ;
        RECT 762.920 252.940 763.420 252.950 ;
        RECT 760.760 252.900 763.420 252.940 ;
        RECT 760.760 252.860 854.100 252.900 ;
        RECT 866.280 252.890 867.340 253.740 ;
        RECT 742.950 252.650 743.330 252.730 ;
        RECT 738.330 252.590 742.660 252.650 ;
        RECT 738.470 252.060 739.060 252.590 ;
        RECT 745.270 252.490 745.960 252.730 ;
        RECT 750.740 252.520 751.340 252.750 ;
        RECT 752.900 252.730 753.380 252.750 ;
        RECT 760.760 252.790 854.290 252.860 ;
        RECT 752.970 252.710 753.230 252.730 ;
        RECT 760.760 252.710 761.140 252.790 ;
        RECT 763.300 252.600 854.290 252.790 ;
        RECT 643.470 251.200 643.890 251.400 ;
        RECT 644.900 251.200 645.880 251.510 ;
        RECT 643.470 250.990 645.880 251.200 ;
        RECT 643.470 250.720 643.890 250.990 ;
        RECT 644.900 250.730 645.880 250.990 ;
        RECT 628.080 250.030 628.260 250.170 ;
        RECT 629.670 250.030 629.850 250.170 ;
        RECT 639.090 250.150 639.350 250.260 ;
        RECT 624.450 249.990 624.600 250.000 ;
        RECT 621.260 249.850 624.690 249.990 ;
        RECT 628.040 249.870 629.880 250.030 ;
        RECT 639.120 249.880 639.350 250.150 ;
        RECT 643.160 250.140 643.400 250.310 ;
        RECT 643.170 249.930 643.400 250.140 ;
        RECT 607.020 249.150 607.170 249.300 ;
        RECT 608.600 249.150 608.750 249.300 ;
        RECT 609.980 249.150 610.160 249.350 ;
        RECT 602.860 248.650 603.310 249.090 ;
        RECT 606.970 249.000 610.160 249.150 ;
        RECT 610.720 249.190 610.890 249.350 ;
        RECT 612.320 249.190 612.490 249.350 ;
        RECT 613.770 249.300 614.000 249.680 ;
        RECT 615.350 249.300 615.580 249.680 ;
        RECT 616.930 249.300 617.160 249.680 ;
        RECT 617.530 249.320 617.760 249.700 ;
        RECT 618.320 249.530 618.550 249.700 ;
        RECT 618.310 249.320 618.550 249.530 ;
        RECT 619.110 249.320 619.340 249.700 ;
        RECT 619.900 249.320 620.130 249.700 ;
        RECT 620.690 249.520 620.920 249.700 ;
        RECT 621.300 249.680 621.450 249.850 ;
        RECT 622.890 249.680 623.040 249.850 ;
        RECT 624.450 249.680 624.600 249.850 ;
        RECT 620.690 249.320 620.930 249.520 ;
        RECT 613.770 249.190 613.970 249.300 ;
        RECT 610.720 249.080 613.970 249.190 ;
        RECT 608.740 248.970 610.160 249.000 ;
        RECT 610.660 249.050 613.970 249.080 ;
        RECT 610.660 249.040 612.560 249.050 ;
        RECT 610.660 248.740 611.070 249.040 ;
        RECT 613.770 248.680 613.970 249.050 ;
        RECT 616.940 249.150 617.160 249.300 ;
        RECT 618.310 249.160 618.480 249.320 ;
        RECT 619.910 249.160 620.080 249.320 ;
        RECT 618.310 249.150 620.150 249.160 ;
        RECT 616.940 249.070 620.150 249.150 ;
        RECT 620.730 249.110 620.930 249.320 ;
        RECT 621.280 249.300 621.510 249.680 ;
        RECT 622.070 249.300 622.300 249.680 ;
        RECT 622.860 249.300 623.090 249.680 ;
        RECT 623.650 249.300 623.880 249.680 ;
        RECT 624.440 249.300 624.670 249.680 ;
        RECT 622.110 249.150 622.260 249.300 ;
        RECT 623.690 249.150 623.840 249.300 ;
        RECT 622.060 249.110 623.880 249.150 ;
        RECT 616.940 249.010 620.190 249.070 ;
        RECT 616.940 248.980 618.700 249.010 ;
        RECT 619.790 248.710 620.190 249.010 ;
        RECT 620.730 249.000 623.880 249.110 ;
        RECT 620.730 248.950 622.220 249.000 ;
        RECT 628.780 248.520 628.990 249.870 ;
        RECT 853.990 248.890 854.290 252.600 ;
        RECT 857.020 250.940 857.410 251.000 ;
        RECT 857.000 250.530 857.430 250.940 ;
        RECT 857.020 250.470 857.410 250.530 ;
        RECT 856.870 248.890 857.560 249.130 ;
        RECT 853.990 248.660 857.560 248.890 ;
        RECT 856.870 248.550 857.560 248.660 ;
        RECT 628.610 248.170 629.230 248.520 ;
        RECT 717.680 248.230 717.940 248.320 ;
        RECT 724.370 248.230 725.620 248.290 ;
        RECT 682.880 248.110 683.140 248.200 ;
        RECT 689.570 248.110 690.820 248.170 ;
        RECT 682.880 247.890 690.820 248.110 ;
        RECT 682.880 247.750 683.140 247.890 ;
        RECT 689.570 247.880 690.820 247.890 ;
        RECT 700.110 248.130 700.370 248.220 ;
        RECT 706.800 248.130 708.050 248.190 ;
        RECT 700.110 247.910 708.050 248.130 ;
        RECT 717.680 248.010 725.620 248.230 ;
        RECT 688.550 247.290 688.870 247.440 ;
        RECT 685.750 247.180 686.040 247.220 ;
        RECT 680.910 246.450 681.370 246.960 ;
        RECT 685.700 246.700 686.130 247.180 ;
        RECT 688.550 247.150 689.750 247.290 ;
        RECT 690.640 247.210 690.810 247.880 ;
        RECT 700.110 247.770 700.370 247.910 ;
        RECT 706.800 247.900 708.050 247.910 ;
        RECT 694.020 247.320 695.500 247.350 ;
        RECT 686.630 246.900 687.050 246.960 ;
        RECT 688.550 246.930 688.870 247.150 ;
        RECT 686.610 246.320 687.070 246.900 ;
        RECT 689.590 246.710 689.740 247.150 ;
        RECT 690.640 247.130 692.590 247.210 ;
        RECT 690.640 247.030 692.800 247.130 ;
        RECT 691.450 246.710 691.860 246.860 ;
        RECT 692.390 246.800 692.800 247.030 ;
        RECT 693.890 247.070 695.500 247.320 ;
        RECT 705.780 247.310 706.100 247.460 ;
        RECT 702.980 247.200 703.270 247.240 ;
        RECT 693.890 246.940 694.140 247.070 ;
        RECT 689.590 246.530 691.860 246.710 ;
        RECT 689.590 246.510 691.700 246.530 ;
        RECT 698.140 246.470 698.600 246.980 ;
        RECT 702.930 246.720 703.360 247.200 ;
        RECT 705.780 247.170 706.980 247.310 ;
        RECT 707.870 247.230 708.040 247.900 ;
        RECT 711.020 247.370 711.480 248.010 ;
        RECT 717.680 247.870 717.940 248.010 ;
        RECT 724.370 248.000 725.620 248.010 ;
        RECT 734.850 248.260 735.110 248.350 ;
        RECT 752.660 248.320 752.920 248.410 ;
        RECT 759.350 248.320 760.600 248.380 ;
        RECT 741.540 248.260 742.790 248.320 ;
        RECT 734.850 248.040 742.790 248.260 ;
        RECT 723.350 247.410 723.670 247.560 ;
        RECT 703.860 246.920 704.280 246.980 ;
        RECT 705.780 246.950 706.100 247.170 ;
        RECT 703.840 246.340 704.300 246.920 ;
        RECT 706.820 246.730 706.970 247.170 ;
        RECT 707.870 247.150 709.820 247.230 ;
        RECT 711.020 247.210 712.730 247.370 ;
        RECT 720.550 247.300 720.840 247.340 ;
        RECT 707.870 247.050 710.030 247.150 ;
        RECT 708.680 246.730 709.090 246.880 ;
        RECT 709.620 246.820 710.030 247.050 ;
        RECT 711.120 247.090 712.730 247.210 ;
        RECT 711.120 246.960 711.370 247.090 ;
        RECT 706.820 246.550 709.090 246.730 ;
        RECT 715.710 246.570 716.170 247.080 ;
        RECT 720.500 246.820 720.930 247.300 ;
        RECT 723.350 247.270 724.550 247.410 ;
        RECT 725.440 247.330 725.610 248.000 ;
        RECT 734.850 247.900 735.110 248.040 ;
        RECT 741.540 248.030 742.790 248.040 ;
        RECT 728.820 247.440 730.300 247.470 ;
        RECT 721.430 247.020 721.850 247.080 ;
        RECT 723.350 247.050 723.670 247.270 ;
        RECT 706.820 246.530 708.930 246.550 ;
        RECT 721.410 246.440 721.870 247.020 ;
        RECT 724.390 246.830 724.540 247.270 ;
        RECT 725.440 247.250 727.390 247.330 ;
        RECT 728.690 247.250 730.300 247.440 ;
        RECT 740.520 247.440 740.840 247.590 ;
        RECT 737.720 247.330 738.010 247.370 ;
        RECT 725.440 247.150 727.600 247.250 ;
        RECT 726.250 246.830 726.660 246.980 ;
        RECT 727.190 246.920 727.600 247.150 ;
        RECT 728.570 247.190 730.300 247.250 ;
        RECT 724.390 246.650 726.660 246.830 ;
        RECT 724.390 246.630 726.500 246.650 ;
        RECT 721.430 246.380 721.850 246.440 ;
        RECT 728.570 246.390 729.100 247.190 ;
        RECT 732.880 246.600 733.340 247.110 ;
        RECT 737.670 246.850 738.100 247.330 ;
        RECT 740.520 247.300 741.720 247.440 ;
        RECT 742.610 247.360 742.780 248.030 ;
        RECT 745.790 247.500 746.200 248.250 ;
        RECT 752.660 248.100 760.600 248.320 ;
        RECT 752.660 247.960 752.920 248.100 ;
        RECT 759.350 248.090 760.600 248.100 ;
        RECT 758.330 247.500 758.650 247.650 ;
        RECT 738.600 247.050 739.020 247.110 ;
        RECT 740.520 247.080 740.840 247.300 ;
        RECT 738.580 246.470 739.040 247.050 ;
        RECT 741.560 246.860 741.710 247.300 ;
        RECT 742.610 247.280 744.560 247.360 ;
        RECT 745.790 247.350 747.470 247.500 ;
        RECT 755.530 247.390 755.820 247.430 ;
        RECT 742.610 247.180 744.770 247.280 ;
        RECT 743.420 246.860 743.830 247.010 ;
        RECT 744.360 246.950 744.770 247.180 ;
        RECT 745.860 247.220 747.470 247.350 ;
        RECT 745.860 247.090 746.110 247.220 ;
        RECT 741.560 246.680 743.830 246.860 ;
        RECT 741.560 246.660 743.670 246.680 ;
        RECT 750.690 246.660 751.150 247.170 ;
        RECT 755.480 246.910 755.910 247.390 ;
        RECT 758.330 247.360 759.530 247.500 ;
        RECT 760.420 247.420 760.590 248.090 ;
        RECT 763.800 247.530 765.280 247.560 ;
        RECT 758.330 247.140 758.650 247.360 ;
        RECT 759.370 246.920 759.520 247.360 ;
        RECT 760.420 247.340 762.370 247.420 ;
        RECT 763.670 247.410 765.280 247.530 ;
        RECT 760.420 247.240 762.580 247.340 ;
        RECT 761.230 246.920 761.640 247.070 ;
        RECT 762.170 247.010 762.580 247.240 ;
        RECT 763.600 247.280 765.280 247.410 ;
        RECT 759.370 246.740 761.640 246.920 ;
        RECT 763.600 246.750 764.050 247.280 ;
        RECT 759.370 246.720 761.480 246.740 ;
        RECT 738.600 246.410 739.020 246.470 ;
        RECT 686.630 246.260 687.050 246.320 ;
        RECT 703.860 246.280 704.280 246.340 ;
        RECT 378.570 236.540 381.890 238.950 ;
        RECT 365.250 233.360 368.420 234.410 ;
        RECT 386.320 233.360 388.100 240.010 ;
        RECT 365.250 233.180 388.100 233.360 ;
        RECT 402.990 233.180 404.770 233.360 ;
        RECT 365.250 231.020 404.770 233.180 ;
        RECT 365.250 230.100 368.420 231.020 ;
        RECT 338.660 218.070 340.190 218.140 ;
        RECT 338.660 216.980 341.140 218.070 ;
        RECT 331.480 214.630 331.710 215.610 ;
        RECT 338.060 214.630 338.290 215.610 ;
        RECT 344.640 214.630 344.870 215.610 ;
        RECT 395.800 215.520 399.400 217.890 ;
        RECT 397.120 215.500 398.640 215.520 ;
        RECT 397.120 215.420 398.040 215.500 ;
        RECT 331.480 211.160 331.710 212.140 ;
        RECT 338.060 211.160 338.290 212.140 ;
        RECT 344.640 211.160 344.870 212.140 ;
        RECT 331.480 207.690 331.710 208.670 ;
        RECT 338.060 207.690 338.290 208.670 ;
        RECT 344.640 207.690 344.870 208.670 ;
        RECT 397.120 207.110 397.690 215.420 ;
        RECT 402.990 207.880 404.770 231.020 ;
        RECT 397.110 205.980 400.940 207.110 ;
        RECT 331.480 204.220 331.710 205.200 ;
        RECT 338.060 204.220 338.290 205.200 ;
        RECT 344.640 204.220 344.870 205.200 ;
        RECT 331.480 200.750 331.710 201.730 ;
        RECT 338.060 200.750 338.290 201.730 ;
        RECT 344.640 200.750 344.870 201.730 ;
        RECT 400.530 197.370 400.940 205.980 ;
        RECT 402.990 197.910 404.760 207.880 ;
        RECT 400.530 197.350 402.650 197.370 ;
        RECT 402.990 197.350 405.700 197.910 ;
        RECT 400.530 197.050 402.670 197.350 ;
        RECT 402.200 195.500 402.670 197.050 ;
        RECT 404.230 196.950 405.700 197.350 ;
        RECT 402.200 195.250 402.680 195.500 ;
        RECT 402.450 194.520 402.680 195.250 ;
        RECT 409.030 194.520 409.260 195.500 ;
        RECT 415.610 194.520 415.840 195.500 ;
        RECT 402.450 191.050 402.680 192.030 ;
        RECT 409.030 191.050 409.260 192.030 ;
        RECT 415.610 191.050 415.840 192.030 ;
        RECT 402.450 187.580 402.680 188.560 ;
        RECT 409.030 187.580 409.260 188.560 ;
        RECT 415.610 187.580 415.840 188.560 ;
        RECT 402.450 184.110 402.680 185.090 ;
        RECT 409.030 184.110 409.260 185.090 ;
        RECT 415.610 184.110 415.840 185.090 ;
        RECT 402.450 180.640 402.680 181.620 ;
        RECT 409.030 180.640 409.260 181.620 ;
        RECT 415.610 180.640 415.840 181.620 ;
        RECT 402.450 177.170 402.680 178.150 ;
        RECT 409.030 177.170 409.260 178.150 ;
        RECT 415.610 177.170 415.840 178.150 ;
      LAYER via ;
        RECT 839.055 353.265 839.315 353.525 ;
        RECT 653.030 352.470 653.290 352.730 ;
        RECT 653.030 352.150 653.290 352.410 ;
        RECT 672.050 352.525 672.310 352.785 ;
        RECT 690.115 352.455 690.375 352.715 ;
        RECT 707.700 352.600 707.960 352.860 ;
        RECT 725.550 352.505 725.810 352.765 ;
        RECT 743.820 352.560 744.080 352.820 ;
        RECT 761.590 352.550 761.850 352.810 ;
        RECT 779.595 352.485 779.855 352.745 ;
        RECT 797.760 352.545 798.020 352.805 ;
        RECT 816.140 352.570 816.400 352.830 ;
        RECT 829.015 351.715 829.275 351.975 ;
        RECT 656.085 349.620 656.665 350.200 ;
        RECT 832.190 348.140 834.050 349.360 ;
        RECT 837.430 347.235 838.970 348.455 ;
        RECT 845.810 347.095 847.030 348.315 ;
        RECT 780.270 343.450 780.850 344.670 ;
        RECT 824.880 343.620 825.140 343.880 ;
        RECT 831.355 337.030 834.815 338.890 ;
        RECT 855.765 338.775 856.345 339.355 ;
        RECT 851.400 337.810 851.660 338.070 ;
        RECT 851.400 337.490 851.660 337.750 ;
        RECT 632.280 333.685 633.180 334.265 ;
        RECT 194.365 325.630 199.745 329.410 ;
        RECT 608.755 329.205 609.015 329.465 ;
        RECT 597.175 327.995 597.755 328.575 ;
        RECT 594.385 326.425 594.645 326.685 ;
        RECT 594.705 326.425 594.965 326.685 ;
        RECT 608.755 328.885 609.015 329.145 ;
        RECT 607.365 328.030 607.945 328.610 ;
        RECT 604.120 326.430 604.380 326.690 ;
        RECT 604.440 326.430 604.700 326.690 ;
        RECT 608.720 327.820 608.980 328.080 ;
        RECT 609.695 326.375 609.955 326.635 ;
        RECT 621.335 327.805 621.595 328.065 ;
        RECT 623.215 329.120 623.475 329.380 ;
        RECT 623.535 329.120 623.795 329.380 ;
        RECT 622.315 327.800 622.575 328.060 ;
        RECT 622.635 327.800 622.895 328.060 ;
        RECT 621.300 326.310 621.560 326.570 ;
        RECT 639.455 328.855 639.715 329.115 ;
        RECT 645.485 328.675 645.745 328.935 ;
        RECT 641.940 328.230 642.200 328.490 ;
        RECT 634.085 327.590 634.665 328.170 ;
        RECT 657.790 327.675 658.050 327.935 ;
        RECT 631.735 327.130 631.995 327.390 ;
        RECT 632.055 327.130 632.315 327.390 ;
        RECT 629.410 326.325 629.670 326.585 ;
        RECT 639.320 326.160 639.580 326.420 ;
        RECT 639.640 326.160 639.900 326.420 ;
        RECT 643.515 326.360 643.775 326.620 ;
        RECT 643.515 326.040 643.775 326.300 ;
        RECT 645.530 324.380 646.110 324.960 ;
        RECT 657.645 323.625 658.225 324.205 ;
        RECT 663.370 329.790 663.630 330.050 ;
        RECT 668.920 329.795 669.180 330.055 ;
        RECT 664.325 329.480 664.585 329.740 ;
        RECT 669.940 329.535 670.200 329.795 ;
        RECT 682.265 329.615 682.525 329.875 ;
        RECT 683.210 329.415 683.470 329.675 ;
        RECT 663.420 327.105 663.680 327.365 ;
        RECT 664.470 326.850 664.730 327.110 ;
        RECT 662.460 323.645 663.040 324.225 ;
        RECT 665.615 323.780 665.875 324.040 ;
        RECT 603.385 322.290 603.645 322.550 ;
        RECT 611.165 322.330 611.425 322.590 ;
        RECT 620.290 322.310 620.550 322.570 ;
        RECT 602.330 321.920 602.590 322.180 ;
        RECT 602.650 321.920 602.910 322.180 ;
        RECT 629.220 321.765 629.480 322.025 ;
        RECT 591.365 320.015 592.585 321.235 ;
        RECT 665.615 323.460 665.875 323.720 ;
        RECT 667.195 323.855 667.455 324.115 ;
        RECT 667.515 323.855 667.775 324.115 ;
        RECT 669.305 323.515 669.565 323.775 ;
        RECT 669.990 323.630 670.570 324.210 ;
        RECT 671.805 323.710 672.065 323.970 ;
        RECT 673.815 323.405 674.075 323.665 ;
        RECT 682.195 323.800 682.455 324.060 ;
        RECT 682.195 323.480 682.455 323.740 ;
        RECT 664.805 318.805 665.065 319.065 ;
        RECT 678.185 323.095 678.445 323.355 ;
        RECT 683.145 323.330 683.405 323.590 ;
        RECT 671.415 318.180 671.675 318.440 ;
        RECT 668.320 317.620 668.580 317.880 ;
        RECT 673.780 317.665 674.040 317.925 ;
        RECT 662.945 317.200 663.205 317.460 ;
        RECT 684.440 317.270 684.700 317.530 ;
        RECT 692.385 317.445 692.965 318.025 ;
        RECT 632.675 315.580 633.255 316.160 ;
        RECT 869.805 333.170 870.385 333.750 ;
        RECT 862.030 326.680 862.290 326.940 ;
        RECT 864.460 326.405 865.040 327.305 ;
        RECT 885.530 322.860 888.670 324.400 ;
        RECT 872.910 321.625 873.170 321.885 ;
        RECT 608.605 311.035 608.865 311.295 ;
        RECT 597.025 309.825 597.605 310.405 ;
        RECT 594.235 308.255 594.495 308.515 ;
        RECT 594.555 308.255 594.815 308.515 ;
        RECT 608.605 310.715 608.865 310.975 ;
        RECT 607.215 309.860 607.795 310.440 ;
        RECT 603.970 308.260 604.230 308.520 ;
        RECT 604.290 308.260 604.550 308.520 ;
        RECT 591.650 306.125 592.550 307.025 ;
        RECT 608.570 309.650 608.830 309.910 ;
        RECT 609.545 308.205 609.805 308.465 ;
        RECT 621.185 309.635 621.445 309.895 ;
        RECT 623.065 310.950 623.325 311.210 ;
        RECT 623.385 310.950 623.645 311.210 ;
        RECT 779.355 311.485 780.575 313.345 ;
        RECT 622.165 309.630 622.425 309.890 ;
        RECT 622.485 309.630 622.745 309.890 ;
        RECT 621.150 308.140 621.410 308.400 ;
        RECT 639.305 310.685 639.565 310.945 ;
        RECT 645.335 310.505 645.595 310.765 ;
        RECT 641.790 310.060 642.050 310.320 ;
        RECT 633.935 309.420 634.515 310.000 ;
        RECT 631.785 308.725 632.365 309.305 ;
        RECT 629.260 308.155 629.520 308.415 ;
        RECT 639.170 307.990 639.430 308.250 ;
        RECT 639.490 307.990 639.750 308.250 ;
        RECT 643.365 308.190 643.625 308.450 ;
        RECT 643.365 307.870 643.625 308.130 ;
        RECT 666.275 307.945 667.495 309.165 ;
        RECT 645.380 306.210 645.960 306.790 ;
        RECT 296.255 284.350 297.475 286.210 ;
        RECT 155.010 277.150 156.230 278.690 ;
        RECT 602.305 303.855 602.565 304.115 ;
        RECT 603.235 304.120 603.495 304.380 ;
        RECT 611.015 304.160 611.275 304.420 ;
        RECT 620.140 304.140 620.400 304.400 ;
        RECT 629.070 303.595 629.330 303.855 ;
        RECT 591.690 300.715 592.590 301.615 ;
        RECT 696.500 300.915 697.400 302.135 ;
        RECT 712.505 297.435 712.765 297.695 ;
        RECT 695.020 297.090 695.280 297.350 ;
        RECT 712.505 297.115 712.765 297.375 ;
        RECT 730.095 297.405 730.355 297.665 ;
        RECT 730.095 297.085 730.355 297.345 ;
        RECT 747.810 297.510 748.070 297.770 ;
        RECT 747.810 297.190 748.070 297.450 ;
        RECT 765.540 297.440 765.800 297.700 ;
        RECT 765.540 297.120 765.800 297.380 ;
        RECT 632.580 296.275 633.480 296.855 ;
        RECT 794.595 305.035 795.815 306.255 ;
        RECT 813.180 306.055 813.440 306.315 ;
        RECT 799.915 304.965 800.175 305.225 ;
        RECT 832.815 304.970 833.075 305.230 ;
        RECT 683.505 295.795 683.765 296.055 ;
        RECT 700.995 295.840 701.255 296.100 ;
        RECT 700.910 293.825 701.490 294.405 ;
        RECT 608.555 291.855 608.815 292.115 ;
        RECT 596.975 290.645 597.555 291.225 ;
        RECT 594.185 289.075 594.445 289.335 ;
        RECT 594.505 289.075 594.765 289.335 ;
        RECT 608.555 291.535 608.815 291.795 ;
        RECT 607.165 290.680 607.745 291.260 ;
        RECT 603.920 289.080 604.180 289.340 ;
        RECT 604.240 289.080 604.500 289.340 ;
        RECT 591.385 287.180 592.605 288.400 ;
        RECT 608.520 290.470 608.780 290.730 ;
        RECT 609.495 289.025 609.755 289.285 ;
        RECT 621.135 290.455 621.395 290.715 ;
        RECT 623.015 291.770 623.275 292.030 ;
        RECT 623.335 291.770 623.595 292.030 ;
        RECT 854.170 295.325 854.430 295.585 ;
        RECT 856.945 295.165 857.205 295.425 ;
        RECT 843.890 294.200 844.150 294.460 ;
        RECT 622.115 290.450 622.375 290.710 ;
        RECT 622.435 290.450 622.695 290.710 ;
        RECT 621.100 288.960 621.360 289.220 ;
        RECT 639.255 291.505 639.515 291.765 ;
        RECT 645.285 291.325 645.545 291.585 ;
        RECT 641.740 290.880 642.000 291.140 ;
        RECT 633.885 290.240 634.465 290.820 ;
        RECT 631.410 289.835 631.670 290.095 ;
        RECT 631.730 289.835 631.990 290.095 ;
        RECT 629.210 288.975 629.470 289.235 ;
        RECT 639.120 288.810 639.380 289.070 ;
        RECT 639.440 288.810 639.700 289.070 ;
        RECT 643.315 289.010 643.575 289.270 ;
        RECT 643.315 288.690 643.575 288.950 ;
        RECT 645.330 287.030 645.910 287.610 ;
        RECT 602.120 284.650 602.380 284.910 ;
        RECT 602.440 284.650 602.700 284.910 ;
        RECT 603.185 284.940 603.445 285.200 ;
        RECT 610.965 284.980 611.225 285.240 ;
        RECT 620.090 284.960 620.350 285.220 ;
        RECT 629.020 284.415 629.280 284.675 ;
        RECT 591.325 281.640 592.545 282.860 ;
        RECT 632.655 277.720 633.235 278.620 ;
        RECT 852.715 293.090 853.615 293.670 ;
        RECT 694.855 288.610 696.075 290.470 ;
        RECT 820.070 290.535 820.330 290.795 ;
        RECT 799.710 281.050 799.970 281.310 ;
        RECT 802.055 280.605 802.955 281.505 ;
        RECT 683.305 279.230 683.565 279.490 ;
        RECT 695.070 279.305 695.650 279.885 ;
        RECT 700.765 279.400 701.025 279.660 ;
        RECT 700.765 279.080 701.025 279.340 ;
        RECT 713.430 279.300 714.010 279.880 ;
        RECT 718.360 279.145 718.620 279.405 ;
        RECT 727.235 279.240 727.815 279.820 ;
        RECT 735.605 279.190 735.865 279.450 ;
        RECT 747.505 279.260 748.085 279.840 ;
        RECT 753.070 279.160 753.330 279.420 ;
        RECT 833.380 288.705 833.640 288.965 ;
        RECT 843.920 292.560 844.180 292.820 ;
        RECT 843.920 292.240 844.180 292.500 ;
        RECT 849.165 291.865 849.745 292.445 ;
        RECT 868.235 291.845 868.495 292.105 ;
        RECT 868.555 291.845 868.815 292.105 ;
        RECT 868.875 291.845 869.135 292.105 ;
        RECT 856.985 289.695 857.245 289.955 ;
        RECT 840.535 288.205 840.795 288.465 ;
        RECT 814.465 286.255 815.045 286.835 ;
        RECT 840.485 286.515 840.745 286.775 ;
        RECT 819.095 285.510 819.355 285.770 ;
        RECT 816.360 284.680 817.260 285.260 ;
        RECT 832.995 285.345 834.215 286.245 ;
        RECT 821.790 281.085 822.050 281.345 ;
        RECT 853.025 283.565 853.285 283.825 ;
        RECT 853.025 283.245 853.285 283.505 ;
        RECT 841.130 281.235 841.390 281.495 ;
        RECT 820.870 280.585 821.130 280.845 ;
        RECT 828.135 280.370 828.395 280.630 ;
        RECT 829.090 280.340 829.350 280.600 ;
        RECT 836.695 280.610 836.955 280.870 ;
        RECT 849.750 280.670 850.010 280.930 ;
        RECT 829.090 280.020 829.350 280.280 ;
        RECT 841.105 280.305 841.365 280.565 ;
        RECT 842.010 279.960 842.270 280.220 ;
        RECT 852.005 280.240 852.585 280.820 ;
        RECT 836.550 278.310 836.810 278.570 ;
        RECT 836.870 278.310 837.130 278.570 ;
        RECT 840.690 278.330 840.950 278.590 ;
        RECT 841.010 278.330 841.270 278.590 ;
        RECT 853.160 277.705 853.420 277.965 ;
        RECT 834.615 276.155 834.875 276.415 ;
        RECT 834.935 276.155 835.195 276.415 ;
        RECT 608.475 273.385 608.735 273.645 ;
        RECT 596.895 272.175 597.475 272.755 ;
        RECT 594.105 270.605 594.365 270.865 ;
        RECT 594.425 270.605 594.685 270.865 ;
        RECT 608.475 273.065 608.735 273.325 ;
        RECT 607.085 272.210 607.665 272.790 ;
        RECT 603.840 270.610 604.100 270.870 ;
        RECT 604.160 270.610 604.420 270.870 ;
        RECT 591.325 269.050 592.545 269.950 ;
        RECT 608.440 272.000 608.700 272.260 ;
        RECT 609.415 270.555 609.675 270.815 ;
        RECT 621.055 271.985 621.315 272.245 ;
        RECT 679.940 274.510 680.200 274.770 ;
        RECT 685.555 274.505 685.815 274.765 ;
        RECT 622.935 273.300 623.195 273.560 ;
        RECT 623.255 273.300 623.515 273.560 ;
        RECT 681.150 273.905 681.410 274.165 ;
        RECT 683.235 274.100 683.495 274.360 ;
        RECT 685.555 274.185 685.815 274.445 ;
        RECT 686.685 273.880 686.945 274.140 ;
        RECT 686.685 273.560 686.945 273.820 ;
        RECT 692.870 273.830 693.450 274.410 ;
        RECT 698.380 273.925 698.640 274.185 ;
        RECT 700.475 274.145 700.735 274.405 ;
        RECT 702.785 274.525 703.045 274.785 ;
        RECT 720.355 274.625 720.615 274.885 ;
        RECT 702.785 274.205 703.045 274.465 ;
        RECT 703.915 273.900 704.175 274.160 ;
        RECT 703.915 273.580 704.175 273.840 ;
        RECT 710.070 273.640 710.970 274.540 ;
        RECT 715.950 274.025 716.210 274.285 ;
        RECT 718.080 274.230 718.340 274.490 ;
        RECT 720.355 274.305 720.615 274.565 ;
        RECT 721.485 274.000 721.745 274.260 ;
        RECT 721.485 273.680 721.745 273.940 ;
        RECT 727.740 273.980 728.320 274.560 ;
        RECT 737.525 274.655 737.785 274.915 ;
        RECT 733.120 274.055 733.380 274.315 ;
        RECT 735.205 274.240 735.465 274.500 ;
        RECT 737.525 274.335 737.785 274.595 ;
        RECT 738.655 274.030 738.915 274.290 ;
        RECT 738.655 273.710 738.915 273.970 ;
        RECT 745.005 273.870 745.905 274.770 ;
        RECT 755.335 274.715 755.595 274.975 ;
        RECT 750.930 274.115 751.190 274.375 ;
        RECT 753.030 274.290 753.290 274.550 ;
        RECT 755.335 274.395 755.595 274.655 ;
        RECT 762.655 273.970 763.555 274.870 ;
        RECT 797.680 273.745 798.260 274.325 ;
        RECT 815.945 273.905 816.525 274.485 ;
        RECT 834.705 274.185 834.965 274.445 ;
        RECT 622.035 271.980 622.295 272.240 ;
        RECT 622.355 271.980 622.615 272.240 ;
        RECT 621.020 270.490 621.280 270.750 ;
        RECT 639.175 273.035 639.435 273.295 ;
        RECT 645.205 272.855 645.465 273.115 ;
        RECT 641.660 272.410 641.920 272.670 ;
        RECT 633.805 271.770 634.385 272.350 ;
        RECT 784.405 272.295 784.665 272.555 ;
        RECT 803.310 272.335 803.570 272.595 ;
        RECT 822.150 272.340 822.410 272.600 ;
        RECT 837.105 273.775 837.365 274.035 ;
        RECT 837.105 273.455 837.365 273.715 ;
        RECT 836.825 272.740 837.085 273.000 ;
        RECT 837.145 272.740 837.405 273.000 ;
        RECT 631.630 271.280 631.890 271.540 ;
        RECT 629.130 270.505 629.390 270.765 ;
        RECT 639.040 270.340 639.300 270.600 ;
        RECT 639.360 270.340 639.620 270.600 ;
        RECT 643.235 270.540 643.495 270.800 ;
        RECT 822.175 270.575 822.435 270.835 ;
        RECT 865.310 281.230 865.890 282.130 ;
        RECT 857.060 278.945 857.320 279.205 ;
        RECT 853.120 271.665 853.380 271.925 ;
        RECT 643.235 270.220 643.495 270.480 ;
        RECT 645.250 268.560 645.830 269.140 ;
        RECT 680.105 268.310 680.365 268.570 ;
        RECT 681.030 268.105 681.290 268.365 ;
        RECT 685.805 268.340 686.065 268.600 ;
        RECT 686.730 268.170 686.990 268.430 ;
        RECT 686.730 267.850 686.990 268.110 ;
        RECT 698.260 268.125 698.520 268.385 ;
        RECT 703.035 268.360 703.295 268.620 ;
        RECT 711.140 269.170 711.400 269.430 ;
        RECT 711.140 268.850 711.400 269.110 ;
        RECT 703.960 268.190 704.220 268.450 ;
        RECT 703.960 267.870 704.220 268.130 ;
        RECT 715.830 268.225 716.090 268.485 ;
        RECT 720.605 268.460 720.865 268.720 ;
        RECT 721.530 268.290 721.790 268.550 ;
        RECT 721.530 267.970 721.790 268.230 ;
        RECT 728.725 268.380 728.985 268.640 ;
        RECT 728.725 268.060 728.985 268.320 ;
        RECT 733.000 268.255 733.260 268.515 ;
        RECT 737.775 268.490 738.035 268.750 ;
        RECT 745.885 269.520 746.145 269.780 ;
        RECT 745.885 269.200 746.145 269.460 ;
        RECT 738.700 268.320 738.960 268.580 ;
        RECT 738.700 268.000 738.960 268.260 ;
        RECT 745.885 268.880 746.145 269.140 ;
        RECT 750.810 268.315 751.070 268.575 ;
        RECT 755.585 268.550 755.845 268.810 ;
        RECT 763.715 268.640 763.975 268.900 ;
        RECT 763.715 268.320 763.975 268.580 ;
        RECT 601.520 266.190 601.780 266.450 ;
        RECT 601.840 266.190 602.100 266.450 ;
        RECT 602.160 266.190 602.420 266.450 ;
        RECT 603.105 266.470 603.365 266.730 ;
        RECT 610.885 266.510 611.145 266.770 ;
        RECT 620.010 266.490 620.270 266.750 ;
        RECT 797.685 266.620 798.265 267.200 ;
        RECT 816.265 266.520 816.845 267.100 ;
        RECT 628.940 265.945 629.200 266.205 ;
        RECT 784.430 264.815 784.690 265.075 ;
        RECT 802.955 264.850 803.215 265.110 ;
        RECT 591.195 263.675 592.415 264.575 ;
        RECT 632.510 260.220 633.410 260.800 ;
        RECT 692.555 263.650 693.775 264.550 ;
        RECT 837.005 267.480 837.265 267.740 ;
        RECT 839.535 266.755 839.795 267.015 ;
        RECT 850.995 267.045 851.575 267.625 ;
        RECT 853.225 264.920 853.485 265.180 ;
        RECT 850.885 261.600 851.785 262.180 ;
        RECT 852.575 261.810 853.155 262.390 ;
        RECT 853.505 261.305 853.765 261.565 ;
        RECT 683.285 257.700 683.545 257.960 ;
        RECT 694.495 257.815 695.075 258.395 ;
        RECT 700.745 257.870 701.005 258.130 ;
        RECT 712.830 257.990 713.090 258.250 ;
        RECT 713.150 257.990 713.410 258.250 ;
        RECT 700.745 257.550 701.005 257.810 ;
        RECT 718.340 257.615 718.600 257.875 ;
        RECT 730.025 257.815 730.605 258.395 ;
        RECT 735.585 257.660 735.845 257.920 ;
        RECT 747.615 257.815 748.195 258.395 ;
        RECT 846.745 258.290 847.325 259.190 ;
        RECT 853.495 258.855 853.755 259.115 ;
        RECT 753.050 257.630 753.310 257.890 ;
        RECT 608.325 255.655 608.585 255.915 ;
        RECT 334.240 229.925 336.100 233.385 ;
        RECT 596.745 254.445 597.325 255.025 ;
        RECT 593.955 252.875 594.215 253.135 ;
        RECT 594.275 252.875 594.535 253.135 ;
        RECT 608.325 255.335 608.585 255.595 ;
        RECT 606.935 254.480 607.515 255.060 ;
        RECT 603.690 252.880 603.950 253.140 ;
        RECT 604.010 252.880 604.270 253.140 ;
        RECT 591.265 250.270 592.165 251.490 ;
        RECT 608.290 254.270 608.550 254.530 ;
        RECT 609.265 252.825 609.525 253.085 ;
        RECT 620.905 254.255 621.165 254.515 ;
        RECT 622.785 255.570 623.045 255.830 ;
        RECT 623.105 255.570 623.365 255.830 ;
        RECT 856.075 256.730 856.335 256.990 ;
        RECT 751.670 255.730 752.250 256.310 ;
        RECT 851.030 255.910 851.610 256.490 ;
        RECT 621.885 254.250 622.145 254.510 ;
        RECT 622.205 254.250 622.465 254.510 ;
        RECT 620.870 252.760 621.130 253.020 ;
        RECT 639.025 255.305 639.285 255.565 ;
        RECT 645.055 255.125 645.315 255.385 ;
        RECT 641.510 254.680 641.770 254.940 ;
        RECT 852.805 254.745 853.385 255.325 ;
        RECT 633.655 254.040 634.235 254.620 ;
        RECT 631.515 253.610 631.775 253.870 ;
        RECT 628.980 252.775 629.240 253.035 ;
        RECT 638.890 252.610 639.150 252.870 ;
        RECT 639.210 252.610 639.470 252.870 ;
        RECT 643.085 252.810 643.345 253.070 ;
        RECT 685.535 252.975 685.795 253.235 ;
        RECT 643.085 252.490 643.345 252.750 ;
        RECT 681.130 252.375 681.390 252.635 ;
        RECT 683.215 252.570 683.475 252.830 ;
        RECT 685.535 252.655 685.795 252.915 ;
        RECT 686.665 252.350 686.925 252.610 ;
        RECT 686.665 252.030 686.925 252.290 ;
        RECT 693.380 252.180 693.960 253.080 ;
        RECT 698.360 252.395 698.620 252.655 ;
        RECT 700.455 252.615 700.715 252.875 ;
        RECT 702.765 252.995 703.025 253.255 ;
        RECT 720.335 253.095 720.595 253.355 ;
        RECT 702.765 252.675 703.025 252.935 ;
        RECT 703.895 252.370 704.155 252.630 ;
        RECT 703.895 252.050 704.155 252.310 ;
        RECT 710.470 252.245 711.050 252.825 ;
        RECT 715.930 252.495 716.190 252.755 ;
        RECT 718.060 252.700 718.320 252.960 ;
        RECT 720.335 252.775 720.595 253.035 ;
        RECT 721.465 252.470 721.725 252.730 ;
        RECT 737.505 253.125 737.765 253.385 ;
        RECT 755.315 253.185 755.575 253.445 ;
        RECT 733.100 252.525 733.360 252.785 ;
        RECT 735.185 252.710 735.445 252.970 ;
        RECT 737.505 252.805 737.765 253.065 ;
        RECT 738.635 252.500 738.895 252.760 ;
        RECT 721.465 252.150 721.725 252.410 ;
        RECT 745.325 252.490 745.905 253.070 ;
        RECT 750.910 252.585 751.170 252.845 ;
        RECT 753.010 252.760 753.270 253.020 ;
        RECT 755.315 252.865 755.575 253.125 ;
        RECT 866.360 253.025 867.260 253.605 ;
        RECT 738.635 252.180 738.895 252.440 ;
        RECT 645.100 250.830 645.680 251.410 ;
        RECT 602.955 248.740 603.215 249.000 ;
        RECT 610.735 248.780 610.995 249.040 ;
        RECT 619.860 248.760 620.120 249.020 ;
        RECT 857.085 250.605 857.345 250.865 ;
        RECT 856.925 248.550 857.505 249.130 ;
        RECT 628.790 248.215 629.050 248.475 ;
        RECT 681.010 246.575 681.270 246.835 ;
        RECT 685.785 246.810 686.045 247.070 ;
        RECT 686.710 246.640 686.970 246.900 ;
        RECT 686.710 246.320 686.970 246.580 ;
        RECT 698.240 246.595 698.500 246.855 ;
        RECT 703.015 246.830 703.275 247.090 ;
        RECT 711.120 247.640 711.380 247.900 ;
        RECT 711.120 247.320 711.380 247.580 ;
        RECT 703.940 246.660 704.200 246.920 ;
        RECT 703.940 246.340 704.200 246.600 ;
        RECT 715.810 246.695 716.070 246.955 ;
        RECT 720.585 246.930 720.845 247.190 ;
        RECT 721.510 246.760 721.770 247.020 ;
        RECT 721.510 246.440 721.770 246.700 ;
        RECT 728.705 246.850 728.965 247.110 ;
        RECT 728.705 246.530 728.965 246.790 ;
        RECT 732.980 246.725 733.240 246.985 ;
        RECT 737.755 246.960 738.015 247.220 ;
        RECT 745.865 247.990 746.125 248.250 ;
        RECT 745.865 247.670 746.125 247.930 ;
        RECT 738.680 246.790 738.940 247.050 ;
        RECT 738.680 246.470 738.940 246.730 ;
        RECT 745.865 247.350 746.125 247.610 ;
        RECT 750.790 246.785 751.050 247.045 ;
        RECT 755.565 247.020 755.825 247.280 ;
        RECT 763.695 247.110 763.955 247.370 ;
        RECT 763.695 246.790 763.955 247.050 ;
        RECT 378.660 236.655 381.800 238.835 ;
        RECT 365.425 230.205 368.245 234.305 ;
        RECT 395.870 215.615 399.330 217.795 ;
      LAYER met2 ;
        RECT 839.000 353.080 839.370 353.710 ;
        RECT 707.680 353.010 707.980 353.060 ;
        RECT 652.900 352.100 653.420 352.780 ;
        RECT 671.930 352.290 672.430 352.980 ;
        RECT 690.060 352.250 690.480 352.930 ;
        RECT 707.640 352.320 708.030 353.010 ;
        RECT 725.520 352.350 725.890 352.940 ;
        RECT 743.790 352.400 744.140 353.020 ;
        RECT 761.520 352.380 761.920 352.980 ;
        RECT 725.540 352.330 725.820 352.350 ;
        RECT 779.540 352.340 779.920 352.900 ;
        RECT 797.680 352.430 798.100 352.950 ;
        RECT 816.070 352.430 816.470 352.980 ;
        RECT 828.900 351.610 829.390 352.080 ;
        RECT 829.060 350.410 829.200 351.610 ;
        RECT 656.060 349.480 656.690 350.340 ;
        RECT 828.800 349.650 829.470 350.410 ;
        RECT 832.110 347.980 834.130 349.520 ;
        RECT 780.120 343.340 781.000 344.780 ;
        RECT 824.850 344.060 825.170 344.070 ;
        RECT 824.800 343.410 825.220 344.060 ;
        RECT 832.380 339.040 833.860 347.980 ;
        RECT 837.310 347.820 839.090 348.630 ;
        RECT 845.710 347.820 847.130 348.470 ;
        RECT 837.310 347.310 847.130 347.820 ;
        RECT 837.310 347.060 839.090 347.310 ;
        RECT 845.710 346.940 847.130 347.310 ;
        RECT 194.240 334.650 199.610 338.700 ;
        RECT 831.230 336.880 834.940 339.040 ;
        RECT 855.630 338.630 856.480 339.500 ;
        RECT 851.270 337.420 851.790 338.140 ;
        RECT 195.760 329.460 197.690 334.650 ;
        RECT 632.250 333.570 633.210 334.380 ;
        RECT 194.240 325.580 199.870 329.460 ;
        RECT 608.600 329.290 609.170 329.650 ;
        RECT 663.300 329.610 663.690 330.230 ;
        RECT 623.130 329.290 623.880 329.520 ;
        RECT 664.250 329.370 664.670 329.890 ;
        RECT 668.810 329.630 669.240 330.250 ;
        RECT 669.850 329.350 670.270 329.980 ;
        RECT 682.130 329.410 682.640 330.050 ;
        RECT 608.600 329.060 623.880 329.290 ;
        RECT 683.130 329.270 683.550 329.820 ;
        RECT 597.150 328.520 597.780 328.760 ;
        RECT 608.600 328.700 609.170 329.060 ;
        RECT 623.130 328.980 623.880 329.060 ;
        RECT 639.400 328.960 639.770 329.260 ;
        RECT 639.360 328.710 639.770 328.960 ;
        RECT 607.270 328.520 608.040 328.690 ;
        RECT 597.150 328.150 608.040 328.520 ;
        RECT 597.150 327.810 597.780 328.150 ;
        RECT 607.270 327.950 608.040 328.150 ;
        RECT 608.580 328.000 609.120 328.210 ;
        RECT 621.260 328.000 621.670 328.130 ;
        RECT 608.580 327.830 621.670 328.000 ;
        RECT 608.580 327.690 609.120 327.830 ;
        RECT 621.260 327.740 621.670 327.830 ;
        RECT 622.310 328.070 622.900 328.210 ;
        RECT 634.020 328.070 634.730 328.270 ;
        RECT 622.310 327.760 634.730 328.070 ;
        RECT 622.310 327.650 622.900 327.760 ;
        RECT 631.690 326.970 632.360 327.550 ;
        RECT 634.020 327.490 634.730 327.760 ;
        RECT 639.360 326.960 639.600 328.710 ;
        RECT 645.460 328.580 645.770 329.030 ;
        RECT 856.090 328.980 856.450 338.630 ;
        RECT 869.720 333.060 870.470 333.860 ;
        RECT 641.880 328.150 642.260 328.570 ;
        RECT 639.360 326.910 639.790 326.960 ;
        RECT 645.490 326.920 645.710 328.580 ;
        RECT 657.720 327.890 658.120 328.040 ;
        RECT 677.980 327.900 678.350 327.920 ;
        RECT 673.000 327.890 678.350 327.900 ;
        RECT 657.720 327.690 678.350 327.890 ;
        RECT 657.720 327.570 658.120 327.690 ;
        RECT 677.980 327.680 678.350 327.690 ;
        RECT 663.370 327.440 663.730 327.500 ;
        RECT 642.700 326.910 645.710 326.920 ;
        RECT 594.360 326.370 594.990 326.740 ;
        RECT 603.980 326.590 604.840 326.890 ;
        RECT 609.550 326.590 610.100 326.840 ;
        RECT 639.360 326.740 645.710 326.910 ;
        RECT 663.300 326.800 663.790 327.440 ;
        RECT 642.700 326.720 645.710 326.740 ;
        RECT 603.980 326.380 610.100 326.590 ;
        RECT 591.340 319.920 592.610 321.330 ;
        RECT 594.490 321.270 594.900 326.370 ;
        RECT 603.980 326.230 604.840 326.380 ;
        RECT 609.550 326.170 610.100 326.380 ;
        RECT 621.240 326.530 621.620 326.630 ;
        RECT 629.310 326.530 629.770 326.680 ;
        RECT 621.240 326.340 629.770 326.530 ;
        RECT 639.500 326.520 639.710 326.530 ;
        RECT 621.240 326.250 621.620 326.340 ;
        RECT 629.310 326.230 629.770 326.340 ;
        RECT 639.310 326.390 639.910 326.520 ;
        RECT 641.850 326.390 642.280 326.550 ;
        RECT 639.310 326.180 642.280 326.390 ;
        RECT 639.310 326.060 639.910 326.180 ;
        RECT 641.850 326.020 642.280 326.180 ;
        RECT 643.410 325.940 643.880 326.720 ;
        RECT 664.260 326.640 664.920 327.310 ;
        RECT 645.380 324.230 646.260 325.110 ;
        RECT 603.340 322.460 603.690 322.690 ;
        RECT 611.140 322.460 611.450 322.680 ;
        RECT 603.340 322.280 611.450 322.460 ;
        RECT 602.330 321.820 602.910 322.280 ;
        RECT 603.340 322.150 603.690 322.280 ;
        RECT 611.140 322.240 611.450 322.280 ;
        RECT 620.270 322.210 620.570 322.670 ;
        RECT 620.360 321.990 620.510 322.210 ;
        RECT 629.090 321.990 629.610 322.120 ;
        RECT 620.360 321.790 629.610 321.990 ;
        RECT 629.090 321.670 629.610 321.790 ;
        RECT 645.620 321.320 645.840 324.230 ;
        RECT 657.600 323.450 658.270 324.380 ;
        RECT 662.330 323.550 663.170 324.320 ;
        RECT 662.680 323.300 662.910 323.550 ;
        RECT 665.470 323.340 666.020 324.160 ;
        RECT 667.060 323.650 667.910 324.320 ;
        RECT 669.260 323.470 669.610 323.970 ;
        RECT 669.990 323.570 670.570 324.270 ;
        RECT 671.680 323.480 672.190 324.280 ;
        RECT 660.500 323.290 662.910 323.300 ;
        RECT 657.110 323.230 662.910 323.290 ;
        RECT 656.890 323.070 662.910 323.230 ;
        RECT 667.370 323.320 669.610 323.470 ;
        RECT 667.370 323.180 669.540 323.320 ;
        RECT 656.890 323.060 662.900 323.070 ;
        RECT 656.890 323.050 660.740 323.060 ;
        RECT 656.890 322.390 657.350 323.050 ;
        RECT 636.280 321.300 645.850 321.320 ;
        RECT 614.050 321.270 645.850 321.300 ;
        RECT 594.490 320.970 645.850 321.270 ;
        RECT 667.410 321.140 667.580 323.180 ;
        RECT 662.970 321.070 667.610 321.140 ;
        RECT 594.490 320.890 637.260 320.970 ;
        RECT 662.950 320.910 667.610 321.070 ;
        RECT 671.830 321.060 671.970 323.480 ;
        RECT 673.770 323.310 674.120 323.760 ;
        RECT 678.190 323.480 678.350 327.680 ;
        RECT 668.350 320.960 671.970 321.060 ;
        RECT 668.340 320.910 671.970 320.960 ;
        RECT 594.490 320.860 617.700 320.890 ;
        RECT 662.950 317.590 663.120 320.910 ;
        RECT 667.410 320.890 667.580 320.910 ;
        RECT 668.340 320.900 671.940 320.910 ;
        RECT 664.800 319.020 665.070 319.240 ;
        RECT 666.060 319.020 666.270 319.050 ;
        RECT 664.800 318.820 666.270 319.020 ;
        RECT 664.800 318.630 665.070 318.820 ;
        RECT 662.850 317.070 663.300 317.590 ;
        RECT 632.540 316.230 633.390 316.240 ;
        RECT 632.540 315.500 633.490 316.230 ;
        RECT 632.640 315.490 633.490 315.500 ;
        RECT 666.060 315.580 666.270 318.820 ;
        RECT 668.340 318.670 668.490 320.900 ;
        RECT 668.230 318.020 668.680 318.670 ;
        RECT 671.340 318.020 671.750 318.600 ;
        RECT 673.850 318.040 673.990 323.310 ;
        RECT 678.140 322.970 678.490 323.480 ;
        RECT 682.070 323.370 682.580 324.170 ;
        RECT 683.070 323.130 683.480 323.790 ;
        RECT 856.090 321.830 856.390 328.980 ;
        RECT 861.940 326.850 862.380 327.140 ;
        RECT 864.330 326.850 865.170 327.390 ;
        RECT 861.940 326.620 865.170 326.850 ;
        RECT 861.940 326.610 863.440 326.620 ;
        RECT 861.940 326.480 862.380 326.610 ;
        RECT 864.330 326.320 865.170 326.620 ;
        RECT 885.390 322.690 888.810 324.570 ;
        RECT 872.860 321.830 873.220 322.090 ;
        RECT 856.080 321.820 856.390 321.830 ;
        RECT 863.080 321.820 873.220 321.830 ;
        RECT 856.080 321.540 873.220 321.820 ;
        RECT 856.080 321.530 856.390 321.540 ;
        RECT 863.080 321.530 873.220 321.540 ;
        RECT 856.090 321.440 856.390 321.530 ;
        RECT 872.860 321.420 873.220 321.530 ;
        RECT 668.300 317.490 668.600 318.020 ;
        RECT 673.770 317.550 674.050 318.040 ;
        RECT 684.440 317.130 684.700 317.670 ;
        RECT 692.320 317.350 693.030 318.120 ;
        RECT 666.060 315.570 683.750 315.580 ;
        RECT 684.470 315.570 684.680 317.130 ;
        RECT 666.060 315.390 684.680 315.570 ;
        RECT 684.470 315.380 684.680 315.390 ;
        RECT 608.450 311.120 609.020 311.480 ;
        RECT 622.980 311.120 623.730 311.350 ;
        RECT 608.450 310.890 623.730 311.120 ;
        RECT 597.000 310.350 597.630 310.590 ;
        RECT 608.450 310.530 609.020 310.890 ;
        RECT 622.980 310.810 623.730 310.890 ;
        RECT 639.250 310.790 639.620 311.090 ;
        RECT 639.210 310.540 639.620 310.790 ;
        RECT 607.120 310.350 607.890 310.520 ;
        RECT 597.000 309.980 607.890 310.350 ;
        RECT 597.000 309.640 597.630 309.980 ;
        RECT 607.120 309.780 607.890 309.980 ;
        RECT 608.430 309.830 608.970 310.040 ;
        RECT 621.110 309.830 621.520 309.960 ;
        RECT 608.430 309.660 621.520 309.830 ;
        RECT 608.430 309.520 608.970 309.660 ;
        RECT 621.110 309.570 621.520 309.660 ;
        RECT 622.160 309.900 622.750 310.040 ;
        RECT 633.870 309.900 634.580 310.100 ;
        RECT 622.160 309.590 634.580 309.900 ;
        RECT 622.160 309.480 622.750 309.590 ;
        RECT 594.210 308.200 594.840 308.570 ;
        RECT 603.830 308.420 604.690 308.720 ;
        RECT 609.400 308.420 609.950 308.670 ;
        RECT 631.720 308.660 632.430 309.370 ;
        RECT 633.870 309.320 634.580 309.590 ;
        RECT 639.210 308.790 639.450 310.540 ;
        RECT 645.310 310.410 645.620 310.860 ;
        RECT 641.730 309.980 642.110 310.400 ;
        RECT 639.210 308.740 639.640 308.790 ;
        RECT 645.340 308.750 645.560 310.410 ;
        RECT 642.550 308.740 645.560 308.750 ;
        RECT 639.210 308.570 645.560 308.740 ;
        RECT 642.550 308.550 645.560 308.570 ;
        RECT 603.830 308.210 609.950 308.420 ;
        RECT 591.550 305.940 592.650 307.210 ;
        RECT 594.340 303.100 594.750 308.200 ;
        RECT 603.830 308.060 604.690 308.210 ;
        RECT 609.400 308.000 609.950 308.210 ;
        RECT 621.090 308.360 621.470 308.460 ;
        RECT 629.160 308.360 629.620 308.510 ;
        RECT 621.090 308.170 629.620 308.360 ;
        RECT 639.350 308.350 639.560 308.360 ;
        RECT 621.090 308.080 621.470 308.170 ;
        RECT 629.160 308.060 629.620 308.170 ;
        RECT 639.160 308.220 639.760 308.350 ;
        RECT 641.700 308.220 642.130 308.380 ;
        RECT 639.160 308.010 642.130 308.220 ;
        RECT 639.160 307.890 639.760 308.010 ;
        RECT 641.700 307.850 642.130 308.010 ;
        RECT 643.260 307.770 643.730 308.550 ;
        RECT 666.230 307.780 667.540 309.330 ;
        RECT 645.230 306.060 646.110 306.940 ;
        RECT 603.190 304.290 603.540 304.520 ;
        RECT 610.990 304.290 611.300 304.510 ;
        RECT 602.140 303.730 602.740 304.250 ;
        RECT 603.190 304.110 611.300 304.290 ;
        RECT 603.190 303.980 603.540 304.110 ;
        RECT 610.990 304.070 611.300 304.110 ;
        RECT 620.120 304.040 620.420 304.500 ;
        RECT 620.210 303.820 620.360 304.040 ;
        RECT 628.940 303.820 629.460 303.950 ;
        RECT 620.210 303.620 629.460 303.820 ;
        RECT 628.940 303.500 629.460 303.620 ;
        RECT 645.470 303.150 645.690 306.060 ;
        RECT 692.340 303.360 692.830 317.350 ;
        RECT 779.340 312.570 780.590 313.440 ;
        RECT 813.190 312.570 813.470 312.600 ;
        RECT 779.340 312.140 813.470 312.570 ;
        RECT 779.340 311.390 780.590 312.140 ;
        RECT 813.190 306.430 813.470 312.140 ;
        RECT 794.470 304.980 795.940 306.310 ;
        RECT 813.120 305.940 813.500 306.430 ;
        RECT 799.900 304.840 800.190 305.350 ;
        RECT 692.340 303.340 700.440 303.360 ;
        RECT 700.980 303.340 701.270 303.390 ;
        RECT 636.130 303.130 645.700 303.150 ;
        RECT 613.900 303.100 645.700 303.130 ;
        RECT 594.340 302.800 645.700 303.100 ;
        RECT 692.340 302.930 701.270 303.340 ;
        RECT 799.930 303.150 800.170 304.840 ;
        RECT 832.740 304.770 833.150 305.430 ;
        RECT 832.940 303.150 833.150 304.770 ;
        RECT 799.930 302.970 833.170 303.150 ;
        RECT 832.940 302.960 833.150 302.970 ;
        RECT 594.340 302.720 637.110 302.800 ;
        RECT 594.340 302.690 617.550 302.720 ;
        RECT 591.590 300.530 592.690 301.800 ;
        RECT 696.400 301.340 697.500 302.260 ;
        RECT 683.570 301.020 697.500 301.340 ;
        RECT 632.560 296.160 633.500 296.970 ;
        RECT 683.570 296.110 683.750 301.020 ;
        RECT 696.400 300.790 697.500 301.020 ;
        RECT 694.940 296.930 695.340 297.510 ;
        RECT 700.980 296.180 701.270 302.930 ;
        RECT 712.470 296.970 712.800 297.840 ;
        RECT 730.080 296.950 730.370 297.800 ;
        RECT 747.750 297.000 748.140 297.980 ;
        RECT 765.510 297.450 765.830 297.760 ;
        RECT 765.510 297.060 765.880 297.450 ;
        RECT 683.470 295.740 683.800 296.110 ;
        RECT 700.950 295.760 701.300 296.180 ;
        RECT 683.520 294.390 683.740 295.740 ;
        RECT 701.030 294.510 701.200 295.760 ;
        RECT 700.820 293.720 701.580 294.510 ;
        RECT 729.960 292.450 731.040 292.650 ;
        RECT 608.400 291.940 608.970 292.300 ;
        RECT 622.930 291.940 623.680 292.170 ;
        RECT 728.470 292.100 731.040 292.450 ;
        RECT 608.400 291.710 623.680 291.940 ;
        RECT 728.430 291.950 731.040 292.100 ;
        RECT 596.950 291.170 597.580 291.410 ;
        RECT 608.400 291.350 608.970 291.710 ;
        RECT 622.930 291.630 623.680 291.710 ;
        RECT 639.200 291.610 639.570 291.910 ;
        RECT 639.160 291.360 639.570 291.610 ;
        RECT 607.070 291.170 607.840 291.340 ;
        RECT 596.950 290.800 607.840 291.170 ;
        RECT 596.950 290.460 597.580 290.800 ;
        RECT 607.070 290.600 607.840 290.800 ;
        RECT 608.380 290.650 608.920 290.860 ;
        RECT 621.060 290.650 621.470 290.780 ;
        RECT 608.380 290.480 621.470 290.650 ;
        RECT 608.380 290.340 608.920 290.480 ;
        RECT 621.060 290.390 621.470 290.480 ;
        RECT 622.110 290.720 622.700 290.860 ;
        RECT 633.820 290.720 634.530 290.920 ;
        RECT 622.110 290.410 634.530 290.720 ;
        RECT 622.110 290.300 622.700 290.410 ;
        RECT 631.400 289.730 632.000 290.200 ;
        RECT 633.820 290.140 634.530 290.410 ;
        RECT 639.160 289.610 639.400 291.360 ;
        RECT 645.260 291.230 645.570 291.680 ;
        RECT 641.680 290.800 642.060 291.220 ;
        RECT 639.160 289.560 639.590 289.610 ;
        RECT 645.290 289.570 645.510 291.230 ;
        RECT 709.360 290.800 710.000 290.840 ;
        RECT 711.950 290.800 713.630 291.490 ;
        RECT 642.500 289.560 645.510 289.570 ;
        RECT 594.160 289.020 594.790 289.390 ;
        RECT 603.780 289.240 604.640 289.540 ;
        RECT 609.350 289.240 609.900 289.490 ;
        RECT 639.160 289.390 645.510 289.560 ;
        RECT 642.500 289.370 645.510 289.390 ;
        RECT 603.780 289.030 609.900 289.240 ;
        RECT 591.300 287.120 592.690 288.460 ;
        RECT 296.180 285.870 297.550 286.360 ;
        RECT 302.600 285.870 304.660 286.410 ;
        RECT 296.180 284.780 304.660 285.870 ;
        RECT 296.180 284.200 297.550 284.780 ;
        RECT 302.600 283.850 304.660 284.780 ;
        RECT 594.290 283.920 594.700 289.020 ;
        RECT 603.780 288.880 604.640 289.030 ;
        RECT 609.350 288.820 609.900 289.030 ;
        RECT 621.040 289.180 621.420 289.280 ;
        RECT 629.110 289.180 629.570 289.330 ;
        RECT 621.040 288.990 629.570 289.180 ;
        RECT 639.300 289.170 639.510 289.180 ;
        RECT 621.040 288.900 621.420 288.990 ;
        RECT 629.110 288.880 629.570 288.990 ;
        RECT 639.110 289.040 639.710 289.170 ;
        RECT 641.650 289.040 642.080 289.200 ;
        RECT 639.110 288.830 642.080 289.040 ;
        RECT 639.110 288.710 639.710 288.830 ;
        RECT 641.650 288.670 642.080 288.830 ;
        RECT 643.210 288.590 643.680 289.370 ;
        RECT 694.770 288.500 696.160 290.580 ;
        RECT 709.360 290.300 713.630 290.800 ;
        RECT 645.180 286.880 646.060 287.760 ;
        RECT 709.360 287.440 710.000 290.300 ;
        RECT 711.950 289.980 713.630 290.300 ;
        RECT 728.430 289.750 728.790 291.950 ;
        RECT 729.960 291.900 731.040 291.950 ;
        RECT 713.530 289.410 728.790 289.750 ;
        RECT 713.530 289.380 728.720 289.410 ;
        RECT 603.140 285.110 603.490 285.340 ;
        RECT 610.940 285.110 611.250 285.330 ;
        RECT 602.050 284.580 602.770 284.980 ;
        RECT 603.140 284.930 611.250 285.110 ;
        RECT 603.140 284.800 603.490 284.930 ;
        RECT 610.940 284.890 611.250 284.930 ;
        RECT 620.070 284.860 620.370 285.320 ;
        RECT 620.160 284.640 620.310 284.860 ;
        RECT 628.890 284.640 629.410 284.770 ;
        RECT 620.160 284.440 629.410 284.640 ;
        RECT 628.890 284.320 629.410 284.440 ;
        RECT 645.420 283.970 645.640 286.880 ;
        RECT 695.190 286.870 710.000 287.440 ;
        RECT 695.190 284.350 695.660 286.870 ;
        RECT 636.080 283.950 645.650 283.970 ;
        RECT 613.850 283.920 645.650 283.950 ;
        RECT 594.290 283.620 645.650 283.920 ;
        RECT 594.290 283.540 637.060 283.620 ;
        RECT 594.290 283.510 617.500 283.540 ;
        RECT 591.240 281.580 592.630 282.920 ;
        RECT 695.210 280.020 695.560 284.350 ;
        RECT 683.190 279.060 683.680 279.660 ;
        RECT 694.930 279.170 695.790 280.020 ;
        RECT 713.550 280.010 713.940 289.380 ;
        RECT 726.790 286.450 728.240 287.580 ;
        RECT 700.690 279.150 701.100 279.770 ;
        RECT 713.380 279.170 714.060 280.010 ;
        RECT 727.250 279.910 727.660 286.450 ;
        RECT 765.580 286.180 765.880 297.060 ;
        RECT 854.050 295.590 854.550 295.740 ;
        RECT 852.050 295.300 854.550 295.590 ;
        RECT 843.810 294.080 844.230 294.580 ;
        RECT 843.880 292.870 844.090 294.080 ;
        RECT 843.790 292.190 844.310 292.870 ;
        RECT 849.040 291.730 849.870 292.580 ;
        RECT 820.030 290.420 820.370 290.910 ;
        RECT 820.110 288.990 820.310 290.420 ;
        RECT 820.110 288.830 823.520 288.990 ;
        RECT 779.440 286.680 781.260 287.260 ;
        RECT 779.440 286.660 812.200 286.680 ;
        RECT 814.450 286.660 815.060 286.920 ;
        RECT 779.440 286.410 815.060 286.660 ;
        RECT 747.610 285.610 765.920 286.180 ;
        RECT 779.440 285.700 781.260 286.410 ;
        RECT 811.400 286.390 815.060 286.410 ;
        RECT 814.450 286.170 815.060 286.390 ;
        RECT 747.620 279.970 747.990 285.610 ;
        RECT 816.300 284.500 817.320 285.440 ;
        RECT 819.020 285.350 819.430 285.930 ;
        RECT 799.690 281.250 799.990 281.380 ;
        RECT 797.850 281.220 799.990 281.250 ;
        RECT 797.840 281.060 799.990 281.220 ;
        RECT 718.270 279.220 718.710 279.550 ;
        RECT 154.900 278.150 156.340 278.740 ;
        RECT 157.270 278.150 158.270 278.880 ;
        RECT 154.900 277.620 158.270 278.150 ;
        RECT 632.560 277.660 633.330 278.680 ;
        RECT 154.900 277.100 156.340 277.620 ;
        RECT 157.270 276.990 158.270 277.620 ;
        RECT 679.840 274.340 680.300 274.940 ;
        RECT 683.270 274.530 683.430 279.060 ;
        RECT 700.520 278.970 701.100 279.150 ;
        RECT 718.100 279.000 718.710 279.220 ;
        RECT 727.180 279.150 727.870 279.910 ;
        RECT 735.570 279.310 735.900 279.540 ;
        RECT 735.370 279.100 735.900 279.310 ;
        RECT 747.460 279.130 748.130 279.970 ;
        RECT 608.320 273.470 608.890 273.830 ;
        RECT 622.850 273.470 623.600 273.700 ;
        RECT 608.320 273.240 623.600 273.470 ;
        RECT 596.870 272.700 597.500 272.940 ;
        RECT 608.320 272.880 608.890 273.240 ;
        RECT 622.850 273.160 623.600 273.240 ;
        RECT 639.120 273.140 639.490 273.440 ;
        RECT 639.080 272.890 639.490 273.140 ;
        RECT 606.990 272.700 607.760 272.870 ;
        RECT 596.870 272.330 607.760 272.700 ;
        RECT 596.870 271.990 597.500 272.330 ;
        RECT 606.990 272.130 607.760 272.330 ;
        RECT 608.300 272.180 608.840 272.390 ;
        RECT 620.980 272.180 621.390 272.310 ;
        RECT 608.300 272.010 621.390 272.180 ;
        RECT 608.300 271.870 608.840 272.010 ;
        RECT 620.980 271.920 621.390 272.010 ;
        RECT 622.030 272.250 622.620 272.390 ;
        RECT 633.740 272.250 634.450 272.450 ;
        RECT 622.030 271.940 634.450 272.250 ;
        RECT 622.030 271.830 622.620 271.940 ;
        RECT 631.550 271.140 631.970 271.680 ;
        RECT 633.740 271.670 634.450 271.940 ;
        RECT 639.080 271.140 639.320 272.890 ;
        RECT 645.180 272.760 645.490 273.210 ;
        RECT 641.600 272.330 641.980 272.750 ;
        RECT 639.080 271.090 639.510 271.140 ;
        RECT 645.210 271.100 645.430 272.760 ;
        RECT 642.420 271.090 645.430 271.100 ;
        RECT 594.080 270.550 594.710 270.920 ;
        RECT 603.700 270.770 604.560 271.070 ;
        RECT 609.270 270.770 609.820 271.020 ;
        RECT 639.080 270.920 645.430 271.090 ;
        RECT 642.420 270.900 645.430 270.920 ;
        RECT 603.700 270.560 609.820 270.770 ;
        RECT 591.300 268.930 592.570 270.070 ;
        RECT 594.210 265.450 594.620 270.550 ;
        RECT 603.700 270.410 604.560 270.560 ;
        RECT 609.270 270.350 609.820 270.560 ;
        RECT 620.960 270.710 621.340 270.810 ;
        RECT 629.030 270.710 629.490 270.860 ;
        RECT 620.960 270.520 629.490 270.710 ;
        RECT 639.220 270.700 639.430 270.710 ;
        RECT 620.960 270.430 621.340 270.520 ;
        RECT 629.030 270.410 629.490 270.520 ;
        RECT 639.030 270.570 639.630 270.700 ;
        RECT 641.570 270.570 642.000 270.730 ;
        RECT 639.030 270.360 642.000 270.570 ;
        RECT 639.030 270.240 639.630 270.360 ;
        RECT 641.570 270.200 642.000 270.360 ;
        RECT 643.130 270.120 643.600 270.900 ;
        RECT 645.100 268.410 645.980 269.290 ;
        RECT 680.090 268.710 680.270 274.340 ;
        RECT 681.030 273.790 681.530 274.280 ;
        RECT 683.200 273.930 683.530 274.530 ;
        RECT 685.480 274.080 685.890 274.870 ;
        RECT 700.520 274.600 700.820 278.970 ;
        RECT 603.060 266.640 603.410 266.870 ;
        RECT 610.860 266.640 611.170 266.860 ;
        RECT 601.480 266.100 602.460 266.540 ;
        RECT 603.060 266.460 611.170 266.640 ;
        RECT 603.060 266.330 603.410 266.460 ;
        RECT 610.860 266.420 611.170 266.460 ;
        RECT 619.990 266.390 620.290 266.850 ;
        RECT 620.080 266.170 620.230 266.390 ;
        RECT 628.810 266.170 629.330 266.300 ;
        RECT 620.080 265.970 629.330 266.170 ;
        RECT 628.810 265.850 629.330 265.970 ;
        RECT 645.340 265.500 645.560 268.410 ;
        RECT 680.030 268.170 680.440 268.710 ;
        RECT 681.070 268.540 681.290 273.790 ;
        RECT 685.650 268.760 685.840 274.080 ;
        RECT 686.570 273.390 687.060 274.310 ;
        RECT 692.820 273.680 693.500 274.560 ;
        RECT 700.420 274.380 700.820 274.600 ;
        RECT 698.260 273.810 698.760 274.300 ;
        RECT 700.420 273.950 700.790 274.380 ;
        RECT 702.710 274.100 703.120 274.890 ;
        RECT 718.100 274.600 718.350 279.000 ;
        RECT 686.730 269.610 686.900 273.390 ;
        RECT 680.980 267.930 681.340 268.540 ;
        RECT 685.650 268.530 686.100 268.760 ;
        RECT 686.670 268.710 687.030 269.610 ;
        RECT 685.770 268.180 686.100 268.530 ;
        RECT 686.730 268.480 686.900 268.710 ;
        RECT 686.680 267.800 687.040 268.480 ;
        RECT 636.000 265.480 645.570 265.500 ;
        RECT 613.770 265.450 645.570 265.480 ;
        RECT 594.210 265.150 645.570 265.450 ;
        RECT 594.210 265.070 636.980 265.150 ;
        RECT 594.210 265.040 617.420 265.070 ;
        RECT 693.010 264.750 693.440 273.680 ;
        RECT 698.300 268.560 698.520 273.810 ;
        RECT 702.880 268.780 703.070 274.100 ;
        RECT 703.800 273.410 704.290 274.330 ;
        RECT 710.070 273.590 710.970 274.590 ;
        RECT 715.830 273.910 716.330 274.400 ;
        RECT 718.040 274.120 718.380 274.600 ;
        RECT 720.280 274.200 720.690 274.990 ;
        RECT 698.210 267.950 698.570 268.560 ;
        RECT 702.880 268.550 703.330 268.780 ;
        RECT 703.960 268.680 704.130 273.410 ;
        RECT 703.000 268.200 703.330 268.550 ;
        RECT 703.860 267.720 704.290 268.680 ;
        RECT 591.100 263.540 592.510 264.710 ;
        RECT 692.400 263.450 693.930 264.750 ;
        RECT 710.180 264.740 710.680 273.590 ;
        RECT 711.090 268.690 711.450 269.590 ;
        RECT 715.870 268.660 716.090 273.910 ;
        RECT 720.450 268.880 720.640 274.200 ;
        RECT 721.370 273.510 721.860 274.430 ;
        RECT 727.600 274.270 728.460 274.720 ;
        RECT 735.370 274.590 735.660 279.100 ;
        RECT 753.010 279.080 753.390 279.500 ;
        RECT 735.170 274.440 735.660 274.590 ;
        RECT 727.530 273.820 728.460 274.270 ;
        RECT 733.000 273.940 733.500 274.430 ;
        RECT 735.170 274.150 735.500 274.440 ;
        RECT 737.450 274.230 737.860 275.020 ;
        RECT 721.530 269.840 721.700 273.510 ;
        RECT 715.780 268.050 716.140 268.660 ;
        RECT 720.450 268.650 720.900 268.880 ;
        RECT 721.450 268.860 721.920 269.840 ;
        RECT 720.570 268.300 720.900 268.650 ;
        RECT 721.530 268.600 721.700 268.860 ;
        RECT 721.480 267.920 721.840 268.600 ;
        RECT 694.650 264.140 710.710 264.740 ;
        RECT 727.530 264.250 728.110 273.820 ;
        RECT 728.640 267.870 729.070 268.830 ;
        RECT 733.040 268.690 733.260 273.940 ;
        RECT 737.620 268.910 737.810 274.230 ;
        RECT 738.540 273.540 739.030 274.460 ;
        RECT 744.910 273.790 746.000 274.850 ;
        RECT 753.050 274.630 753.210 279.080 ;
        RECT 797.840 278.320 798.230 281.060 ;
        RECT 799.690 280.980 799.990 281.060 ;
        RECT 802.040 280.510 802.970 281.600 ;
        RECT 797.440 277.390 798.560 278.320 ;
        RECT 797.830 276.780 798.120 277.390 ;
        RECT 816.000 277.260 816.260 277.340 ;
        RECT 816.420 277.260 816.780 284.500 ;
        RECT 818.020 281.290 818.650 281.480 ;
        RECT 819.020 281.290 819.280 285.350 ;
        RECT 823.330 284.260 823.520 288.830 ;
        RECT 833.270 288.600 833.750 289.070 ;
        RECT 833.360 286.340 833.650 288.600 ;
        RECT 840.520 288.100 840.810 288.570 ;
        RECT 840.520 286.880 840.710 288.100 ;
        RECT 840.330 286.410 840.910 286.880 ;
        RECT 832.940 285.250 834.270 286.340 ;
        RECT 840.520 286.230 840.710 286.410 ;
        RECT 823.330 283.930 850.020 284.260 ;
        RECT 821.730 281.290 822.110 281.410 ;
        RECT 841.080 281.370 841.440 281.570 ;
        RECT 818.020 281.060 822.110 281.290 ;
        RECT 839.680 281.220 841.440 281.370 ;
        RECT 818.020 280.830 818.650 281.060 ;
        RECT 821.730 281.020 822.110 281.060 ;
        RECT 820.840 280.740 821.160 280.900 ;
        RECT 818.830 280.730 821.160 280.740 ;
        RECT 818.780 280.530 821.160 280.730 ;
        RECT 818.780 280.520 821.060 280.530 ;
        RECT 818.780 277.260 819.030 280.520 ;
        RECT 828.010 280.200 828.470 280.820 ;
        RECT 829.050 279.950 829.390 280.670 ;
        RECT 836.600 280.490 837.090 280.990 ;
        RECT 829.080 277.260 829.240 279.950 ;
        RECT 836.640 278.750 836.920 280.490 ;
        RECT 836.540 278.130 837.140 278.750 ;
        RECT 839.700 277.270 839.900 281.220 ;
        RECT 841.080 281.160 841.440 281.220 ;
        RECT 849.690 281.060 849.990 283.930 ;
        RECT 840.990 280.190 841.420 280.710 ;
        RECT 849.690 280.620 850.020 281.060 ;
        RECT 852.080 280.920 852.330 295.300 ;
        RECT 854.050 295.170 854.550 295.300 ;
        RECT 856.910 295.080 857.240 295.510 ;
        RECT 857.020 294.270 857.220 295.080 ;
        RECT 852.960 294.030 857.220 294.270 ;
        RECT 852.970 293.830 853.240 294.030 ;
        RECT 852.670 292.930 853.660 293.830 ;
        RECT 852.970 283.900 853.240 292.930 ;
        RECT 868.180 291.640 869.190 292.310 ;
        RECT 856.960 289.570 857.270 290.080 ;
        RECT 857.050 288.480 857.200 289.570 ;
        RECT 852.930 283.170 853.380 283.900 ;
        RECT 857.040 282.660 857.200 288.480 ;
        RECT 853.210 282.650 857.230 282.660 ;
        RECT 853.150 282.470 857.230 282.650 ;
        RECT 849.710 280.540 850.020 280.620 ;
        RECT 841.830 279.780 842.430 280.420 ;
        RECT 840.640 278.750 840.800 279.700 ;
        RECT 840.640 278.650 841.280 278.750 ;
        RECT 840.680 278.170 841.280 278.650 ;
        RECT 836.040 277.260 839.900 277.270 ;
        RECT 816.000 277.060 839.900 277.260 ;
        RECT 797.830 276.600 798.130 276.780 ;
        RECT 816.000 276.720 816.260 277.060 ;
        RECT 836.040 277.050 839.900 277.060 ;
        RECT 816.000 276.630 816.270 276.720 ;
        RECT 750.810 274.000 751.310 274.490 ;
        RECT 752.970 274.210 753.350 274.630 ;
        RECT 755.260 274.290 755.670 275.080 ;
        RECT 732.950 268.080 733.310 268.690 ;
        RECT 737.620 268.680 738.070 268.910 ;
        RECT 737.740 268.330 738.070 268.680 ;
        RECT 738.700 268.660 738.870 273.540 ;
        RECT 745.210 270.200 745.760 273.790 ;
        RECT 745.210 268.930 745.690 270.200 ;
        RECT 745.830 269.830 746.140 270.070 ;
        RECT 745.830 269.070 746.170 269.830 ;
        RECT 745.210 268.690 745.700 268.930 ;
        RECT 745.860 268.830 746.170 269.070 ;
        RECT 750.850 268.750 751.070 274.000 ;
        RECT 755.430 268.970 755.620 274.290 ;
        RECT 762.620 273.900 763.590 274.940 ;
        RECT 797.850 274.500 798.130 276.600 ;
        RECT 816.010 274.630 816.270 276.630 ;
        RECT 834.590 276.050 835.220 276.520 ;
        RECT 834.740 274.650 835.020 276.050 ;
        RECT 738.660 268.630 739.010 268.660 ;
        RECT 738.650 267.950 739.010 268.630 ;
        RECT 738.660 267.900 739.010 267.950 ;
        RECT 745.210 264.270 745.760 268.690 ;
        RECT 750.760 268.140 751.120 268.750 ;
        RECT 755.430 268.740 755.880 268.970 ;
        RECT 755.550 268.390 755.880 268.740 ;
        RECT 694.620 263.800 710.710 264.140 ;
        RECT 693.030 261.670 693.870 262.630 ;
        RECT 632.390 260.110 633.530 260.910 ;
        RECT 683.170 257.530 683.660 258.130 ;
        RECT 608.170 255.740 608.740 256.100 ;
        RECT 622.700 255.740 623.450 255.970 ;
        RECT 608.170 255.510 623.450 255.740 ;
        RECT 596.720 254.970 597.350 255.210 ;
        RECT 608.170 255.150 608.740 255.510 ;
        RECT 622.700 255.430 623.450 255.510 ;
        RECT 638.970 255.410 639.340 255.710 ;
        RECT 638.930 255.160 639.340 255.410 ;
        RECT 606.840 254.970 607.610 255.140 ;
        RECT 596.720 254.600 607.610 254.970 ;
        RECT 596.720 254.260 597.350 254.600 ;
        RECT 606.840 254.400 607.610 254.600 ;
        RECT 608.150 254.450 608.690 254.660 ;
        RECT 620.830 254.450 621.240 254.580 ;
        RECT 608.150 254.280 621.240 254.450 ;
        RECT 608.150 254.140 608.690 254.280 ;
        RECT 620.830 254.190 621.240 254.280 ;
        RECT 621.880 254.520 622.470 254.660 ;
        RECT 633.590 254.520 634.300 254.720 ;
        RECT 621.880 254.210 634.300 254.520 ;
        RECT 621.880 254.100 622.470 254.210 ;
        RECT 631.360 253.480 631.930 254.000 ;
        RECT 633.590 253.940 634.300 254.210 ;
        RECT 638.930 253.410 639.170 255.160 ;
        RECT 645.030 255.030 645.340 255.480 ;
        RECT 641.450 254.600 641.830 255.020 ;
        RECT 638.930 253.360 639.360 253.410 ;
        RECT 645.060 253.370 645.280 255.030 ;
        RECT 642.270 253.360 645.280 253.370 ;
        RECT 593.930 252.820 594.560 253.190 ;
        RECT 603.550 253.040 604.410 253.340 ;
        RECT 609.120 253.040 609.670 253.290 ;
        RECT 638.930 253.190 645.280 253.360 ;
        RECT 642.270 253.170 645.280 253.190 ;
        RECT 603.550 252.830 609.670 253.040 ;
        RECT 591.240 250.110 592.190 251.650 ;
        RECT 594.060 247.720 594.470 252.820 ;
        RECT 603.550 252.680 604.410 252.830 ;
        RECT 609.120 252.620 609.670 252.830 ;
        RECT 620.810 252.980 621.190 253.080 ;
        RECT 628.880 252.980 629.340 253.130 ;
        RECT 620.810 252.790 629.340 252.980 ;
        RECT 639.070 252.970 639.280 252.980 ;
        RECT 620.810 252.700 621.190 252.790 ;
        RECT 628.880 252.680 629.340 252.790 ;
        RECT 638.880 252.840 639.480 252.970 ;
        RECT 641.420 252.840 641.850 253.000 ;
        RECT 638.880 252.630 641.850 252.840 ;
        RECT 638.880 252.510 639.480 252.630 ;
        RECT 641.420 252.470 641.850 252.630 ;
        RECT 642.980 252.390 643.450 253.170 ;
        RECT 683.250 253.000 683.410 257.530 ;
        RECT 681.010 252.260 681.510 252.750 ;
        RECT 683.180 252.400 683.510 253.000 ;
        RECT 685.460 252.550 685.870 253.340 ;
        RECT 693.320 253.190 693.600 261.670 ;
        RECT 694.620 258.470 694.850 263.800 ;
        RECT 712.860 263.750 728.110 264.250 ;
        RECT 694.480 257.740 695.090 258.470 ;
        RECT 712.870 258.450 713.360 263.750 ;
        RECT 727.530 263.650 728.110 263.750 ;
        RECT 730.160 263.820 745.760 264.270 ;
        RECT 762.690 264.240 763.390 273.900 ;
        RECT 797.530 273.570 798.410 274.500 ;
        RECT 815.820 273.760 816.650 274.630 ;
        RECT 834.600 273.980 835.070 274.650 ;
        RECT 836.080 272.910 836.260 277.050 ;
        RECT 839.700 277.030 839.900 277.050 ;
        RECT 849.710 276.660 849.980 280.540 ;
        RECT 851.940 280.140 852.650 280.920 ;
        RECT 853.150 278.160 853.370 282.470 ;
        RECT 865.220 281.150 865.980 282.210 ;
        RECT 857.040 278.810 857.340 279.340 ;
        RECT 853.060 277.510 853.520 278.160 ;
        RECT 857.130 276.950 857.270 278.810 ;
        RECT 851.070 276.690 857.280 276.950 ;
        RECT 844.000 276.390 849.980 276.660 ;
        RECT 837.020 273.390 837.450 274.100 ;
        RECT 836.770 272.910 837.460 273.130 ;
        RECT 784.370 272.200 784.700 272.650 ;
        RECT 784.480 271.050 784.680 272.200 ;
        RECT 803.300 272.190 803.580 272.740 ;
        RECT 836.080 272.710 837.460 272.910 ;
        RECT 822.140 272.230 822.420 272.710 ;
        RECT 836.770 272.610 837.460 272.710 ;
        RECT 784.180 270.370 784.950 271.050 ;
        RECT 803.320 271.020 803.560 272.190 ;
        RECT 802.970 270.450 803.860 271.020 ;
        RECT 822.170 270.970 822.360 272.230 ;
        RECT 822.090 270.440 822.520 270.970 ;
        RECT 763.670 268.230 764.020 268.990 ;
        RECT 797.610 268.350 798.470 269.390 ;
        RECT 797.780 267.340 798.070 268.350 ;
        RECT 836.900 267.350 837.370 267.870 ;
        RECT 797.550 266.480 798.400 267.340 ;
        RECT 816.130 266.950 816.980 267.240 ;
        RECT 821.650 266.950 822.590 267.240 ;
        RECT 816.130 266.540 822.590 266.950 ;
        RECT 816.130 266.380 816.980 266.540 ;
        RECT 821.650 266.200 822.590 266.540 ;
        RECT 837.060 266.960 837.680 267.070 ;
        RECT 839.520 266.980 839.810 267.130 ;
        RECT 844.000 266.980 844.320 276.390 ;
        RECT 851.090 267.720 851.380 276.690 ;
        RECT 853.000 271.460 853.500 272.130 ;
        RECT 853.080 270.610 853.360 271.460 ;
        RECT 839.520 266.960 844.330 266.980 ;
        RECT 837.060 266.740 844.330 266.960 ;
        RECT 850.870 266.950 851.700 267.720 ;
        RECT 837.060 266.490 837.680 266.740 ;
        RECT 839.520 266.640 839.810 266.740 ;
        RECT 844.000 266.700 844.320 266.740 ;
        RECT 853.080 266.080 853.380 270.610 ;
        RECT 853.100 265.360 853.380 266.080 ;
        RECT 784.420 264.690 784.700 265.200 ;
        RECT 802.950 264.730 803.220 265.230 ;
        RECT 853.100 265.040 853.580 265.360 ;
        RECT 853.130 264.740 853.580 265.040 ;
        RECT 747.780 264.000 763.390 264.240 ;
        RECT 730.160 263.720 745.730 263.820 ;
        RECT 730.190 258.470 730.500 263.720 ;
        RECT 747.760 263.700 763.390 264.000 ;
        RECT 747.760 258.470 748.110 263.700 ;
        RECT 762.690 263.610 763.390 263.700 ;
        RECT 784.480 263.190 784.670 264.690 ;
        RECT 802.970 263.520 803.160 264.730 ;
        RECT 784.200 262.500 784.950 263.190 ;
        RECT 802.590 262.820 803.680 263.520 ;
        RECT 850.870 261.460 851.800 262.320 ;
        RECT 852.520 261.730 853.210 262.470 ;
        RECT 700.670 257.620 701.080 258.240 ;
        RECT 712.750 257.790 713.490 258.450 ;
        RECT 718.250 257.690 718.690 258.020 ;
        RECT 729.930 257.740 730.700 258.470 ;
        RECT 735.550 257.780 735.880 258.010 ;
        RECT 700.500 257.440 701.080 257.620 ;
        RECT 718.080 257.470 718.690 257.690 ;
        RECT 735.350 257.570 735.880 257.780 ;
        RECT 747.500 257.740 748.310 258.470 ;
        RECT 846.620 258.140 847.450 259.340 ;
        RECT 644.950 250.680 645.830 251.560 ;
        RECT 602.910 248.910 603.260 249.140 ;
        RECT 610.710 248.910 611.020 249.130 ;
        RECT 602.910 248.730 611.020 248.910 ;
        RECT 602.910 248.600 603.260 248.730 ;
        RECT 610.710 248.690 611.020 248.730 ;
        RECT 619.840 248.660 620.140 249.120 ;
        RECT 619.930 248.440 620.080 248.660 ;
        RECT 628.660 248.440 629.180 248.570 ;
        RECT 619.930 248.240 629.180 248.440 ;
        RECT 628.660 248.120 629.180 248.240 ;
        RECT 645.190 247.770 645.410 250.680 ;
        RECT 635.850 247.750 645.420 247.770 ;
        RECT 613.620 247.720 645.420 247.750 ;
        RECT 594.060 247.420 645.420 247.720 ;
        RECT 594.060 247.340 636.830 247.420 ;
        RECT 594.060 247.310 617.270 247.340 ;
        RECT 681.050 247.010 681.270 252.260 ;
        RECT 685.630 247.230 685.820 252.550 ;
        RECT 686.550 251.860 687.040 252.780 ;
        RECT 693.290 252.070 694.050 253.190 ;
        RECT 700.500 253.070 700.800 257.440 ;
        RECT 700.400 252.850 700.800 253.070 ;
        RECT 698.240 252.280 698.740 252.770 ;
        RECT 700.400 252.420 700.770 252.850 ;
        RECT 702.690 252.570 703.100 253.360 ;
        RECT 718.080 253.070 718.330 257.470 ;
        RECT 686.710 248.080 686.880 251.860 ;
        RECT 680.960 246.400 681.320 247.010 ;
        RECT 685.630 247.000 686.080 247.230 ;
        RECT 686.650 247.180 687.010 248.080 ;
        RECT 685.750 246.650 686.080 247.000 ;
        RECT 686.710 246.950 686.880 247.180 ;
        RECT 698.280 247.030 698.500 252.280 ;
        RECT 702.860 247.250 703.050 252.570 ;
        RECT 703.780 251.880 704.270 252.800 ;
        RECT 710.330 252.120 711.190 252.950 ;
        RECT 715.810 252.380 716.310 252.870 ;
        RECT 718.020 252.590 718.360 253.070 ;
        RECT 720.260 252.670 720.670 253.460 ;
        RECT 735.350 253.060 735.640 257.570 ;
        RECT 752.990 257.550 753.370 257.970 ;
        RECT 745.580 256.190 745.850 256.320 ;
        RECT 751.670 256.190 752.250 256.370 ;
        RECT 745.580 255.940 752.250 256.190 ;
        RECT 735.150 252.910 735.640 253.060 ;
        RECT 686.660 246.270 687.020 246.950 ;
        RECT 698.190 246.420 698.550 247.030 ;
        RECT 702.860 247.020 703.310 247.250 ;
        RECT 703.940 247.150 704.110 251.880 ;
        RECT 711.070 247.160 711.430 248.060 ;
        RECT 702.980 246.670 703.310 247.020 ;
        RECT 703.840 246.190 704.270 247.150 ;
        RECT 715.850 247.130 716.070 252.380 ;
        RECT 720.430 247.350 720.620 252.670 ;
        RECT 721.350 251.980 721.840 252.900 ;
        RECT 732.980 252.410 733.480 252.900 ;
        RECT 735.150 252.620 735.480 252.910 ;
        RECT 737.430 252.700 737.840 253.490 ;
        RECT 745.580 253.120 745.850 255.940 ;
        RECT 751.670 255.670 752.250 255.940 ;
        RECT 721.510 248.310 721.680 251.980 ;
        RECT 715.760 246.520 716.120 247.130 ;
        RECT 720.430 247.120 720.880 247.350 ;
        RECT 721.430 247.330 721.900 248.310 ;
        RECT 720.550 246.770 720.880 247.120 ;
        RECT 721.510 247.070 721.680 247.330 ;
        RECT 721.460 246.390 721.820 247.070 ;
        RECT 728.620 246.340 729.050 247.300 ;
        RECT 733.020 247.160 733.240 252.410 ;
        RECT 737.600 247.380 737.790 252.700 ;
        RECT 738.520 252.010 739.010 252.930 ;
        RECT 745.320 252.440 745.910 253.120 ;
        RECT 753.030 253.100 753.190 257.550 ;
        RECT 776.160 257.360 776.990 257.750 ;
        RECT 846.790 257.360 847.110 258.140 ;
        RECT 851.090 257.610 851.380 261.460 ;
        RECT 851.090 257.410 851.430 257.610 ;
        RECT 776.160 256.980 847.110 257.360 ;
        RECT 776.160 256.760 776.990 256.980 ;
        RECT 846.790 256.920 847.110 256.980 ;
        RECT 851.110 256.690 851.430 257.410 ;
        RECT 852.700 256.910 852.870 261.730 ;
        RECT 853.400 261.170 853.870 261.700 ;
        RECT 853.540 259.280 853.760 261.170 ;
        RECT 853.360 258.690 853.890 259.280 ;
        RECT 856.040 256.910 856.370 257.060 ;
        RECT 852.680 256.750 856.370 256.910 ;
        RECT 852.700 256.730 852.870 256.750 ;
        RECT 850.970 255.710 851.670 256.690 ;
        RECT 856.040 256.660 856.370 256.750 ;
        RECT 852.730 254.580 853.460 255.490 ;
        RECT 750.790 252.470 751.290 252.960 ;
        RECT 752.950 252.680 753.330 253.100 ;
        RECT 755.240 252.760 755.650 253.550 ;
        RECT 866.340 252.870 867.280 253.760 ;
        RECT 732.930 246.550 733.290 247.160 ;
        RECT 737.600 247.150 738.050 247.380 ;
        RECT 737.720 246.800 738.050 247.150 ;
        RECT 738.680 247.130 738.850 252.010 ;
        RECT 745.810 248.300 746.120 248.540 ;
        RECT 745.810 247.540 746.150 248.300 ;
        RECT 745.840 247.300 746.150 247.540 ;
        RECT 750.830 247.220 751.050 252.470 ;
        RECT 755.410 247.440 755.600 252.760 ;
        RECT 857.050 250.480 857.380 250.990 ;
        RECT 857.080 249.180 857.310 250.480 ;
        RECT 856.920 248.500 857.510 249.180 ;
        RECT 738.640 247.100 738.990 247.130 ;
        RECT 738.630 246.420 738.990 247.100 ;
        RECT 750.740 246.610 751.100 247.220 ;
        RECT 755.410 247.210 755.860 247.440 ;
        RECT 755.530 246.860 755.860 247.210 ;
        RECT 763.650 246.700 764.000 247.460 ;
        RECT 738.640 246.370 738.990 246.420 ;
        RECT 378.620 236.490 381.840 239.000 ;
        RECT 334.120 232.890 336.220 233.490 ;
        RECT 365.300 232.890 368.370 234.460 ;
        RECT 334.120 231.060 368.370 232.890 ;
        RECT 334.120 229.820 336.220 231.060 ;
        RECT 365.300 230.050 368.370 231.060 ;
        RECT 379.420 229.520 380.940 236.490 ;
        RECT 379.280 229.290 384.790 229.520 ;
        RECT 389.610 229.290 393.820 230.020 ;
        RECT 379.140 228.250 393.820 229.290 ;
        RECT 379.280 227.800 393.820 228.250 ;
        RECT 379.280 225.900 380.910 227.800 ;
        RECT 381.990 227.720 393.820 227.800 ;
        RECT 389.610 226.400 393.820 227.720 ;
        RECT 379.280 225.380 381.140 225.900 ;
        RECT 379.280 225.270 380.940 225.380 ;
        RECT 379.330 217.320 380.940 225.270 ;
        RECT 395.850 217.320 399.350 217.940 ;
        RECT 379.330 216.000 399.350 217.320 ;
        RECT 379.330 215.950 380.940 216.000 ;
        RECT 395.850 215.500 399.350 216.000 ;
        RECT 395.850 215.470 398.040 215.500 ;
        RECT 398.990 215.470 399.350 215.500 ;
      LAYER via2 ;
        RECT 839.045 353.255 839.325 353.535 ;
        RECT 653.020 352.300 653.300 352.580 ;
        RECT 672.040 352.495 672.320 352.775 ;
        RECT 690.130 352.450 690.410 352.730 ;
        RECT 707.695 352.525 707.975 352.805 ;
        RECT 725.565 352.505 725.845 352.785 ;
        RECT 743.825 352.570 744.105 352.850 ;
        RECT 761.580 352.540 761.860 352.820 ;
        RECT 779.590 352.480 779.870 352.760 ;
        RECT 797.750 352.550 798.030 352.830 ;
        RECT 816.130 352.565 816.410 352.845 ;
        RECT 656.235 349.970 656.515 350.250 ;
        RECT 656.235 349.570 656.515 349.850 ;
        RECT 828.995 349.890 829.275 350.170 ;
        RECT 780.220 343.520 780.900 344.600 ;
        RECT 824.870 343.595 825.150 343.875 ;
        RECT 194.385 334.735 199.465 338.615 ;
        RECT 851.390 337.640 851.670 337.920 ;
        RECT 632.390 333.635 633.070 334.315 ;
        RECT 663.355 329.780 663.635 330.060 ;
        RECT 664.320 329.490 664.600 329.770 ;
        RECT 668.885 329.800 669.165 330.080 ;
        RECT 669.920 329.525 670.200 329.805 ;
        RECT 682.245 329.590 682.525 329.870 ;
        RECT 683.200 329.405 683.480 329.685 ;
        RECT 631.885 327.120 632.165 327.400 ;
        RECT 869.755 333.120 870.435 333.800 ;
        RECT 641.930 328.220 642.210 328.500 ;
        RECT 663.405 326.980 663.685 327.260 ;
        RECT 664.450 326.835 664.730 327.115 ;
        RECT 591.435 320.085 592.515 321.165 ;
        RECT 641.925 326.145 642.205 326.425 ;
        RECT 602.480 321.910 602.760 322.190 ;
        RECT 657.795 323.975 658.075 324.255 ;
        RECT 657.795 323.575 658.075 323.855 ;
        RECT 665.605 323.810 665.885 324.090 ;
        RECT 665.605 323.410 665.885 323.690 ;
        RECT 667.145 323.845 667.425 324.125 ;
        RECT 667.545 323.845 667.825 324.125 ;
        RECT 670.140 323.780 670.420 324.060 ;
        RECT 671.795 323.940 672.075 324.220 ;
        RECT 671.795 323.540 672.075 323.820 ;
        RECT 656.980 322.870 657.260 323.150 ;
        RECT 656.980 322.470 657.260 322.750 ;
        RECT 682.185 323.830 682.465 324.110 ;
        RECT 632.725 315.720 633.005 316.000 ;
        RECT 633.125 315.720 633.405 316.000 ;
        RECT 668.315 318.205 668.595 318.485 ;
        RECT 671.405 318.170 671.685 318.450 ;
        RECT 682.185 323.430 682.465 323.710 ;
        RECT 683.135 323.320 683.415 323.600 ;
        RECT 885.560 322.890 888.640 324.370 ;
        RECT 631.735 308.875 632.015 309.155 ;
        RECT 632.135 308.875 632.415 309.155 ;
        RECT 641.780 310.050 642.060 310.330 ;
        RECT 591.560 306.035 592.640 307.115 ;
        RECT 641.775 307.975 642.055 308.255 ;
        RECT 666.345 308.015 667.425 309.095 ;
        RECT 602.300 303.850 602.580 304.130 ;
        RECT 794.665 305.105 795.745 306.185 ;
        RECT 591.600 300.625 592.680 301.705 ;
        RECT 632.690 296.225 633.370 296.905 ;
        RECT 695.000 297.080 695.280 297.360 ;
        RECT 712.495 297.465 712.775 297.745 ;
        RECT 712.495 297.065 712.775 297.345 ;
        RECT 730.085 297.435 730.365 297.715 ;
        RECT 730.085 297.035 730.365 297.315 ;
        RECT 747.805 297.550 748.085 297.830 ;
        RECT 747.805 297.150 748.085 297.430 ;
        RECT 729.960 292.135 730.240 292.415 ;
        RECT 730.360 292.135 730.640 292.415 ;
        RECT 730.760 292.135 731.040 292.415 ;
        RECT 631.560 289.825 631.840 290.105 ;
        RECT 641.730 290.870 642.010 291.150 ;
        RECT 591.455 287.250 592.535 288.330 ;
        RECT 302.690 283.990 304.570 286.270 ;
        RECT 641.725 288.795 642.005 289.075 ;
        RECT 694.925 288.600 696.005 290.480 ;
        RECT 712.050 290.195 713.530 291.275 ;
        RECT 602.070 284.640 602.350 284.920 ;
        RECT 602.470 284.640 602.750 284.920 ;
        RECT 591.395 281.710 592.475 282.790 ;
        RECT 726.975 286.675 728.055 287.355 ;
        RECT 849.115 291.815 849.795 292.495 ;
        RECT 779.610 285.940 781.090 287.020 ;
        RECT 157.430 277.195 158.110 278.675 ;
        RECT 632.605 277.830 633.285 278.510 ;
        RECT 631.620 271.270 631.900 271.550 ;
        RECT 641.650 272.400 641.930 272.680 ;
        RECT 591.395 269.160 592.475 269.840 ;
        RECT 641.645 270.325 641.925 270.605 ;
        RECT 601.630 266.180 601.910 266.460 ;
        RECT 602.030 266.180 602.310 266.460 ;
        RECT 686.710 269.220 686.990 269.500 ;
        RECT 686.710 268.820 686.990 269.100 ;
        RECT 703.935 268.260 704.215 268.540 ;
        RECT 703.935 267.860 704.215 268.140 ;
        RECT 591.265 263.785 592.345 264.465 ;
        RECT 711.130 269.200 711.410 269.480 ;
        RECT 711.130 268.800 711.410 269.080 ;
        RECT 721.545 269.410 721.825 269.690 ;
        RECT 721.545 269.010 721.825 269.290 ;
        RECT 802.165 280.715 802.845 281.395 ;
        RECT 797.460 277.515 798.540 278.195 ;
        RECT 818.195 281.015 818.475 281.295 ;
        RECT 833.065 285.455 834.145 286.135 ;
        RECT 828.100 280.370 828.380 280.650 ;
        RECT 836.705 280.600 836.985 280.880 ;
        RECT 868.345 291.835 868.625 292.115 ;
        RECT 868.745 291.835 869.025 292.115 ;
        RECT 841.065 280.310 841.345 280.590 ;
        RECT 841.990 279.960 842.270 280.240 ;
        RECT 840.840 278.320 841.120 278.600 ;
        RECT 728.715 268.410 728.995 268.690 ;
        RECT 728.715 268.010 728.995 268.290 ;
        RECT 745.845 269.630 746.125 269.910 ;
        RECT 745.845 269.230 746.125 269.510 ;
        RECT 738.695 268.140 738.975 268.420 ;
        RECT 693.110 261.810 693.790 262.490 ;
        RECT 632.420 260.170 633.500 260.850 ;
        RECT 631.505 253.600 631.785 253.880 ;
        RECT 641.500 254.670 641.780 254.950 ;
        RECT 591.375 250.340 592.055 251.420 ;
        RECT 641.495 252.595 641.775 252.875 ;
        RECT 865.260 281.340 865.940 282.020 ;
        RECT 837.095 273.605 837.375 273.885 ;
        RECT 784.225 270.570 784.505 270.850 ;
        RECT 784.625 270.570 784.905 270.850 ;
        RECT 803.075 270.595 803.355 270.875 ;
        RECT 803.475 270.595 803.755 270.875 ;
        RECT 763.705 268.470 763.985 268.750 ;
        RECT 797.700 268.530 798.380 269.210 ;
        RECT 836.995 267.470 837.275 267.750 ;
        RECT 821.780 266.380 822.460 267.060 ;
        RECT 837.230 266.640 837.510 266.920 ;
        RECT 784.235 262.705 784.515 262.985 ;
        RECT 784.635 262.705 784.915 262.985 ;
        RECT 802.595 263.030 802.875 263.310 ;
        RECT 802.995 263.030 803.275 263.310 ;
        RECT 803.395 263.030 803.675 263.310 ;
        RECT 686.690 247.690 686.970 247.970 ;
        RECT 686.690 247.290 686.970 247.570 ;
        RECT 710.420 252.195 711.100 252.875 ;
        RECT 711.110 247.670 711.390 247.950 ;
        RECT 711.110 247.270 711.390 247.550 ;
        RECT 721.525 247.880 721.805 248.160 ;
        RECT 721.525 247.480 721.805 247.760 ;
        RECT 703.915 246.730 704.195 247.010 ;
        RECT 703.915 246.330 704.195 246.610 ;
        RECT 776.235 256.915 776.915 257.595 ;
        RECT 852.755 254.695 853.435 255.375 ;
        RECT 866.470 252.975 867.150 253.655 ;
        RECT 728.695 246.880 728.975 247.160 ;
        RECT 728.695 246.480 728.975 246.760 ;
        RECT 745.825 248.100 746.105 248.380 ;
        RECT 745.825 247.700 746.105 247.980 ;
        RECT 738.675 246.610 738.955 246.890 ;
        RECT 763.685 246.940 763.965 247.220 ;
        RECT 389.775 226.470 393.655 229.950 ;
      LAYER met3 ;
        RECT 838.950 353.620 839.420 353.685 ;
        RECT 672.050 353.580 839.420 353.620 ;
        RECT 672.040 353.300 839.420 353.580 ;
        RECT 672.040 353.290 744.070 353.300 ;
        RECT 744.490 353.290 839.420 353.300 ;
        RECT 672.040 352.955 672.360 353.290 ;
        RECT 652.850 352.125 653.470 352.755 ;
        RECT 671.880 352.315 672.480 352.955 ;
        RECT 690.060 352.905 690.370 353.290 ;
        RECT 707.660 352.985 707.960 353.290 ;
        RECT 690.010 352.275 690.530 352.905 ;
        RECT 707.590 352.345 708.080 352.985 ;
        RECT 725.530 352.915 725.840 353.290 ;
        RECT 743.740 352.995 744.070 353.290 ;
        RECT 725.470 352.375 725.940 352.915 ;
        RECT 743.740 352.425 744.190 352.995 ;
        RECT 761.480 352.955 761.820 353.290 ;
        RECT 761.470 352.405 761.970 352.955 ;
        RECT 779.590 352.875 779.890 353.290 ;
        RECT 797.730 352.925 798.030 353.290 ;
        RECT 816.160 352.955 816.460 353.290 ;
        RECT 838.950 353.105 839.420 353.290 ;
        RECT 725.490 352.355 725.870 352.375 ;
        RECT 779.490 352.365 779.970 352.875 ;
        RECT 797.630 352.455 798.150 352.925 ;
        RECT 816.020 352.455 816.520 352.955 ;
        RECT 652.920 349.190 653.270 352.125 ;
        RECT 656.010 349.505 656.740 350.315 ;
        RECT 828.750 349.675 829.520 350.385 ;
        RECT 828.890 349.200 829.240 349.675 ;
        RECT 656.410 349.190 829.240 349.200 ;
        RECT 652.870 348.890 829.240 349.190 ;
        RECT 652.870 348.870 656.600 348.890 ;
        RECT 824.260 348.880 825.280 348.890 ;
        RECT 824.360 347.710 825.330 348.180 ;
        RECT 195.120 341.250 198.160 346.540 ;
        RECT 780.070 343.365 781.050 344.755 ;
        RECT 824.820 344.035 825.130 347.710 ;
        RECT 824.750 343.435 825.270 344.035 ;
        RECT 780.500 342.350 781.000 343.365 ;
        RECT 632.640 341.980 781.000 342.350 ;
        RECT 632.610 341.530 781.000 341.980 ;
        RECT 632.610 341.500 780.970 341.530 ;
        RECT 195.920 338.675 197.440 341.250 ;
        RECT 194.190 334.675 199.660 338.675 ;
        RECT 632.610 334.355 633.090 341.500 ;
        RECT 851.220 337.445 851.840 338.115 ;
        RECT 851.490 337.030 851.790 337.445 ;
        RECT 865.000 337.030 868.990 337.040 ;
        RECT 869.850 337.030 870.220 337.050 ;
        RECT 851.480 336.690 870.220 337.030 ;
        RECT 865.000 336.680 868.990 336.690 ;
        RECT 632.200 333.595 633.260 334.355 ;
        RECT 869.850 333.835 870.220 336.690 ;
        RECT 631.640 326.995 632.410 327.525 ;
        RECT 602.280 321.845 602.960 322.255 ;
        RECT 591.290 319.945 592.660 321.305 ;
        RECT 602.480 320.470 602.800 321.845 ;
        RECT 591.810 319.500 592.400 319.945 ;
        RECT 602.450 319.500 602.830 320.470 ;
        RECT 591.760 319.000 602.830 319.500 ;
        RECT 631.860 319.430 632.210 326.995 ;
        RECT 591.810 318.390 592.400 319.000 ;
        RECT 602.450 318.960 602.830 319.000 ;
        RECT 630.920 318.800 632.210 319.430 ;
        RECT 632.730 319.400 633.080 333.595 ;
        RECT 869.670 333.085 870.520 333.835 ;
        RECT 663.250 329.635 663.740 330.205 ;
        RECT 641.830 328.175 642.310 328.545 ;
        RECT 641.910 326.525 642.230 328.175 ;
        RECT 663.420 327.415 663.730 329.635 ;
        RECT 664.200 329.630 664.720 329.865 ;
        RECT 668.760 329.655 669.290 330.225 ;
        RECT 664.200 329.395 664.730 329.630 ;
        RECT 663.250 326.825 663.840 327.415 ;
        RECT 664.400 327.285 664.730 329.395 ;
        RECT 668.800 328.250 669.170 329.655 ;
        RECT 669.800 329.650 670.320 329.955 ;
        RECT 682.080 329.730 682.690 330.025 ;
        RECT 669.800 329.375 670.330 329.650 ;
        RECT 665.530 327.950 669.220 328.250 ;
        RECT 664.210 326.665 664.970 327.285 ;
        RECT 650.550 326.530 653.620 326.540 ;
        RECT 641.800 326.520 642.330 326.525 ;
        RECT 650.550 326.520 653.630 326.530 ;
        RECT 641.800 326.120 653.680 326.520 ;
        RECT 641.800 326.045 642.330 326.120 ;
        RECT 650.550 326.110 653.680 326.120 ;
        RECT 653.360 324.080 653.680 326.110 ;
        RECT 657.550 324.080 658.320 324.355 ;
        RECT 665.570 324.135 665.930 327.950 ;
        RECT 653.360 323.750 658.320 324.080 ;
        RECT 657.550 323.475 658.320 323.750 ;
        RECT 665.420 323.365 666.070 324.135 ;
        RECT 667.010 323.675 667.960 324.295 ;
        RECT 669.980 324.245 670.330 329.375 ;
        RECT 682.040 329.435 682.690 329.730 ;
        RECT 656.840 322.950 657.400 323.205 ;
        RECT 653.760 322.610 657.400 322.950 ;
        RECT 591.800 318.180 592.400 318.390 ;
        RECT 591.800 307.185 592.360 318.180 ;
        RECT 631.860 317.780 632.210 318.800 ;
        RECT 632.610 318.630 633.860 319.400 ;
        RECT 631.860 317.490 632.220 317.780 ;
        RECT 631.880 309.345 632.220 317.490 ;
        RECT 632.730 316.610 633.080 318.630 ;
        RECT 632.720 316.205 633.080 316.610 ;
        RECT 632.590 315.515 633.540 316.205 ;
        RECT 632.720 315.100 633.080 315.515 ;
        RECT 632.730 309.650 633.080 315.100 ;
        RECT 641.680 310.005 642.160 310.375 ;
        RECT 631.670 309.010 632.480 309.345 ;
        RECT 631.600 308.685 632.480 309.010 ;
        RECT 591.500 305.965 592.700 307.185 ;
        RECT 602.090 303.755 602.790 304.225 ;
        RECT 591.540 301.290 592.740 301.775 ;
        RECT 602.210 301.290 602.550 303.755 ;
        RECT 591.540 300.830 602.560 301.290 ;
        RECT 591.540 300.555 592.740 300.830 ;
        RECT 591.700 289.600 592.290 300.555 ;
        RECT 631.600 290.175 632.070 308.685 ;
        RECT 632.780 308.390 633.080 309.650 ;
        RECT 632.730 296.945 633.080 308.390 ;
        RECT 641.760 308.355 642.080 310.005 ;
        RECT 641.650 308.320 642.180 308.355 ;
        RECT 648.500 308.320 649.220 308.360 ;
        RECT 641.650 308.260 650.050 308.320 ;
        RECT 653.780 308.260 654.220 322.610 ;
        RECT 656.840 322.415 657.400 322.610 ;
        RECT 657.190 313.850 657.790 313.870 ;
        RECT 667.340 313.850 667.670 323.675 ;
        RECT 669.940 323.595 670.620 324.245 ;
        RECT 671.630 324.130 672.240 324.255 ;
        RECT 682.040 324.145 682.490 329.435 ;
        RECT 683.080 329.295 683.600 329.795 ;
        RECT 682.020 324.130 682.630 324.145 ;
        RECT 671.630 323.790 682.630 324.130 ;
        RECT 671.630 323.505 672.240 323.790 ;
        RECT 682.020 323.395 682.630 323.790 ;
        RECT 683.180 323.765 683.510 329.295 ;
        RECT 683.020 323.155 683.530 323.765 ;
        RECT 683.170 320.950 683.490 323.155 ;
        RECT 885.340 322.715 888.860 324.545 ;
        RECT 682.060 320.940 683.490 320.950 ;
        RECT 671.390 320.820 683.490 320.940 ;
        RECT 671.380 320.630 683.490 320.820 ;
        RECT 671.380 320.600 683.440 320.630 ;
        RECT 671.380 320.590 682.210 320.600 ;
        RECT 668.180 318.300 668.730 318.645 ;
        RECT 671.380 318.575 671.700 320.590 ;
        RECT 668.170 318.260 668.730 318.300 ;
        RECT 668.000 317.960 668.900 318.260 ;
        RECT 671.290 318.045 671.800 318.575 ;
        RECT 668.170 317.540 668.900 317.960 ;
        RECT 657.160 313.350 667.690 313.850 ;
        RECT 641.650 307.930 654.220 308.260 ;
        RECT 641.650 307.875 642.180 307.930 ;
        RECT 648.500 307.900 649.220 307.930 ;
        RECT 653.780 307.840 654.220 307.930 ;
        RECT 657.190 306.820 657.790 313.350 ;
        RECT 667.340 313.340 667.670 313.350 ;
        RECT 668.170 311.700 668.720 317.540 ;
        RECT 660.050 311.690 668.720 311.700 ;
        RECT 659.960 311.130 668.720 311.690 ;
        RECT 657.230 306.280 657.790 306.820 ;
        RECT 659.970 311.070 668.720 311.130 ;
        RECT 632.510 296.185 633.550 296.945 ;
        RECT 631.350 289.960 632.070 290.175 ;
        RECT 631.350 289.755 632.050 289.960 ;
        RECT 591.690 289.290 592.290 289.600 ;
        RECT 591.690 288.435 592.280 289.290 ;
        RECT 591.250 287.145 592.740 288.435 ;
        RECT 302.550 285.740 304.710 286.385 ;
        RECT 305.140 285.740 306.910 286.180 ;
        RECT 302.550 284.640 306.910 285.740 ;
        RECT 602.000 284.810 602.820 284.955 ;
        RECT 302.550 283.875 304.710 284.640 ;
        RECT 305.140 283.900 306.910 284.640 ;
        RECT 601.930 284.605 602.820 284.810 ;
        RECT 591.190 282.330 592.680 282.895 ;
        RECT 601.930 282.860 602.270 284.605 ;
        RECT 601.900 282.330 602.300 282.860 ;
        RECT 591.190 281.870 602.300 282.330 ;
        RECT 591.190 281.860 602.280 281.870 ;
        RECT 591.190 281.605 592.680 281.860 ;
        RECT 631.590 281.830 631.920 289.755 ;
        RECT 631.550 281.610 631.920 281.830 ;
        RECT 157.220 278.220 158.320 278.855 ;
        RECT 158.800 278.220 160.190 278.830 ;
        RECT 157.220 277.540 160.190 278.220 ;
        RECT 157.220 277.015 158.320 277.540 ;
        RECT 158.800 276.930 160.190 277.540 ;
        RECT 591.770 270.660 592.180 281.605 ;
        RECT 631.550 280.860 631.910 281.610 ;
        RECT 631.550 280.760 631.920 280.860 ;
        RECT 631.590 271.655 631.920 280.760 ;
        RECT 632.730 278.655 633.080 296.185 ;
        RECT 641.630 290.825 642.110 291.195 ;
        RECT 641.710 289.175 642.030 290.825 ;
        RECT 641.600 289.100 642.130 289.175 ;
        RECT 648.410 289.160 649.540 289.170 ;
        RECT 648.410 289.120 651.600 289.160 ;
        RECT 657.090 289.150 657.860 306.280 ;
        RECT 652.060 289.120 657.860 289.150 ;
        RECT 648.410 289.100 657.860 289.120 ;
        RECT 641.600 288.790 657.860 289.100 ;
        RECT 641.600 288.780 649.540 288.790 ;
        RECT 641.600 288.695 642.130 288.780 ;
        RECT 648.410 288.760 649.540 288.780 ;
        RECT 652.060 288.600 657.860 288.790 ;
        RECT 652.060 288.570 657.470 288.600 ;
        RECT 632.510 277.685 633.380 278.655 ;
        RECT 631.500 271.520 632.020 271.655 ;
        RECT 591.750 270.045 592.180 270.660 ;
        RECT 631.430 271.165 632.020 271.520 ;
        RECT 591.250 268.955 592.620 270.045 ;
        RECT 601.430 266.125 602.510 266.515 ;
        RECT 591.050 264.140 592.560 264.685 ;
        RECT 601.710 264.140 602.190 266.125 ;
        RECT 591.050 263.770 602.200 264.140 ;
        RECT 591.050 263.565 592.560 263.770 ;
        RECT 591.420 255.760 592.060 263.565 ;
        RECT 591.390 255.150 592.060 255.760 ;
        RECT 591.390 251.625 592.000 255.150 ;
        RECT 631.430 253.975 631.870 271.165 ;
        RECT 632.730 260.885 633.080 277.685 ;
        RECT 641.550 272.355 642.030 272.725 ;
        RECT 641.630 270.705 641.950 272.355 ;
        RECT 659.970 270.840 660.760 311.070 ;
        RECT 668.180 311.050 668.720 311.070 ;
        RECT 666.180 307.805 667.590 309.305 ;
        RECT 641.520 270.700 642.050 270.705 ;
        RECT 641.520 270.690 648.450 270.700 ;
        RECT 649.000 270.690 660.850 270.840 ;
        RECT 641.520 270.340 660.850 270.690 ;
        RECT 641.520 270.225 642.050 270.340 ;
        RECT 648.330 270.320 660.850 270.340 ;
        RECT 649.000 270.060 660.850 270.320 ;
        RECT 659.970 269.930 660.760 270.060 ;
        RECT 632.340 260.135 633.580 260.885 ;
        RECT 641.400 254.625 641.880 254.995 ;
        RECT 631.310 253.505 631.980 253.975 ;
        RECT 591.190 250.135 592.240 251.625 ;
        RECT 631.340 234.750 631.740 253.505 ;
        RECT 641.480 252.990 641.800 254.625 ;
        RECT 666.590 253.080 667.160 307.805 ;
        RECT 794.420 305.900 795.990 306.285 ;
        RECT 794.420 305.030 796.020 305.900 ;
        RECT 794.420 305.005 795.990 305.030 ;
        RECT 849.070 298.640 849.620 298.660 ;
        RECT 785.430 298.500 786.190 298.570 ;
        RECT 843.880 298.500 849.650 298.640 ;
        RECT 694.890 296.955 695.390 297.485 ;
        RECT 712.420 296.995 712.850 297.815 ;
        RECT 694.950 294.570 695.310 296.955 ;
        RECT 694.950 292.590 695.330 294.570 ;
        RECT 694.970 290.555 695.330 292.590 ;
        RECT 712.430 291.465 712.800 296.995 ;
        RECT 730.030 296.975 730.420 297.775 ;
        RECT 747.700 297.025 748.190 297.955 ;
        RECT 785.350 297.930 849.650 298.500 ;
        RECT 730.110 292.625 730.420 296.975 ;
        RECT 729.910 291.925 731.090 292.625 ;
        RECT 694.720 288.525 696.210 290.555 ;
        RECT 711.900 290.005 713.680 291.465 ;
        RECT 726.740 287.360 728.290 287.555 ;
        RECT 747.750 287.360 748.180 297.025 ;
        RECT 726.740 286.750 748.200 287.360 ;
        RECT 779.390 286.810 781.310 287.235 ;
        RECT 726.740 286.740 747.220 286.750 ;
        RECT 726.740 286.475 728.290 286.740 ;
        RECT 774.600 286.320 781.310 286.810 ;
        RECT 745.780 269.900 746.190 270.045 ;
        RECT 721.610 269.815 746.190 269.900 ;
        RECT 686.620 269.440 687.080 269.585 ;
        RECT 711.040 269.440 711.500 269.565 ;
        RECT 686.620 269.080 711.500 269.440 ;
        RECT 686.620 268.735 687.080 269.080 ;
        RECT 711.040 268.715 711.500 269.080 ;
        RECT 721.400 269.490 746.190 269.815 ;
        RECT 721.400 268.885 721.970 269.490 ;
        RECT 745.780 269.095 746.190 269.490 ;
        RECT 703.810 268.300 704.340 268.655 ;
        RECT 728.590 268.300 729.120 268.805 ;
        RECT 703.810 267.920 729.120 268.300 ;
        RECT 738.610 268.570 739.060 268.635 ;
        RECT 763.620 268.570 764.070 268.965 ;
        RECT 738.610 268.255 764.070 268.570 ;
        RECT 738.610 268.180 763.830 268.255 ;
        RECT 738.610 267.925 739.060 268.180 ;
        RECT 703.810 267.745 704.340 267.920 ;
        RECT 728.590 267.895 729.120 267.920 ;
        RECT 692.980 262.540 693.920 262.605 ;
        RECT 774.640 262.540 775.130 286.320 ;
        RECT 779.390 285.725 781.310 286.320 ;
        RECT 785.430 285.320 786.190 297.930 ;
        RECT 843.880 297.920 849.650 297.930 ;
        RECT 849.070 292.555 849.620 297.920 ;
        RECT 848.990 291.755 849.920 292.555 ;
        RECT 868.130 291.665 869.240 292.285 ;
        RECT 785.420 284.920 786.190 285.320 ;
        RECT 832.890 285.275 834.320 286.315 ;
        RECT 777.630 271.070 778.240 271.080 ;
        RECT 777.630 271.025 784.540 271.070 ;
        RECT 777.630 270.690 785.000 271.025 ;
        RECT 692.980 262.030 775.220 262.540 ;
        RECT 692.980 261.695 693.920 262.030 ;
        RECT 776.110 257.430 777.040 257.725 ;
        RECT 710.770 257.020 777.040 257.430 ;
        RECT 649.410 253.040 667.720 253.080 ;
        RECT 648.590 252.990 667.720 253.040 ;
        RECT 641.480 252.975 667.720 252.990 ;
        RECT 641.370 252.600 667.720 252.975 ;
        RECT 710.770 252.925 711.240 257.020 ;
        RECT 776.110 256.785 777.040 257.020 ;
        RECT 641.370 252.495 641.900 252.600 ;
        RECT 648.590 252.580 667.720 252.600 ;
        RECT 649.410 252.390 667.720 252.580 ;
        RECT 710.280 252.145 711.240 252.925 ;
        RECT 745.760 248.370 746.170 248.515 ;
        RECT 721.590 248.285 746.170 248.370 ;
        RECT 686.600 247.910 687.060 248.055 ;
        RECT 711.020 247.910 711.480 248.035 ;
        RECT 686.600 247.550 711.480 247.910 ;
        RECT 686.600 247.205 687.060 247.550 ;
        RECT 711.020 247.185 711.480 247.550 ;
        RECT 721.380 247.960 746.170 248.285 ;
        RECT 721.380 247.355 721.950 247.960 ;
        RECT 745.760 247.565 746.170 247.960 ;
        RECT 703.790 246.770 704.320 247.125 ;
        RECT 728.570 246.770 729.100 247.275 ;
        RECT 703.790 246.390 729.100 246.770 ;
        RECT 738.590 247.040 739.040 247.105 ;
        RECT 763.600 247.040 764.050 247.435 ;
        RECT 738.590 246.725 764.050 247.040 ;
        RECT 738.590 246.650 763.810 246.725 ;
        RECT 738.590 246.395 739.040 246.650 ;
        RECT 703.790 246.215 704.320 246.390 ;
        RECT 728.570 246.365 729.100 246.390 ;
        RECT 777.630 246.290 778.240 270.690 ;
        RECT 784.130 270.395 785.000 270.690 ;
        RECT 784.150 263.040 785.000 263.165 ;
        RECT 785.420 263.040 786.100 284.920 ;
        RECT 801.990 280.535 803.020 281.575 ;
        RECT 817.970 281.050 818.700 281.455 ;
        RECT 865.170 281.175 866.030 282.185 ;
        RECT 817.950 280.855 818.700 281.050 ;
        RECT 836.960 281.020 837.920 281.030 ;
        RECT 836.740 280.980 841.370 281.020 ;
        RECT 836.740 280.965 841.390 280.980 ;
        RECT 817.950 278.320 818.270 280.855 ;
        RECT 827.960 280.225 828.520 280.795 ;
        RECT 836.550 280.720 841.390 280.965 ;
        RECT 836.550 280.515 837.140 280.720 ;
        RECT 840.940 280.685 841.390 280.720 ;
        RECT 827.970 278.320 828.300 280.225 ;
        RECT 836.580 279.360 836.900 280.515 ;
        RECT 840.940 280.215 841.470 280.685 ;
        RECT 841.780 279.805 842.480 280.395 ;
        RECT 841.830 278.790 842.280 279.805 ;
        RECT 841.130 278.725 842.280 278.790 ;
        RECT 840.630 278.500 842.280 278.725 ;
        RECT 840.630 278.490 842.160 278.500 ;
        RECT 836.580 278.320 836.900 278.340 ;
        RECT 798.000 278.295 837.300 278.320 ;
        RECT 797.390 278.270 837.300 278.295 ;
        RECT 797.390 278.020 837.310 278.270 ;
        RECT 840.630 278.195 841.330 278.490 ;
        RECT 797.390 277.415 798.610 278.020 ;
        RECT 837.000 276.520 837.310 278.020 ;
        RECT 840.790 276.520 841.140 278.195 ;
        RECT 837.000 276.190 841.140 276.520 ;
        RECT 837.000 276.180 841.020 276.190 ;
        RECT 837.000 274.075 837.310 276.180 ;
        RECT 836.970 273.415 837.500 274.075 ;
        RECT 802.920 270.830 803.910 270.995 ;
        RECT 865.460 270.830 865.760 281.175 ;
        RECT 802.920 270.530 865.760 270.830 ;
        RECT 802.920 270.475 803.910 270.530 ;
        RECT 797.560 269.130 798.520 269.365 ;
        RECT 833.130 269.130 834.240 269.590 ;
        RECT 797.560 268.830 837.400 269.130 ;
        RECT 797.560 268.375 798.520 268.830 ;
        RECT 833.130 268.440 834.240 268.830 ;
        RECT 837.000 267.845 837.380 268.830 ;
        RECT 836.850 267.375 837.420 267.845 ;
        RECT 821.600 266.790 822.640 267.215 ;
        RECT 837.010 266.810 837.730 267.045 ;
        RECT 835.820 266.790 837.730 266.810 ;
        RECT 821.600 266.515 837.730 266.790 ;
        RECT 821.600 266.490 837.310 266.515 ;
        RECT 821.600 266.225 822.640 266.490 ;
        RECT 868.630 263.530 869.020 291.665 ;
        RECT 803.110 263.495 869.100 263.530 ;
        RECT 784.150 262.680 786.100 263.040 ;
        RECT 802.540 262.960 869.100 263.495 ;
        RECT 802.540 262.845 803.730 262.960 ;
        RECT 868.630 262.930 869.020 262.960 ;
        RECT 784.150 262.660 785.880 262.680 ;
        RECT 784.150 262.525 785.000 262.660 ;
        RECT 852.680 254.605 853.510 255.465 ;
        RECT 866.290 252.895 867.330 253.735 ;
        RECT 866.610 246.290 867.030 252.895 ;
        RECT 777.630 245.320 867.040 246.290 ;
        RECT 630.890 233.320 632.270 234.750 ;
        RECT 389.560 229.090 393.870 229.995 ;
        RECT 406.300 229.090 409.730 230.950 ;
        RECT 389.560 227.040 409.730 229.090 ;
        RECT 389.560 226.425 393.870 227.040 ;
        RECT 406.300 226.350 409.730 227.040 ;
      LAYER via3 ;
        RECT 656.215 349.950 656.535 350.270 ;
        RECT 656.215 349.550 656.535 349.870 ;
        RECT 824.485 347.785 824.805 348.105 ;
        RECT 824.885 347.785 825.205 348.105 ;
        RECT 195.280 341.335 198.000 346.455 ;
        RECT 885.540 322.870 888.660 324.390 ;
        RECT 305.265 284.080 306.785 286.000 ;
        RECT 158.935 277.120 160.055 278.640 ;
        RECT 794.660 305.085 795.780 306.205 ;
        RECT 833.045 285.435 834.165 286.155 ;
        RECT 802.145 280.695 802.865 281.415 ;
        RECT 833.325 268.455 834.045 269.575 ;
        RECT 852.735 254.675 853.455 255.395 ;
        RECT 631.020 233.475 632.140 234.595 ;
        RECT 406.455 226.490 409.575 230.810 ;
      LAYER met4 ;
        RECT 656.055 349.800 656.695 350.295 ;
        RECT 656.055 349.630 825.180 349.800 ;
        RECT 656.055 349.525 825.190 349.630 ;
        RECT 656.330 349.470 825.190 349.525 ;
        RECT 824.780 348.185 825.190 349.470 ;
        RECT 824.405 347.705 825.285 348.185 ;
        RECT 195.165 346.120 198.115 346.545 ;
        RECT 160.730 343.770 198.115 346.120 ;
        RECT 160.810 333.490 162.580 343.770 ;
        RECT 195.165 341.245 198.115 343.770 ;
        RECT 171.410 333.500 181.300 337.320 ;
        RECT 163.670 333.490 181.300 333.500 ;
        RECT 160.600 333.480 181.300 333.490 ;
        RECT 160.490 331.290 181.300 333.480 ;
        RECT 160.490 312.540 162.700 331.290 ;
        RECT 163.670 331.250 181.300 331.290 ;
        RECT 171.410 328.230 181.300 331.250 ;
        RECT 885.385 322.735 888.815 324.525 ;
        RECT 307.790 315.160 313.290 315.390 ;
        RECT 307.790 315.150 313.330 315.160 ;
        RECT 319.370 315.150 329.260 318.970 ;
        RECT 160.470 312.480 162.990 312.540 ;
        RECT 160.470 310.550 163.010 312.480 ;
        RECT 160.470 310.500 165.360 310.550 ;
        RECT 171.410 310.500 181.300 314.320 ;
        RECT 307.790 312.900 329.260 315.150 ;
        RECT 307.790 312.840 313.330 312.900 ;
        RECT 307.790 312.780 313.290 312.840 ;
        RECT 307.970 310.590 309.840 312.780 ;
        RECT 160.470 308.250 181.300 310.500 ;
        RECT 160.470 308.130 165.360 308.250 ;
        RECT 160.470 291.540 162.990 308.130 ;
        RECT 171.410 305.230 181.300 308.250 ;
        RECT 308.020 308.120 309.790 310.590 ;
        RECT 319.370 309.880 329.260 312.900 ;
        RECT 308.020 292.460 309.860 308.120 ;
        RECT 412.420 306.790 414.220 306.840 ;
        RECT 412.420 306.780 795.000 306.790 ;
        RECT 412.420 306.265 795.160 306.780 ;
        RECT 412.420 306.090 795.945 306.265 ;
        RECT 319.370 292.460 329.260 295.970 ;
        RECT 160.470 288.090 163.050 291.540 ;
        RECT 160.470 287.510 162.990 288.090 ;
        RECT 160.470 287.500 165.370 287.510 ;
        RECT 171.410 287.500 181.300 291.320 ;
        RECT 160.470 285.250 181.300 287.500 ;
        RECT 308.020 289.760 329.260 292.460 ;
        RECT 412.420 291.120 414.220 306.090 ;
        RECT 794.465 305.905 795.945 306.090 ;
        RECT 794.465 305.025 795.975 305.905 ;
        RECT 412.420 290.750 414.380 291.120 ;
        RECT 308.020 289.160 309.860 289.760 ;
        RECT 311.580 289.700 329.260 289.760 ;
        RECT 308.020 286.470 309.930 289.160 ;
        RECT 319.370 286.880 329.260 289.700 ;
        RECT 160.470 285.190 165.370 285.250 ;
        RECT 158.845 278.120 160.145 278.835 ;
        RECT 160.470 278.120 162.990 285.190 ;
        RECT 171.410 282.230 181.300 285.250 ;
        RECT 305.185 285.650 306.865 286.185 ;
        RECT 308.020 285.650 309.860 286.470 ;
        RECT 305.185 284.640 309.860 285.650 ;
        RECT 305.185 283.895 306.865 284.640 ;
        RECT 158.845 277.470 162.990 278.120 ;
        RECT 158.845 276.925 160.145 277.470 ;
        RECT 160.470 269.230 162.990 277.470 ;
        RECT 160.470 267.030 163.030 269.230 ;
        RECT 308.020 269.120 309.860 284.640 ;
        RECT 311.420 269.150 313.130 269.180 ;
        RECT 319.370 269.150 329.260 272.970 ;
        RECT 311.420 269.120 329.260 269.150 ;
        RECT 160.470 264.590 162.990 267.030 ;
        RECT 160.470 264.500 165.390 264.590 ;
        RECT 171.410 264.500 181.300 268.320 ;
        RECT 307.790 266.900 329.260 269.120 ;
        RECT 307.790 266.790 313.660 266.900 ;
        RECT 160.470 262.270 181.300 264.500 ;
        RECT 319.370 263.880 329.260 266.900 ;
        RECT 160.470 245.250 162.990 262.270 ;
        RECT 164.400 262.250 181.300 262.270 ;
        RECT 171.410 259.230 181.300 262.250 ;
        RECT 412.520 252.170 414.380 290.750 ;
        RECT 832.935 285.295 834.275 286.295 ;
        RECT 802.035 280.555 802.975 281.555 ;
        RECT 802.160 275.540 802.790 280.555 ;
        RECT 802.160 260.140 802.820 275.540 ;
        RECT 833.330 269.595 833.750 285.295 ;
        RECT 833.175 268.435 834.195 269.595 ;
        RECT 422.810 252.290 432.700 255.800 ;
        RECT 802.190 255.380 802.820 260.140 ;
        RECT 852.725 255.380 853.465 255.445 ;
        RECT 802.190 254.650 853.465 255.380 ;
        RECT 852.725 254.625 853.465 254.650 ;
        RECT 415.280 252.170 432.700 252.290 ;
        RECT 412.510 250.150 432.700 252.170 ;
        RECT 412.310 249.530 432.700 250.150 ;
        RECT 412.310 249.470 417.910 249.530 ;
        RECT 412.310 247.430 414.680 249.470 ;
        RECT 160.470 241.530 162.970 245.250 ;
        RECT 160.470 241.500 165.170 241.530 ;
        RECT 171.410 241.500 181.300 245.320 ;
        RECT 412.310 241.880 414.540 247.430 ;
        RECT 422.810 246.710 432.700 249.530 ;
        RECT 160.470 239.250 181.300 241.500 ;
        RECT 160.470 239.210 165.170 239.250 ;
        RECT 160.470 239.060 162.970 239.210 ;
        RECT 160.470 239.040 162.790 239.060 ;
        RECT 171.410 236.230 181.300 239.250 ;
        RECT 412.230 237.980 414.540 241.880 ;
        RECT 406.345 230.460 409.685 230.955 ;
        RECT 412.310 230.460 414.540 237.980 ;
        RECT 620.750 234.130 630.530 234.160 ;
        RECT 557.960 234.120 630.530 234.130 ;
        RECT 630.935 234.120 632.225 234.755 ;
        RECT 730.870 234.410 758.320 234.630 ;
        RECT 837.040 234.510 864.490 234.950 ;
        RECT 886.840 234.530 888.110 322.735 ;
        RECT 883.900 234.510 929.540 234.530 ;
        RECT 837.040 234.430 929.540 234.510 ;
        RECT 775.210 234.410 929.540 234.430 ;
        RECT 633.440 234.120 648.200 234.160 ;
        RECT 557.960 234.110 648.200 234.120 ;
        RECT 557.890 234.070 648.200 234.110 ;
        RECT 730.870 234.090 929.540 234.410 ;
        RECT 665.920 234.070 929.540 234.090 ;
        RECT 406.345 229.160 414.540 230.460 ;
        RECT 406.345 228.980 418.680 229.160 ;
        RECT 422.810 228.980 432.700 232.800 ;
        RECT 557.890 232.300 929.540 234.070 ;
        RECT 557.890 232.200 865.290 232.300 ;
        RECT 557.890 231.900 758.320 232.200 ;
        RECT 775.210 232.110 865.290 232.200 ;
        RECT 775.210 231.910 843.060 232.110 ;
        RECT 557.960 231.860 758.320 231.900 ;
        RECT 557.960 231.610 648.200 231.860 ;
        RECT 558.020 230.360 560.590 231.610 ;
        RECT 406.345 228.210 432.700 228.980 ;
        RECT 406.345 226.345 409.685 228.210 ;
        RECT 412.310 226.730 432.700 228.210 ;
        RECT 412.310 226.460 418.680 226.730 ;
        RECT 412.310 225.720 414.680 226.460 ;
        RECT 422.810 223.710 432.700 226.730 ;
        RECT 558.120 217.990 560.590 230.360 ;
        RECT 579.680 217.990 582.150 231.610 ;
        RECT 601.030 217.990 603.500 231.610 ;
        RECT 620.750 231.320 648.200 231.610 ;
        RECT 665.920 231.790 758.320 231.860 ;
        RECT 665.920 231.570 733.210 231.790 ;
        RECT 622.600 217.990 625.070 231.320 ;
        RECT 630.120 231.250 634.450 231.320 ;
        RECT 644.970 230.360 647.530 231.320 ;
        RECT 665.980 230.360 668.540 231.570 ;
        RECT 645.060 217.990 647.530 230.360 ;
        RECT 666.070 217.990 668.540 230.360 ;
        RECT 687.750 217.990 690.220 231.570 ;
        RECT 709.230 230.360 711.790 231.570 ;
        RECT 709.320 217.990 711.790 230.360 ;
        RECT 730.660 217.990 733.130 231.570 ;
        RECT 754.260 230.360 756.830 231.790 ;
        RECT 775.270 230.360 777.840 231.910 ;
        RECT 797.060 231.460 799.260 231.910 ;
        RECT 817.180 231.650 822.740 231.910 ;
        RECT 839.960 231.710 843.060 231.910 ;
        RECT 797.060 230.360 799.500 231.460 ;
        RECT 754.360 217.990 756.830 230.360 ;
        RECT 775.370 217.990 777.840 230.360 ;
        RECT 797.160 218.080 799.500 230.360 ;
        RECT 818.510 218.080 820.850 231.650 ;
        RECT 839.960 218.080 842.300 231.710 ;
        RECT 862.950 218.080 865.290 232.110 ;
        RECT 883.850 232.010 929.540 232.300 ;
        RECT 883.850 218.080 886.190 232.010 ;
        RECT 905.750 230.360 908.130 232.010 ;
        RECT 927.210 231.530 929.540 232.010 ;
        RECT 927.210 230.360 929.590 231.530 ;
        RECT 905.790 218.080 908.130 230.360 ;
        RECT 927.250 218.080 929.590 230.360 ;
        RECT 558.120 212.470 780.840 217.990 ;
        RECT 792.340 217.440 1013.240 218.080 ;
        RECT 558.980 201.030 780.840 212.470 ;
        RECT 791.380 201.120 1013.240 217.440 ;
        RECT 558.980 189.990 573.060 201.030 ;
        RECT 791.380 190.080 805.460 201.120 ;
        RECT 558.980 173.030 780.840 189.990 ;
        RECT 791.380 173.120 1013.240 190.080 ;
        RECT 558.980 161.990 573.060 173.030 ;
        RECT 791.380 162.080 805.460 173.120 ;
        RECT 558.980 161.650 780.840 161.990 ;
        RECT 791.380 161.650 1013.240 162.080 ;
        RECT 558.980 145.120 1013.240 161.650 ;
        RECT 558.980 145.030 805.460 145.120 ;
        RECT 558.980 133.990 573.060 145.030 ;
        RECT 766.580 144.690 805.460 145.030 ;
        RECT 791.380 134.080 805.460 144.690 ;
        RECT 558.980 117.030 780.840 133.990 ;
        RECT 791.380 117.120 1013.240 134.080 ;
        RECT 558.980 107.310 573.060 117.030 ;
        RECT 791.380 107.400 805.460 117.120 ;
        RECT 554.820 105.990 578.600 107.310 ;
        RECT 787.920 106.080 811.000 107.400 ;
        RECT 554.820 89.030 780.840 105.990 ;
        RECT 787.920 89.120 1013.240 106.080 ;
        RECT 554.820 87.190 578.600 89.030 ;
        RECT 787.920 87.280 811.000 89.120 ;
  END
END LVDT
END LIBRARY

