// File goldcode.vhd translated with vhd2vl v2.4 VHDL to Verilog RTL translator
// vhd2vl settings:
//  * Verilog Module Declaration Style: 1995

// vhd2vl is Free (libre) Software:
//   Copyright (C) 2001 Vincenzo Liguori - Ocean Logic Pty Ltd
//     http://www.ocean-logic.com
//   Modifications Copyright (C) 2006 Mark Gonzales - PMC Sierra Inc
//   Modifications (C) 2010 Shankar Giri
//   Modifications Copyright (C) 2002, 2005, 2008-2010 Larry Doolittle - LBNL
//     http://doolittle.icarus.com/~larry/vhd2vl/
//
//   vhd2vl comes with ABSOLUTELY NO WARRANTY.  Always check the resulting
//   Verilog for correctness, ideally with a formal verification tool.
//
//   You are welcome to redistribute vhd2vl under certain conditions.
//   See the license (GPLv2) file included with the source for details.

// The result of translation follows.  Its copyright status should be
// considered unchanged from the original VHDL.

//FILE NAME : goldcode.vhd
//----**********************************************************************
// DESCRIPTION 
//    Gold code is generated by g1 code and g2 code.
//**************************************************************************
//   I/O signals
//   reset    -- used to set the register contents of g1 reg and g2 reg.
//   clk      -- provided by the codectrllogic to generate goldcode.
//   goldcode -- output of the gold code.  	  
//**************************************************************************
// no timescale needed
`timescale 1ns / 1ps
module goldcode(
reset,
clk,
car_change,
epochrx,
code_sel,
goldcode,
gold1,
gold2,
irnss_sel,
irnss_code
);

input reset, clk;
input car_change;
output epochrx;
input [4:0] code_sel;
output goldcode, gold1, gold2;
input irnss_sel;
input [10:1] irnss_code;

wire reset;
wire clk;
wire car_change;
reg epochrx;
wire [4:0] code_sel;
reg goldcode;
reg gold1;
reg gold2;


reg [10:1] g1codereg;
reg [10:1] g2codereg;
reg g1out;
reg g2out;

  always @(negedge reset or posedge clk or posedge car_change) begin
    if(reset == 1'b 0) begin
      g1codereg <= 10'b 1111111111;
    end 
    else if(car_change == 1'b 1) begin
      g1codereg <= 10'b 1111111111;
    end
    else begin
      g1codereg[1] <= g1codereg[3] ^ g1codereg[10];
      g1codereg[10:2] <= g1codereg[9:1];
    end
  end

  always @(negedge clk) begin
    if(g1codereg == 10'b 1111111111) begin
      epochrx <= 1'b 1;
    end
    else begin
      epochrx <= 1'b 0;
    end
  end
  wire [10:1] code_wire;
  assign code_wire = irnss_sel==1'b0 ? 10'b 1111111111 : irnss_code;

  always @(negedge reset or posedge clk or posedge car_change) begin
    if(reset == 1'b 0) begin
      g2codereg <= code_wire;
    end 
    else if(car_change == 1'b 1) begin
      g2codereg <= code_wire;
    end 
    else begin
      g2codereg[1] <= g2codereg[2] ^ g2codereg[3] ^ g2codereg[6] ^ g2codereg[8] ^ g2codereg[9] ^ g2codereg[10];
      g2codereg[10:2] <= g2codereg[9:1];
    end
  end

  always @(reset or g2codereg or code_sel or g1out or g2out or g1codereg) begin
    if(reset == 1'b 0) begin
      g2out <= 1'b 0;
      g1out <= 1'b 0;
      goldcode <= 1'b 0;
    end
    else begin
      // goldcode<='1';
      if(irnss_sel == 1'b0) begin
        case(code_sel)
        5'b 00001 : begin
          g2out <= g2codereg[2] ^ g2codereg[6];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 00010 : begin
          g2out <= g2codereg[3] ^ g2codereg[7];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 00011 : begin
          g2out <= g2codereg[4] ^ g2codereg[8];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 00100 : begin
          g2out <= g2codereg[5] ^ g2codereg[9];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 00101 : begin
          g2out <= g2codereg[1] ^ g2codereg[9];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 00110 : begin
          g2out <= g2codereg[2] ^ g2codereg[10];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 00111 : begin
          g2out <= g2codereg[1] ^ g2codereg[8];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 01000 : begin
          g2out <= g2codereg[2] ^ g2codereg[9];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 01001 : begin
          g2out <= g2codereg[3] ^ g2codereg[10];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 01010 : begin
          g2out <= g2codereg[2] ^ g2codereg[3];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 01011 : begin
          g2out <= g2codereg[3] ^ g2codereg[4];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 01100 : begin
          g2out <= g2codereg[5] ^ g2codereg[6];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 01101 : begin
          g2out <= g2codereg[6] ^ g2codereg[7];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 01110 : begin
          g2out <= g2codereg[7] ^ g2codereg[8];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 01111 : begin
          g2out <= g2codereg[8] ^ g2codereg[9];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 10000 : begin
          g2out <= g2codereg[9] ^ g2codereg[10];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 10001 : begin
          g2out <= g2codereg[1] ^ g2codereg[4];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 10010 : begin
          g2out <= g2codereg[2] ^ g2codereg[5];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 10011 : begin
          g2out <= g2codereg[3] ^ g2codereg[6];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 10100 : begin
          g2out <= g2codereg[4] ^ g2codereg[7];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 10101 : begin
          g2out <= g2codereg[5] ^ g2codereg[8];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 10110 : begin
          g2out <= g2codereg[6] ^ g2codereg[9];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 10111 : begin
          g2out <= g2codereg[1] ^ g2codereg[3];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 11000 : begin
          g2out <= g2codereg[4] ^ g2codereg[6];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 11001 : begin
          g2out <= g2codereg[5] ^ g2codereg[7];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 11010 : begin
          g2out <= g2codereg[6] ^ g2codereg[8];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 11011 : begin
          g2out <= g2codereg[7] ^ g2codereg[9];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 11100 : begin
          g2out <= g2codereg[8] ^ g2codereg[10];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 11101 : begin
          g2out <= g2codereg[1] ^ g2codereg[6];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 11110 : begin
          g2out <= g2codereg[1] ^ g2codereg[7];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 11111 : begin
          g2out <= g2codereg[3] ^ g2codereg[8];
          g1out <= g1codereg[10];
          goldcode <= g1out ^ g2out;
        end
        5'b 00000 : begin
          g2out <= g2codereg[4] ^ g2codereg[9];
          g1out <= g1codereg[10];
          goldcode <= 1'b 1;
        end
        default : begin
          g2out <= 1'b 1;
          //edited intially commented originally '0'
        end
        endcase
      end else begin
        g1out <= g1codereg[10];
        g2out <= g2codereg[10];
        goldcode <= g1out ^ g2out;
      end
      gold1 <= g1out;
      gold2 <= g2out;
    end
  end

    //  g1out    <= g1codereg(10);
  //	g2out    <= g2codereg(5) xor g2codereg(7);
  //	goldcode <= g1out xor g2out;

endmodule
