VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_macro
  CLASS BLOCK ;
  FOREIGN analog_macro ;
  ORIGIN 37.770 44.270 ;
  SIZE 824.770 BY 440.310 ;
  PIN vinit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    ANTENNADIFFAREA 31.900000 ;
    PORT
      LAYER li1 ;
        RECT 688.970 244.190 689.140 249.230 ;
        RECT 691.550 244.190 691.720 249.230 ;
        RECT 694.130 244.190 694.300 249.230 ;
        RECT 696.710 244.190 696.880 249.230 ;
        RECT 699.290 244.190 699.460 249.230 ;
        RECT 701.870 244.190 702.040 249.230 ;
        RECT 704.450 244.190 704.620 249.230 ;
        RECT 707.030 244.190 707.200 249.230 ;
        RECT 709.610 244.190 709.780 249.230 ;
        RECT 712.190 244.190 712.360 249.230 ;
        RECT 714.770 244.190 714.940 249.230 ;
        RECT 739.770 244.360 739.940 249.400 ;
        RECT 742.350 244.360 742.520 249.400 ;
        RECT 744.930 244.360 745.100 249.400 ;
        RECT 747.510 244.360 747.680 249.400 ;
        RECT 750.090 244.360 750.260 249.400 ;
        RECT 752.670 244.360 752.840 249.400 ;
        RECT 755.250 244.360 755.420 249.400 ;
        RECT 757.830 244.360 758.000 249.400 ;
        RECT 760.410 244.360 760.580 249.400 ;
        RECT 762.990 244.360 763.160 249.400 ;
        RECT 765.570 244.360 765.740 249.400 ;
        RECT 132.530 109.675 133.610 109.845 ;
      LAYER mcon ;
        RECT 688.970 244.270 689.140 249.150 ;
        RECT 691.550 244.270 691.720 249.150 ;
        RECT 694.130 244.270 694.300 249.150 ;
        RECT 696.710 244.270 696.880 249.150 ;
        RECT 699.290 244.270 699.460 249.150 ;
        RECT 701.870 244.270 702.040 249.150 ;
        RECT 704.450 244.270 704.620 249.150 ;
        RECT 707.030 244.270 707.200 249.150 ;
        RECT 709.610 244.270 709.780 249.150 ;
        RECT 712.190 244.270 712.360 249.150 ;
        RECT 714.770 244.270 714.940 249.150 ;
        RECT 739.770 244.440 739.940 249.320 ;
        RECT 742.350 244.440 742.520 249.320 ;
        RECT 744.930 244.440 745.100 249.320 ;
        RECT 747.510 244.440 747.680 249.320 ;
        RECT 750.090 244.440 750.260 249.320 ;
        RECT 752.670 244.440 752.840 249.320 ;
        RECT 755.250 244.440 755.420 249.320 ;
        RECT 757.830 244.440 758.000 249.320 ;
        RECT 760.410 244.440 760.580 249.320 ;
        RECT 762.990 244.440 763.160 249.320 ;
        RECT 765.570 244.440 765.740 249.320 ;
        RECT 132.610 109.675 133.530 109.845 ;
      LAYER met1 ;
        RECT 688.940 243.585 689.170 249.210 ;
        RECT 691.520 243.585 691.750 249.210 ;
        RECT 694.100 243.585 694.330 249.210 ;
        RECT 696.680 243.585 696.910 249.210 ;
        RECT 699.260 243.585 699.490 249.210 ;
        RECT 701.840 243.585 702.070 249.210 ;
        RECT 704.420 243.585 704.650 249.210 ;
        RECT 707.000 243.585 707.230 249.210 ;
        RECT 709.580 243.585 709.810 249.210 ;
        RECT 712.160 243.585 712.390 249.210 ;
        RECT 714.740 243.585 714.970 249.210 ;
        RECT 739.740 243.660 739.970 249.380 ;
        RECT 742.320 243.660 742.550 249.380 ;
        RECT 744.900 243.660 745.130 249.380 ;
        RECT 747.480 243.660 747.710 249.380 ;
        RECT 750.060 243.660 750.290 249.380 ;
        RECT 752.640 243.660 752.870 249.380 ;
        RECT 755.220 243.660 755.450 249.380 ;
        RECT 757.800 243.660 758.030 249.380 ;
        RECT 760.380 243.660 760.610 249.380 ;
        RECT 762.960 243.660 763.190 249.380 ;
        RECT 765.540 243.660 765.770 249.380 ;
        RECT 688.220 242.210 715.690 243.585 ;
        RECT 739.020 242.285 766.490 243.660 ;
        RECT 131.600 108.130 140.380 109.960 ;
      LAYER via ;
        RECT 688.730 243.005 689.030 243.305 ;
        RECT 689.330 243.005 689.630 243.305 ;
        RECT 689.930 243.005 690.230 243.305 ;
        RECT 690.530 243.005 690.830 243.305 ;
        RECT 691.130 243.005 691.430 243.305 ;
        RECT 691.730 243.005 692.030 243.305 ;
        RECT 692.330 243.005 692.630 243.305 ;
        RECT 692.930 243.005 693.230 243.305 ;
        RECT 693.530 243.005 693.830 243.305 ;
        RECT 694.130 243.005 694.430 243.305 ;
        RECT 694.730 243.005 695.030 243.305 ;
        RECT 695.330 243.005 695.630 243.305 ;
        RECT 695.930 243.005 696.230 243.305 ;
        RECT 696.530 243.005 696.830 243.305 ;
        RECT 697.130 243.005 697.430 243.305 ;
        RECT 697.730 243.005 698.030 243.305 ;
        RECT 698.330 243.005 698.630 243.305 ;
        RECT 698.930 243.005 699.230 243.305 ;
        RECT 699.530 243.005 699.830 243.305 ;
        RECT 700.130 243.005 700.430 243.305 ;
        RECT 700.730 243.005 701.030 243.305 ;
        RECT 701.330 243.005 701.630 243.305 ;
        RECT 701.930 243.005 702.230 243.305 ;
        RECT 702.530 243.005 702.830 243.305 ;
        RECT 703.130 243.005 703.430 243.305 ;
        RECT 703.730 243.005 704.030 243.305 ;
        RECT 704.330 243.005 704.630 243.305 ;
        RECT 704.930 243.005 705.230 243.305 ;
        RECT 705.530 243.005 705.830 243.305 ;
        RECT 706.130 243.005 706.430 243.305 ;
        RECT 706.730 243.005 707.030 243.305 ;
        RECT 707.330 243.005 707.630 243.305 ;
        RECT 707.930 243.005 708.230 243.305 ;
        RECT 708.530 243.005 708.830 243.305 ;
        RECT 709.130 243.005 709.430 243.305 ;
        RECT 709.730 243.005 710.030 243.305 ;
        RECT 710.330 243.005 710.630 243.305 ;
        RECT 710.930 243.005 711.230 243.305 ;
        RECT 711.530 243.005 711.830 243.305 ;
        RECT 712.130 243.005 712.430 243.305 ;
        RECT 712.730 243.005 713.030 243.305 ;
        RECT 713.330 243.005 713.630 243.305 ;
        RECT 713.930 243.005 714.230 243.305 ;
        RECT 714.530 243.005 714.830 243.305 ;
        RECT 715.130 243.005 715.430 243.305 ;
        RECT 688.730 242.405 689.030 242.705 ;
        RECT 689.330 242.405 689.630 242.705 ;
        RECT 689.930 242.405 690.230 242.705 ;
        RECT 690.530 242.405 690.830 242.705 ;
        RECT 691.130 242.405 691.430 242.705 ;
        RECT 691.730 242.405 692.030 242.705 ;
        RECT 692.330 242.405 692.630 242.705 ;
        RECT 692.930 242.405 693.230 242.705 ;
        RECT 693.530 242.405 693.830 242.705 ;
        RECT 694.130 242.405 694.430 242.705 ;
        RECT 694.730 242.405 695.030 242.705 ;
        RECT 695.330 242.405 695.630 242.705 ;
        RECT 695.930 242.405 696.230 242.705 ;
        RECT 696.530 242.405 696.830 242.705 ;
        RECT 697.130 242.405 697.430 242.705 ;
        RECT 697.730 242.405 698.030 242.705 ;
        RECT 698.330 242.405 698.630 242.705 ;
        RECT 698.930 242.405 699.230 242.705 ;
        RECT 699.530 242.405 699.830 242.705 ;
        RECT 700.130 242.405 700.430 242.705 ;
        RECT 700.730 242.405 701.030 242.705 ;
        RECT 701.330 242.405 701.630 242.705 ;
        RECT 701.930 242.405 702.230 242.705 ;
        RECT 702.530 242.405 702.830 242.705 ;
        RECT 703.130 242.405 703.430 242.705 ;
        RECT 703.730 242.405 704.030 242.705 ;
        RECT 704.330 242.405 704.630 242.705 ;
        RECT 704.930 242.405 705.230 242.705 ;
        RECT 705.530 242.405 705.830 242.705 ;
        RECT 706.130 242.405 706.430 242.705 ;
        RECT 706.730 242.405 707.030 242.705 ;
        RECT 707.330 242.405 707.630 242.705 ;
        RECT 707.930 242.405 708.230 242.705 ;
        RECT 708.530 242.405 708.830 242.705 ;
        RECT 709.130 242.405 709.430 242.705 ;
        RECT 709.730 242.405 710.030 242.705 ;
        RECT 710.330 242.405 710.630 242.705 ;
        RECT 710.930 242.405 711.230 242.705 ;
        RECT 711.530 242.405 711.830 242.705 ;
        RECT 712.130 242.405 712.430 242.705 ;
        RECT 712.730 242.405 713.030 242.705 ;
        RECT 713.330 242.405 713.630 242.705 ;
        RECT 713.930 242.405 714.230 242.705 ;
        RECT 714.530 242.405 714.830 242.705 ;
        RECT 715.130 242.405 715.430 242.705 ;
        RECT 739.280 243.080 739.580 243.380 ;
        RECT 739.880 243.080 740.180 243.380 ;
        RECT 740.480 243.080 740.780 243.380 ;
        RECT 741.080 243.080 741.380 243.380 ;
        RECT 741.680 243.080 741.980 243.380 ;
        RECT 742.280 243.080 742.580 243.380 ;
        RECT 742.880 243.080 743.180 243.380 ;
        RECT 743.480 243.080 743.780 243.380 ;
        RECT 744.080 243.080 744.380 243.380 ;
        RECT 744.680 243.080 744.980 243.380 ;
        RECT 745.280 243.080 745.580 243.380 ;
        RECT 745.880 243.080 746.180 243.380 ;
        RECT 746.480 243.080 746.780 243.380 ;
        RECT 747.080 243.080 747.380 243.380 ;
        RECT 747.680 243.080 747.980 243.380 ;
        RECT 748.280 243.080 748.580 243.380 ;
        RECT 748.880 243.080 749.180 243.380 ;
        RECT 749.480 243.080 749.780 243.380 ;
        RECT 750.080 243.080 750.380 243.380 ;
        RECT 750.680 243.080 750.980 243.380 ;
        RECT 751.280 243.080 751.580 243.380 ;
        RECT 751.880 243.080 752.180 243.380 ;
        RECT 752.480 243.080 752.780 243.380 ;
        RECT 753.080 243.080 753.380 243.380 ;
        RECT 753.680 243.080 753.980 243.380 ;
        RECT 754.280 243.080 754.580 243.380 ;
        RECT 754.880 243.080 755.180 243.380 ;
        RECT 755.480 243.080 755.780 243.380 ;
        RECT 756.080 243.080 756.380 243.380 ;
        RECT 756.680 243.080 756.980 243.380 ;
        RECT 757.280 243.080 757.580 243.380 ;
        RECT 757.880 243.080 758.180 243.380 ;
        RECT 758.480 243.080 758.780 243.380 ;
        RECT 759.080 243.080 759.380 243.380 ;
        RECT 759.680 243.080 759.980 243.380 ;
        RECT 760.280 243.080 760.580 243.380 ;
        RECT 760.880 243.080 761.180 243.380 ;
        RECT 761.480 243.080 761.780 243.380 ;
        RECT 762.080 243.080 762.380 243.380 ;
        RECT 762.680 243.080 762.980 243.380 ;
        RECT 763.280 243.080 763.580 243.380 ;
        RECT 763.880 243.080 764.180 243.380 ;
        RECT 764.480 243.080 764.780 243.380 ;
        RECT 765.080 243.080 765.380 243.380 ;
        RECT 765.680 243.080 765.980 243.380 ;
        RECT 739.280 242.480 739.580 242.780 ;
        RECT 739.880 242.480 740.180 242.780 ;
        RECT 740.480 242.480 740.780 242.780 ;
        RECT 741.080 242.480 741.380 242.780 ;
        RECT 741.680 242.480 741.980 242.780 ;
        RECT 742.280 242.480 742.580 242.780 ;
        RECT 742.880 242.480 743.180 242.780 ;
        RECT 743.480 242.480 743.780 242.780 ;
        RECT 744.080 242.480 744.380 242.780 ;
        RECT 744.680 242.480 744.980 242.780 ;
        RECT 745.280 242.480 745.580 242.780 ;
        RECT 745.880 242.480 746.180 242.780 ;
        RECT 746.480 242.480 746.780 242.780 ;
        RECT 747.080 242.480 747.380 242.780 ;
        RECT 747.680 242.480 747.980 242.780 ;
        RECT 748.280 242.480 748.580 242.780 ;
        RECT 748.880 242.480 749.180 242.780 ;
        RECT 749.480 242.480 749.780 242.780 ;
        RECT 750.080 242.480 750.380 242.780 ;
        RECT 750.680 242.480 750.980 242.780 ;
        RECT 751.280 242.480 751.580 242.780 ;
        RECT 751.880 242.480 752.180 242.780 ;
        RECT 752.480 242.480 752.780 242.780 ;
        RECT 753.080 242.480 753.380 242.780 ;
        RECT 753.680 242.480 753.980 242.780 ;
        RECT 754.280 242.480 754.580 242.780 ;
        RECT 754.880 242.480 755.180 242.780 ;
        RECT 755.480 242.480 755.780 242.780 ;
        RECT 756.080 242.480 756.380 242.780 ;
        RECT 756.680 242.480 756.980 242.780 ;
        RECT 757.280 242.480 757.580 242.780 ;
        RECT 757.880 242.480 758.180 242.780 ;
        RECT 758.480 242.480 758.780 242.780 ;
        RECT 759.080 242.480 759.380 242.780 ;
        RECT 759.680 242.480 759.980 242.780 ;
        RECT 760.280 242.480 760.580 242.780 ;
        RECT 760.880 242.480 761.180 242.780 ;
        RECT 761.480 242.480 761.780 242.780 ;
        RECT 762.080 242.480 762.380 242.780 ;
        RECT 762.680 242.480 762.980 242.780 ;
        RECT 763.280 242.480 763.580 242.780 ;
        RECT 763.880 242.480 764.180 242.780 ;
        RECT 764.480 242.480 764.780 242.780 ;
        RECT 765.080 242.480 765.380 242.780 ;
        RECT 765.680 242.480 765.980 242.780 ;
        RECT 139.570 108.630 140.070 109.490 ;
      LAYER met2 ;
        RECT 335.050 234.320 354.880 250.370 ;
        RECT 688.130 242.105 715.730 243.605 ;
        RECT 738.980 242.180 766.580 243.680 ;
        RECT 339.640 149.930 344.830 234.320 ;
        RECT 242.250 147.890 344.830 149.930 ;
        RECT 241.900 145.060 344.830 147.890 ;
        RECT 241.900 144.750 341.840 145.060 ;
        RECT 241.900 120.430 245.710 144.750 ;
        RECT 226.540 117.450 229.280 119.020 ;
        RECT 152.850 117.410 229.280 117.450 ;
        RECT 152.820 116.160 229.280 117.410 ;
        RECT 139.150 109.660 140.410 109.950 ;
        RECT 152.820 109.660 154.500 116.160 ;
        RECT 226.540 115.180 229.280 116.160 ;
        RECT 139.150 108.380 154.500 109.660 ;
        RECT 139.150 108.275 153.970 108.380 ;
        RECT 139.150 108.260 147.150 108.275 ;
        RECT 139.150 108.100 140.410 108.260 ;
      LAYER via2 ;
        RECT 340.710 236.840 349.210 242.820 ;
        RECT 688.730 243.005 689.030 243.305 ;
        RECT 689.330 243.005 689.630 243.305 ;
        RECT 689.930 243.005 690.230 243.305 ;
        RECT 690.530 243.005 690.830 243.305 ;
        RECT 691.130 243.005 691.430 243.305 ;
        RECT 691.730 243.005 692.030 243.305 ;
        RECT 692.330 243.005 692.630 243.305 ;
        RECT 692.930 243.005 693.230 243.305 ;
        RECT 693.530 243.005 693.830 243.305 ;
        RECT 694.130 243.005 694.430 243.305 ;
        RECT 694.730 243.005 695.030 243.305 ;
        RECT 695.330 243.005 695.630 243.305 ;
        RECT 695.930 243.005 696.230 243.305 ;
        RECT 696.530 243.005 696.830 243.305 ;
        RECT 697.130 243.005 697.430 243.305 ;
        RECT 697.730 243.005 698.030 243.305 ;
        RECT 698.330 243.005 698.630 243.305 ;
        RECT 698.930 243.005 699.230 243.305 ;
        RECT 699.530 243.005 699.830 243.305 ;
        RECT 700.130 243.005 700.430 243.305 ;
        RECT 700.730 243.005 701.030 243.305 ;
        RECT 701.330 243.005 701.630 243.305 ;
        RECT 701.930 243.005 702.230 243.305 ;
        RECT 702.530 243.005 702.830 243.305 ;
        RECT 703.130 243.005 703.430 243.305 ;
        RECT 703.730 243.005 704.030 243.305 ;
        RECT 704.330 243.005 704.630 243.305 ;
        RECT 704.930 243.005 705.230 243.305 ;
        RECT 705.530 243.005 705.830 243.305 ;
        RECT 706.130 243.005 706.430 243.305 ;
        RECT 706.730 243.005 707.030 243.305 ;
        RECT 707.330 243.005 707.630 243.305 ;
        RECT 707.930 243.005 708.230 243.305 ;
        RECT 708.530 243.005 708.830 243.305 ;
        RECT 709.130 243.005 709.430 243.305 ;
        RECT 709.730 243.005 710.030 243.305 ;
        RECT 710.330 243.005 710.630 243.305 ;
        RECT 710.930 243.005 711.230 243.305 ;
        RECT 711.530 243.005 711.830 243.305 ;
        RECT 712.130 243.005 712.430 243.305 ;
        RECT 712.730 243.005 713.030 243.305 ;
        RECT 713.330 243.005 713.630 243.305 ;
        RECT 713.930 243.005 714.230 243.305 ;
        RECT 714.530 243.005 714.830 243.305 ;
        RECT 715.130 243.005 715.430 243.305 ;
        RECT 688.730 242.405 689.030 242.705 ;
        RECT 689.330 242.405 689.630 242.705 ;
        RECT 689.930 242.405 690.230 242.705 ;
        RECT 690.530 242.405 690.830 242.705 ;
        RECT 691.130 242.405 691.430 242.705 ;
        RECT 691.730 242.405 692.030 242.705 ;
        RECT 692.330 242.405 692.630 242.705 ;
        RECT 692.930 242.405 693.230 242.705 ;
        RECT 693.530 242.405 693.830 242.705 ;
        RECT 694.130 242.405 694.430 242.705 ;
        RECT 694.730 242.405 695.030 242.705 ;
        RECT 695.330 242.405 695.630 242.705 ;
        RECT 695.930 242.405 696.230 242.705 ;
        RECT 696.530 242.405 696.830 242.705 ;
        RECT 697.130 242.405 697.430 242.705 ;
        RECT 697.730 242.405 698.030 242.705 ;
        RECT 698.330 242.405 698.630 242.705 ;
        RECT 698.930 242.405 699.230 242.705 ;
        RECT 699.530 242.405 699.830 242.705 ;
        RECT 700.130 242.405 700.430 242.705 ;
        RECT 700.730 242.405 701.030 242.705 ;
        RECT 701.330 242.405 701.630 242.705 ;
        RECT 701.930 242.405 702.230 242.705 ;
        RECT 702.530 242.405 702.830 242.705 ;
        RECT 703.130 242.405 703.430 242.705 ;
        RECT 703.730 242.405 704.030 242.705 ;
        RECT 704.330 242.405 704.630 242.705 ;
        RECT 704.930 242.405 705.230 242.705 ;
        RECT 705.530 242.405 705.830 242.705 ;
        RECT 706.130 242.405 706.430 242.705 ;
        RECT 706.730 242.405 707.030 242.705 ;
        RECT 707.330 242.405 707.630 242.705 ;
        RECT 707.930 242.405 708.230 242.705 ;
        RECT 708.530 242.405 708.830 242.705 ;
        RECT 709.130 242.405 709.430 242.705 ;
        RECT 709.730 242.405 710.030 242.705 ;
        RECT 710.330 242.405 710.630 242.705 ;
        RECT 710.930 242.405 711.230 242.705 ;
        RECT 711.530 242.405 711.830 242.705 ;
        RECT 712.130 242.405 712.430 242.705 ;
        RECT 712.730 242.405 713.030 242.705 ;
        RECT 713.330 242.405 713.630 242.705 ;
        RECT 713.930 242.405 714.230 242.705 ;
        RECT 714.530 242.405 714.830 242.705 ;
        RECT 715.130 242.405 715.430 242.705 ;
        RECT 739.280 243.080 739.580 243.380 ;
        RECT 739.880 243.080 740.180 243.380 ;
        RECT 740.480 243.080 740.780 243.380 ;
        RECT 741.080 243.080 741.380 243.380 ;
        RECT 741.680 243.080 741.980 243.380 ;
        RECT 742.280 243.080 742.580 243.380 ;
        RECT 742.880 243.080 743.180 243.380 ;
        RECT 743.480 243.080 743.780 243.380 ;
        RECT 744.080 243.080 744.380 243.380 ;
        RECT 744.680 243.080 744.980 243.380 ;
        RECT 745.280 243.080 745.580 243.380 ;
        RECT 745.880 243.080 746.180 243.380 ;
        RECT 746.480 243.080 746.780 243.380 ;
        RECT 747.080 243.080 747.380 243.380 ;
        RECT 747.680 243.080 747.980 243.380 ;
        RECT 748.280 243.080 748.580 243.380 ;
        RECT 748.880 243.080 749.180 243.380 ;
        RECT 749.480 243.080 749.780 243.380 ;
        RECT 750.080 243.080 750.380 243.380 ;
        RECT 750.680 243.080 750.980 243.380 ;
        RECT 751.280 243.080 751.580 243.380 ;
        RECT 751.880 243.080 752.180 243.380 ;
        RECT 752.480 243.080 752.780 243.380 ;
        RECT 753.080 243.080 753.380 243.380 ;
        RECT 753.680 243.080 753.980 243.380 ;
        RECT 754.280 243.080 754.580 243.380 ;
        RECT 754.880 243.080 755.180 243.380 ;
        RECT 755.480 243.080 755.780 243.380 ;
        RECT 756.080 243.080 756.380 243.380 ;
        RECT 756.680 243.080 756.980 243.380 ;
        RECT 757.280 243.080 757.580 243.380 ;
        RECT 757.880 243.080 758.180 243.380 ;
        RECT 758.480 243.080 758.780 243.380 ;
        RECT 759.080 243.080 759.380 243.380 ;
        RECT 759.680 243.080 759.980 243.380 ;
        RECT 760.280 243.080 760.580 243.380 ;
        RECT 760.880 243.080 761.180 243.380 ;
        RECT 761.480 243.080 761.780 243.380 ;
        RECT 762.080 243.080 762.380 243.380 ;
        RECT 762.680 243.080 762.980 243.380 ;
        RECT 763.280 243.080 763.580 243.380 ;
        RECT 763.880 243.080 764.180 243.380 ;
        RECT 764.480 243.080 764.780 243.380 ;
        RECT 765.080 243.080 765.380 243.380 ;
        RECT 765.680 243.080 765.980 243.380 ;
        RECT 739.280 242.480 739.580 242.780 ;
        RECT 739.880 242.480 740.180 242.780 ;
        RECT 740.480 242.480 740.780 242.780 ;
        RECT 741.080 242.480 741.380 242.780 ;
        RECT 741.680 242.480 741.980 242.780 ;
        RECT 742.280 242.480 742.580 242.780 ;
        RECT 742.880 242.480 743.180 242.780 ;
        RECT 743.480 242.480 743.780 242.780 ;
        RECT 744.080 242.480 744.380 242.780 ;
        RECT 744.680 242.480 744.980 242.780 ;
        RECT 745.280 242.480 745.580 242.780 ;
        RECT 745.880 242.480 746.180 242.780 ;
        RECT 746.480 242.480 746.780 242.780 ;
        RECT 747.080 242.480 747.380 242.780 ;
        RECT 747.680 242.480 747.980 242.780 ;
        RECT 748.280 242.480 748.580 242.780 ;
        RECT 748.880 242.480 749.180 242.780 ;
        RECT 749.480 242.480 749.780 242.780 ;
        RECT 750.080 242.480 750.380 242.780 ;
        RECT 750.680 242.480 750.980 242.780 ;
        RECT 751.280 242.480 751.580 242.780 ;
        RECT 751.880 242.480 752.180 242.780 ;
        RECT 752.480 242.480 752.780 242.780 ;
        RECT 753.080 242.480 753.380 242.780 ;
        RECT 753.680 242.480 753.980 242.780 ;
        RECT 754.280 242.480 754.580 242.780 ;
        RECT 754.880 242.480 755.180 242.780 ;
        RECT 755.480 242.480 755.780 242.780 ;
        RECT 756.080 242.480 756.380 242.780 ;
        RECT 756.680 242.480 756.980 242.780 ;
        RECT 757.280 242.480 757.580 242.780 ;
        RECT 757.880 242.480 758.180 242.780 ;
        RECT 758.480 242.480 758.780 242.780 ;
        RECT 759.080 242.480 759.380 242.780 ;
        RECT 759.680 242.480 759.980 242.780 ;
        RECT 760.280 242.480 760.580 242.780 ;
        RECT 760.880 242.480 761.180 242.780 ;
        RECT 761.480 242.480 761.780 242.780 ;
        RECT 762.080 242.480 762.380 242.780 ;
        RECT 762.680 242.480 762.980 242.780 ;
        RECT 763.280 242.480 763.580 242.780 ;
        RECT 763.880 242.480 764.180 242.780 ;
        RECT 764.480 242.480 764.780 242.780 ;
        RECT 765.080 242.480 765.380 242.780 ;
        RECT 765.680 242.480 765.980 242.780 ;
        RECT 242.760 121.370 244.480 124.270 ;
        RECT 227.320 115.960 228.970 117.770 ;
      LAYER met3 ;
        RECT 683.800 248.480 687.220 248.700 ;
        RECT 673.820 248.170 687.220 248.480 ;
        RECT 667.260 245.200 687.220 248.170 ;
        RECT 667.260 245.150 768.030 245.200 ;
        RECT 661.490 244.980 768.030 245.150 ;
        RECT 661.490 244.840 776.780 244.980 ;
        RECT 339.420 241.200 776.780 244.840 ;
        RECT 339.420 237.480 687.220 241.200 ;
        RECT 767.260 240.860 776.780 241.200 ;
        RECT 339.420 235.910 675.940 237.480 ;
        RECT 683.800 237.310 687.220 237.480 ;
        RECT 339.420 235.350 673.170 235.910 ;
        RECT 661.490 234.150 673.170 235.350 ;
        RECT 241.580 125.120 245.740 126.930 ;
        RECT 241.580 118.630 245.900 125.120 ;
        RECT 227.010 115.490 245.900 118.630 ;
    END
  END vinit
  PIN vbiasr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 33.300697 ;
    PORT
      LAYER li1 ;
        RECT 258.230 20.020 258.400 20.450 ;
        RECT 258.220 19.280 258.460 20.020 ;
        RECT 258.230 18.590 258.400 19.280 ;
        RECT 258.090 18.140 258.470 18.590 ;
        RECT 258.230 15.580 258.400 18.140 ;
        RECT 694.260 1.470 694.430 6.510 ;
        RECT 696.840 1.470 697.010 6.510 ;
        RECT 699.420 1.470 699.590 6.510 ;
        RECT 702.000 1.470 702.170 6.510 ;
        RECT 704.580 1.470 704.750 6.510 ;
        RECT 707.160 1.470 707.330 6.510 ;
        RECT 709.740 1.470 709.910 6.510 ;
        RECT 712.320 1.470 712.490 6.510 ;
        RECT 714.900 1.470 715.070 6.510 ;
        RECT 717.480 1.470 717.650 6.510 ;
        RECT 720.060 1.470 720.230 6.510 ;
        RECT 745.060 1.640 745.230 6.680 ;
        RECT 747.640 1.640 747.810 6.680 ;
        RECT 750.220 1.640 750.390 6.680 ;
        RECT 752.800 1.640 752.970 6.680 ;
        RECT 755.380 1.640 755.550 6.680 ;
        RECT 757.960 1.640 758.130 6.680 ;
        RECT 760.540 1.640 760.710 6.680 ;
        RECT 763.120 1.640 763.290 6.680 ;
        RECT 765.700 1.640 765.870 6.680 ;
        RECT 768.280 1.640 768.450 6.680 ;
        RECT 770.860 1.640 771.030 6.680 ;
      LAYER mcon ;
        RECT 258.230 15.660 258.400 20.370 ;
        RECT 694.260 1.550 694.430 6.430 ;
        RECT 696.840 1.550 697.010 6.430 ;
        RECT 699.420 1.550 699.590 6.430 ;
        RECT 702.000 1.550 702.170 6.430 ;
        RECT 704.580 1.550 704.750 6.430 ;
        RECT 707.160 1.550 707.330 6.430 ;
        RECT 709.740 1.550 709.910 6.430 ;
        RECT 712.320 1.550 712.490 6.430 ;
        RECT 714.900 1.550 715.070 6.430 ;
        RECT 717.480 1.550 717.650 6.430 ;
        RECT 720.060 1.550 720.230 6.430 ;
        RECT 745.060 1.720 745.230 6.600 ;
        RECT 747.640 1.720 747.810 6.600 ;
        RECT 750.220 1.720 750.390 6.600 ;
        RECT 752.800 1.720 752.970 6.600 ;
        RECT 755.380 1.720 755.550 6.600 ;
        RECT 757.960 1.720 758.130 6.600 ;
        RECT 760.540 1.720 760.710 6.600 ;
        RECT 763.120 1.720 763.290 6.600 ;
        RECT 765.700 1.720 765.870 6.600 ;
        RECT 768.280 1.720 768.450 6.600 ;
        RECT 770.860 1.720 771.030 6.600 ;
      LAYER met1 ;
        RECT 258.140 18.590 258.460 20.420 ;
        RECT 258.090 18.140 258.470 18.590 ;
        RECT 258.140 18.000 258.460 18.140 ;
        RECT 257.750 17.730 258.460 18.000 ;
        RECT 258.140 16.310 258.460 17.730 ;
        RECT 255.750 16.000 258.460 16.310 ;
        RECT 255.750 15.600 258.470 16.000 ;
        RECT 255.750 15.570 258.390 15.600 ;
        RECT 255.770 9.970 256.740 15.570 ;
        RECT 255.770 9.220 256.900 9.970 ;
        RECT 255.720 3.820 257.020 9.220 ;
        RECT 255.780 -0.190 256.900 3.820 ;
        RECT 694.230 0.865 694.460 6.490 ;
        RECT 696.810 0.865 697.040 6.490 ;
        RECT 699.390 0.865 699.620 6.490 ;
        RECT 701.970 0.865 702.200 6.490 ;
        RECT 704.550 0.865 704.780 6.490 ;
        RECT 707.130 0.865 707.360 6.490 ;
        RECT 709.710 0.865 709.940 6.490 ;
        RECT 712.290 0.865 712.520 6.490 ;
        RECT 714.870 0.865 715.100 6.490 ;
        RECT 717.450 0.865 717.680 6.490 ;
        RECT 720.030 0.865 720.260 6.490 ;
        RECT 745.030 0.940 745.260 6.660 ;
        RECT 747.610 0.940 747.840 6.660 ;
        RECT 750.190 0.940 750.420 6.660 ;
        RECT 752.770 0.940 753.000 6.660 ;
        RECT 755.350 0.940 755.580 6.660 ;
        RECT 757.930 0.940 758.160 6.660 ;
        RECT 760.510 0.940 760.740 6.660 ;
        RECT 763.090 0.940 763.320 6.660 ;
        RECT 765.670 0.940 765.900 6.660 ;
        RECT 768.250 0.940 768.480 6.660 ;
        RECT 770.830 0.940 771.060 6.660 ;
        RECT 255.670 -3.990 256.920 -0.190 ;
        RECT 693.510 -0.510 720.980 0.865 ;
        RECT 744.310 -0.435 771.780 0.940 ;
        RECT 254.540 -6.930 260.390 -3.990 ;
      LAYER via ;
        RECT 694.020 0.285 694.320 0.585 ;
        RECT 694.620 0.285 694.920 0.585 ;
        RECT 695.220 0.285 695.520 0.585 ;
        RECT 695.820 0.285 696.120 0.585 ;
        RECT 696.420 0.285 696.720 0.585 ;
        RECT 697.020 0.285 697.320 0.585 ;
        RECT 697.620 0.285 697.920 0.585 ;
        RECT 698.220 0.285 698.520 0.585 ;
        RECT 698.820 0.285 699.120 0.585 ;
        RECT 699.420 0.285 699.720 0.585 ;
        RECT 700.020 0.285 700.320 0.585 ;
        RECT 700.620 0.285 700.920 0.585 ;
        RECT 701.220 0.285 701.520 0.585 ;
        RECT 701.820 0.285 702.120 0.585 ;
        RECT 702.420 0.285 702.720 0.585 ;
        RECT 703.020 0.285 703.320 0.585 ;
        RECT 703.620 0.285 703.920 0.585 ;
        RECT 704.220 0.285 704.520 0.585 ;
        RECT 704.820 0.285 705.120 0.585 ;
        RECT 705.420 0.285 705.720 0.585 ;
        RECT 706.020 0.285 706.320 0.585 ;
        RECT 706.620 0.285 706.920 0.585 ;
        RECT 707.220 0.285 707.520 0.585 ;
        RECT 707.820 0.285 708.120 0.585 ;
        RECT 708.420 0.285 708.720 0.585 ;
        RECT 709.020 0.285 709.320 0.585 ;
        RECT 709.620 0.285 709.920 0.585 ;
        RECT 710.220 0.285 710.520 0.585 ;
        RECT 710.820 0.285 711.120 0.585 ;
        RECT 711.420 0.285 711.720 0.585 ;
        RECT 712.020 0.285 712.320 0.585 ;
        RECT 712.620 0.285 712.920 0.585 ;
        RECT 713.220 0.285 713.520 0.585 ;
        RECT 713.820 0.285 714.120 0.585 ;
        RECT 714.420 0.285 714.720 0.585 ;
        RECT 715.020 0.285 715.320 0.585 ;
        RECT 715.620 0.285 715.920 0.585 ;
        RECT 716.220 0.285 716.520 0.585 ;
        RECT 716.820 0.285 717.120 0.585 ;
        RECT 717.420 0.285 717.720 0.585 ;
        RECT 718.020 0.285 718.320 0.585 ;
        RECT 718.620 0.285 718.920 0.585 ;
        RECT 719.220 0.285 719.520 0.585 ;
        RECT 719.820 0.285 720.120 0.585 ;
        RECT 720.420 0.285 720.720 0.585 ;
        RECT 694.020 -0.315 694.320 -0.015 ;
        RECT 694.620 -0.315 694.920 -0.015 ;
        RECT 695.220 -0.315 695.520 -0.015 ;
        RECT 695.820 -0.315 696.120 -0.015 ;
        RECT 696.420 -0.315 696.720 -0.015 ;
        RECT 697.020 -0.315 697.320 -0.015 ;
        RECT 697.620 -0.315 697.920 -0.015 ;
        RECT 698.220 -0.315 698.520 -0.015 ;
        RECT 698.820 -0.315 699.120 -0.015 ;
        RECT 699.420 -0.315 699.720 -0.015 ;
        RECT 700.020 -0.315 700.320 -0.015 ;
        RECT 700.620 -0.315 700.920 -0.015 ;
        RECT 701.220 -0.315 701.520 -0.015 ;
        RECT 701.820 -0.315 702.120 -0.015 ;
        RECT 702.420 -0.315 702.720 -0.015 ;
        RECT 703.020 -0.315 703.320 -0.015 ;
        RECT 703.620 -0.315 703.920 -0.015 ;
        RECT 704.220 -0.315 704.520 -0.015 ;
        RECT 704.820 -0.315 705.120 -0.015 ;
        RECT 705.420 -0.315 705.720 -0.015 ;
        RECT 706.020 -0.315 706.320 -0.015 ;
        RECT 706.620 -0.315 706.920 -0.015 ;
        RECT 707.220 -0.315 707.520 -0.015 ;
        RECT 707.820 -0.315 708.120 -0.015 ;
        RECT 708.420 -0.315 708.720 -0.015 ;
        RECT 709.020 -0.315 709.320 -0.015 ;
        RECT 709.620 -0.315 709.920 -0.015 ;
        RECT 710.220 -0.315 710.520 -0.015 ;
        RECT 710.820 -0.315 711.120 -0.015 ;
        RECT 711.420 -0.315 711.720 -0.015 ;
        RECT 712.020 -0.315 712.320 -0.015 ;
        RECT 712.620 -0.315 712.920 -0.015 ;
        RECT 713.220 -0.315 713.520 -0.015 ;
        RECT 713.820 -0.315 714.120 -0.015 ;
        RECT 714.420 -0.315 714.720 -0.015 ;
        RECT 715.020 -0.315 715.320 -0.015 ;
        RECT 715.620 -0.315 715.920 -0.015 ;
        RECT 716.220 -0.315 716.520 -0.015 ;
        RECT 716.820 -0.315 717.120 -0.015 ;
        RECT 717.420 -0.315 717.720 -0.015 ;
        RECT 718.020 -0.315 718.320 -0.015 ;
        RECT 718.620 -0.315 718.920 -0.015 ;
        RECT 719.220 -0.315 719.520 -0.015 ;
        RECT 719.820 -0.315 720.120 -0.015 ;
        RECT 720.420 -0.315 720.720 -0.015 ;
        RECT 744.570 0.360 744.870 0.660 ;
        RECT 745.170 0.360 745.470 0.660 ;
        RECT 745.770 0.360 746.070 0.660 ;
        RECT 746.370 0.360 746.670 0.660 ;
        RECT 746.970 0.360 747.270 0.660 ;
        RECT 747.570 0.360 747.870 0.660 ;
        RECT 748.170 0.360 748.470 0.660 ;
        RECT 748.770 0.360 749.070 0.660 ;
        RECT 749.370 0.360 749.670 0.660 ;
        RECT 749.970 0.360 750.270 0.660 ;
        RECT 750.570 0.360 750.870 0.660 ;
        RECT 751.170 0.360 751.470 0.660 ;
        RECT 751.770 0.360 752.070 0.660 ;
        RECT 752.370 0.360 752.670 0.660 ;
        RECT 752.970 0.360 753.270 0.660 ;
        RECT 753.570 0.360 753.870 0.660 ;
        RECT 754.170 0.360 754.470 0.660 ;
        RECT 754.770 0.360 755.070 0.660 ;
        RECT 755.370 0.360 755.670 0.660 ;
        RECT 755.970 0.360 756.270 0.660 ;
        RECT 756.570 0.360 756.870 0.660 ;
        RECT 757.170 0.360 757.470 0.660 ;
        RECT 757.770 0.360 758.070 0.660 ;
        RECT 758.370 0.360 758.670 0.660 ;
        RECT 758.970 0.360 759.270 0.660 ;
        RECT 759.570 0.360 759.870 0.660 ;
        RECT 760.170 0.360 760.470 0.660 ;
        RECT 760.770 0.360 761.070 0.660 ;
        RECT 761.370 0.360 761.670 0.660 ;
        RECT 761.970 0.360 762.270 0.660 ;
        RECT 762.570 0.360 762.870 0.660 ;
        RECT 763.170 0.360 763.470 0.660 ;
        RECT 763.770 0.360 764.070 0.660 ;
        RECT 764.370 0.360 764.670 0.660 ;
        RECT 764.970 0.360 765.270 0.660 ;
        RECT 765.570 0.360 765.870 0.660 ;
        RECT 766.170 0.360 766.470 0.660 ;
        RECT 766.770 0.360 767.070 0.660 ;
        RECT 767.370 0.360 767.670 0.660 ;
        RECT 767.970 0.360 768.270 0.660 ;
        RECT 768.570 0.360 768.870 0.660 ;
        RECT 769.170 0.360 769.470 0.660 ;
        RECT 769.770 0.360 770.070 0.660 ;
        RECT 770.370 0.360 770.670 0.660 ;
        RECT 770.970 0.360 771.270 0.660 ;
        RECT 744.570 -0.240 744.870 0.060 ;
        RECT 745.170 -0.240 745.470 0.060 ;
        RECT 745.770 -0.240 746.070 0.060 ;
        RECT 746.370 -0.240 746.670 0.060 ;
        RECT 746.970 -0.240 747.270 0.060 ;
        RECT 747.570 -0.240 747.870 0.060 ;
        RECT 748.170 -0.240 748.470 0.060 ;
        RECT 748.770 -0.240 749.070 0.060 ;
        RECT 749.370 -0.240 749.670 0.060 ;
        RECT 749.970 -0.240 750.270 0.060 ;
        RECT 750.570 -0.240 750.870 0.060 ;
        RECT 751.170 -0.240 751.470 0.060 ;
        RECT 751.770 -0.240 752.070 0.060 ;
        RECT 752.370 -0.240 752.670 0.060 ;
        RECT 752.970 -0.240 753.270 0.060 ;
        RECT 753.570 -0.240 753.870 0.060 ;
        RECT 754.170 -0.240 754.470 0.060 ;
        RECT 754.770 -0.240 755.070 0.060 ;
        RECT 755.370 -0.240 755.670 0.060 ;
        RECT 755.970 -0.240 756.270 0.060 ;
        RECT 756.570 -0.240 756.870 0.060 ;
        RECT 757.170 -0.240 757.470 0.060 ;
        RECT 757.770 -0.240 758.070 0.060 ;
        RECT 758.370 -0.240 758.670 0.060 ;
        RECT 758.970 -0.240 759.270 0.060 ;
        RECT 759.570 -0.240 759.870 0.060 ;
        RECT 760.170 -0.240 760.470 0.060 ;
        RECT 760.770 -0.240 761.070 0.060 ;
        RECT 761.370 -0.240 761.670 0.060 ;
        RECT 761.970 -0.240 762.270 0.060 ;
        RECT 762.570 -0.240 762.870 0.060 ;
        RECT 763.170 -0.240 763.470 0.060 ;
        RECT 763.770 -0.240 764.070 0.060 ;
        RECT 764.370 -0.240 764.670 0.060 ;
        RECT 764.970 -0.240 765.270 0.060 ;
        RECT 765.570 -0.240 765.870 0.060 ;
        RECT 766.170 -0.240 766.470 0.060 ;
        RECT 766.770 -0.240 767.070 0.060 ;
        RECT 767.370 -0.240 767.670 0.060 ;
        RECT 767.970 -0.240 768.270 0.060 ;
        RECT 768.570 -0.240 768.870 0.060 ;
        RECT 769.170 -0.240 769.470 0.060 ;
        RECT 769.770 -0.240 770.070 0.060 ;
        RECT 770.370 -0.240 770.670 0.060 ;
        RECT 770.970 -0.240 771.270 0.060 ;
        RECT 255.670 -5.880 258.940 -4.350 ;
      LAYER met2 ;
        RECT 693.420 -0.615 721.020 0.885 ;
        RECT 744.270 -0.540 771.870 0.960 ;
        RECT 255.340 -6.160 259.220 -4.100 ;
      LAYER via2 ;
        RECT 694.020 0.285 694.320 0.585 ;
        RECT 694.620 0.285 694.920 0.585 ;
        RECT 695.220 0.285 695.520 0.585 ;
        RECT 695.820 0.285 696.120 0.585 ;
        RECT 696.420 0.285 696.720 0.585 ;
        RECT 697.020 0.285 697.320 0.585 ;
        RECT 697.620 0.285 697.920 0.585 ;
        RECT 698.220 0.285 698.520 0.585 ;
        RECT 698.820 0.285 699.120 0.585 ;
        RECT 699.420 0.285 699.720 0.585 ;
        RECT 700.020 0.285 700.320 0.585 ;
        RECT 700.620 0.285 700.920 0.585 ;
        RECT 701.220 0.285 701.520 0.585 ;
        RECT 701.820 0.285 702.120 0.585 ;
        RECT 702.420 0.285 702.720 0.585 ;
        RECT 703.020 0.285 703.320 0.585 ;
        RECT 703.620 0.285 703.920 0.585 ;
        RECT 704.220 0.285 704.520 0.585 ;
        RECT 704.820 0.285 705.120 0.585 ;
        RECT 705.420 0.285 705.720 0.585 ;
        RECT 706.020 0.285 706.320 0.585 ;
        RECT 706.620 0.285 706.920 0.585 ;
        RECT 707.220 0.285 707.520 0.585 ;
        RECT 707.820 0.285 708.120 0.585 ;
        RECT 708.420 0.285 708.720 0.585 ;
        RECT 709.020 0.285 709.320 0.585 ;
        RECT 709.620 0.285 709.920 0.585 ;
        RECT 710.220 0.285 710.520 0.585 ;
        RECT 710.820 0.285 711.120 0.585 ;
        RECT 711.420 0.285 711.720 0.585 ;
        RECT 712.020 0.285 712.320 0.585 ;
        RECT 712.620 0.285 712.920 0.585 ;
        RECT 713.220 0.285 713.520 0.585 ;
        RECT 713.820 0.285 714.120 0.585 ;
        RECT 714.420 0.285 714.720 0.585 ;
        RECT 715.020 0.285 715.320 0.585 ;
        RECT 715.620 0.285 715.920 0.585 ;
        RECT 716.220 0.285 716.520 0.585 ;
        RECT 716.820 0.285 717.120 0.585 ;
        RECT 717.420 0.285 717.720 0.585 ;
        RECT 718.020 0.285 718.320 0.585 ;
        RECT 718.620 0.285 718.920 0.585 ;
        RECT 719.220 0.285 719.520 0.585 ;
        RECT 719.820 0.285 720.120 0.585 ;
        RECT 720.420 0.285 720.720 0.585 ;
        RECT 694.020 -0.315 694.320 -0.015 ;
        RECT 694.620 -0.315 694.920 -0.015 ;
        RECT 695.220 -0.315 695.520 -0.015 ;
        RECT 695.820 -0.315 696.120 -0.015 ;
        RECT 696.420 -0.315 696.720 -0.015 ;
        RECT 697.020 -0.315 697.320 -0.015 ;
        RECT 697.620 -0.315 697.920 -0.015 ;
        RECT 698.220 -0.315 698.520 -0.015 ;
        RECT 698.820 -0.315 699.120 -0.015 ;
        RECT 699.420 -0.315 699.720 -0.015 ;
        RECT 700.020 -0.315 700.320 -0.015 ;
        RECT 700.620 -0.315 700.920 -0.015 ;
        RECT 701.220 -0.315 701.520 -0.015 ;
        RECT 701.820 -0.315 702.120 -0.015 ;
        RECT 702.420 -0.315 702.720 -0.015 ;
        RECT 703.020 -0.315 703.320 -0.015 ;
        RECT 703.620 -0.315 703.920 -0.015 ;
        RECT 704.220 -0.315 704.520 -0.015 ;
        RECT 704.820 -0.315 705.120 -0.015 ;
        RECT 705.420 -0.315 705.720 -0.015 ;
        RECT 706.020 -0.315 706.320 -0.015 ;
        RECT 706.620 -0.315 706.920 -0.015 ;
        RECT 707.220 -0.315 707.520 -0.015 ;
        RECT 707.820 -0.315 708.120 -0.015 ;
        RECT 708.420 -0.315 708.720 -0.015 ;
        RECT 709.020 -0.315 709.320 -0.015 ;
        RECT 709.620 -0.315 709.920 -0.015 ;
        RECT 710.220 -0.315 710.520 -0.015 ;
        RECT 710.820 -0.315 711.120 -0.015 ;
        RECT 711.420 -0.315 711.720 -0.015 ;
        RECT 712.020 -0.315 712.320 -0.015 ;
        RECT 712.620 -0.315 712.920 -0.015 ;
        RECT 713.220 -0.315 713.520 -0.015 ;
        RECT 713.820 -0.315 714.120 -0.015 ;
        RECT 714.420 -0.315 714.720 -0.015 ;
        RECT 715.020 -0.315 715.320 -0.015 ;
        RECT 715.620 -0.315 715.920 -0.015 ;
        RECT 716.220 -0.315 716.520 -0.015 ;
        RECT 716.820 -0.315 717.120 -0.015 ;
        RECT 717.420 -0.315 717.720 -0.015 ;
        RECT 718.020 -0.315 718.320 -0.015 ;
        RECT 718.620 -0.315 718.920 -0.015 ;
        RECT 719.220 -0.315 719.520 -0.015 ;
        RECT 719.820 -0.315 720.120 -0.015 ;
        RECT 720.420 -0.315 720.720 -0.015 ;
        RECT 744.570 0.360 744.870 0.660 ;
        RECT 745.170 0.360 745.470 0.660 ;
        RECT 745.770 0.360 746.070 0.660 ;
        RECT 746.370 0.360 746.670 0.660 ;
        RECT 746.970 0.360 747.270 0.660 ;
        RECT 747.570 0.360 747.870 0.660 ;
        RECT 748.170 0.360 748.470 0.660 ;
        RECT 748.770 0.360 749.070 0.660 ;
        RECT 749.370 0.360 749.670 0.660 ;
        RECT 749.970 0.360 750.270 0.660 ;
        RECT 750.570 0.360 750.870 0.660 ;
        RECT 751.170 0.360 751.470 0.660 ;
        RECT 751.770 0.360 752.070 0.660 ;
        RECT 752.370 0.360 752.670 0.660 ;
        RECT 752.970 0.360 753.270 0.660 ;
        RECT 753.570 0.360 753.870 0.660 ;
        RECT 754.170 0.360 754.470 0.660 ;
        RECT 754.770 0.360 755.070 0.660 ;
        RECT 755.370 0.360 755.670 0.660 ;
        RECT 755.970 0.360 756.270 0.660 ;
        RECT 756.570 0.360 756.870 0.660 ;
        RECT 757.170 0.360 757.470 0.660 ;
        RECT 757.770 0.360 758.070 0.660 ;
        RECT 758.370 0.360 758.670 0.660 ;
        RECT 758.970 0.360 759.270 0.660 ;
        RECT 759.570 0.360 759.870 0.660 ;
        RECT 760.170 0.360 760.470 0.660 ;
        RECT 760.770 0.360 761.070 0.660 ;
        RECT 761.370 0.360 761.670 0.660 ;
        RECT 761.970 0.360 762.270 0.660 ;
        RECT 762.570 0.360 762.870 0.660 ;
        RECT 763.170 0.360 763.470 0.660 ;
        RECT 763.770 0.360 764.070 0.660 ;
        RECT 764.370 0.360 764.670 0.660 ;
        RECT 764.970 0.360 765.270 0.660 ;
        RECT 765.570 0.360 765.870 0.660 ;
        RECT 766.170 0.360 766.470 0.660 ;
        RECT 766.770 0.360 767.070 0.660 ;
        RECT 767.370 0.360 767.670 0.660 ;
        RECT 767.970 0.360 768.270 0.660 ;
        RECT 768.570 0.360 768.870 0.660 ;
        RECT 769.170 0.360 769.470 0.660 ;
        RECT 769.770 0.360 770.070 0.660 ;
        RECT 770.370 0.360 770.670 0.660 ;
        RECT 770.970 0.360 771.270 0.660 ;
        RECT 744.570 -0.240 744.870 0.060 ;
        RECT 745.170 -0.240 745.470 0.060 ;
        RECT 745.770 -0.240 746.070 0.060 ;
        RECT 746.370 -0.240 746.670 0.060 ;
        RECT 746.970 -0.240 747.270 0.060 ;
        RECT 747.570 -0.240 747.870 0.060 ;
        RECT 748.170 -0.240 748.470 0.060 ;
        RECT 748.770 -0.240 749.070 0.060 ;
        RECT 749.370 -0.240 749.670 0.060 ;
        RECT 749.970 -0.240 750.270 0.060 ;
        RECT 750.570 -0.240 750.870 0.060 ;
        RECT 751.170 -0.240 751.470 0.060 ;
        RECT 751.770 -0.240 752.070 0.060 ;
        RECT 752.370 -0.240 752.670 0.060 ;
        RECT 752.970 -0.240 753.270 0.060 ;
        RECT 753.570 -0.240 753.870 0.060 ;
        RECT 754.170 -0.240 754.470 0.060 ;
        RECT 754.770 -0.240 755.070 0.060 ;
        RECT 755.370 -0.240 755.670 0.060 ;
        RECT 755.970 -0.240 756.270 0.060 ;
        RECT 756.570 -0.240 756.870 0.060 ;
        RECT 757.170 -0.240 757.470 0.060 ;
        RECT 757.770 -0.240 758.070 0.060 ;
        RECT 758.370 -0.240 758.670 0.060 ;
        RECT 758.970 -0.240 759.270 0.060 ;
        RECT 759.570 -0.240 759.870 0.060 ;
        RECT 760.170 -0.240 760.470 0.060 ;
        RECT 760.770 -0.240 761.070 0.060 ;
        RECT 761.370 -0.240 761.670 0.060 ;
        RECT 761.970 -0.240 762.270 0.060 ;
        RECT 762.570 -0.240 762.870 0.060 ;
        RECT 763.170 -0.240 763.470 0.060 ;
        RECT 763.770 -0.240 764.070 0.060 ;
        RECT 764.370 -0.240 764.670 0.060 ;
        RECT 764.970 -0.240 765.270 0.060 ;
        RECT 765.570 -0.240 765.870 0.060 ;
        RECT 766.170 -0.240 766.470 0.060 ;
        RECT 766.770 -0.240 767.070 0.060 ;
        RECT 767.370 -0.240 767.670 0.060 ;
        RECT 767.970 -0.240 768.270 0.060 ;
        RECT 768.570 -0.240 768.870 0.060 ;
        RECT 769.170 -0.240 769.470 0.060 ;
        RECT 769.770 -0.240 770.070 0.060 ;
        RECT 770.370 -0.240 770.670 0.060 ;
        RECT 770.970 -0.240 771.270 0.060 ;
        RECT 255.520 -6.000 259.050 -4.220 ;
      LAYER met3 ;
        RECT 690.750 2.480 692.370 2.520 ;
        RECT 771.950 2.480 787.000 2.770 ;
        RECT 670.670 2.050 677.110 2.140 ;
        RECT 690.750 2.050 787.000 2.480 ;
        RECT 670.670 -1.280 787.000 2.050 ;
        RECT 255.100 -1.520 787.000 -1.280 ;
        RECT 255.100 -2.630 692.370 -1.520 ;
        RECT 771.950 -1.910 787.000 -1.520 ;
        RECT 255.100 -2.800 691.120 -2.630 ;
        RECT 255.100 -6.130 677.110 -2.800 ;
        RECT 255.340 -6.160 259.220 -6.130 ;
        RECT 670.670 -6.400 677.110 -6.130 ;
    END
  END vbiasr
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER li1 ;
        RECT 310.775 131.660 311.080 132.365 ;
        RECT 313.665 132.160 314.110 132.330 ;
        RECT 316.950 132.160 317.240 132.490 ;
        RECT 313.685 132.000 314.110 132.160 ;
        RECT 324.465 131.695 324.770 132.400 ;
        RECT 327.355 132.195 327.800 132.365 ;
        RECT 330.640 132.195 330.930 132.525 ;
        RECT 327.375 132.035 327.800 132.195 ;
        RECT 322.575 125.595 322.880 126.300 ;
        RECT 325.465 126.095 325.910 126.265 ;
        RECT 328.750 126.095 329.040 126.425 ;
        RECT 325.485 125.935 325.910 126.095 ;
      LAYER mcon ;
        RECT 310.785 132.160 310.955 132.330 ;
        RECT 317.025 132.160 317.195 132.330 ;
        RECT 324.475 132.195 324.645 132.365 ;
        RECT 330.715 132.195 330.885 132.365 ;
        RECT 322.585 126.095 322.755 126.265 ;
        RECT 328.825 126.095 328.995 126.265 ;
      LAYER met1 ;
        RECT 310.660 132.315 311.040 132.440 ;
        RECT 313.605 132.315 313.895 132.360 ;
        RECT 316.965 132.315 317.255 132.360 ;
        RECT 310.660 132.175 317.255 132.315 ;
        RECT 310.660 132.090 311.040 132.175 ;
        RECT 313.605 132.130 313.895 132.175 ;
        RECT 316.965 132.130 317.255 132.175 ;
        RECT 324.280 132.350 324.810 132.530 ;
        RECT 327.295 132.350 327.585 132.395 ;
        RECT 330.655 132.350 330.945 132.395 ;
        RECT 324.280 132.210 330.945 132.350 ;
        RECT 324.280 132.080 324.810 132.210 ;
        RECT 327.295 132.165 327.585 132.210 ;
        RECT 330.655 132.165 330.945 132.210 ;
        RECT 322.350 126.250 322.930 126.430 ;
        RECT 325.405 126.250 325.695 126.295 ;
        RECT 328.765 126.250 329.055 126.295 ;
        RECT 322.350 126.110 329.055 126.250 ;
        RECT 322.350 125.950 322.930 126.110 ;
        RECT 325.405 126.065 325.695 126.110 ;
        RECT 328.765 126.065 329.055 126.110 ;
      LAYER via ;
        RECT 310.710 132.120 311.000 132.390 ;
        RECT 324.350 132.140 324.750 132.480 ;
        RECT 322.400 126.000 322.890 126.380 ;
      LAYER met2 ;
        RECT 320.120 371.560 323.250 392.160 ;
        RECT 320.120 368.130 324.600 371.560 ;
        RECT 320.180 366.170 324.600 368.130 ;
        RECT 320.840 285.850 324.540 366.170 ;
        RECT 320.140 221.850 325.130 285.850 ;
        RECT 320.270 220.110 325.130 221.850 ;
        RECT 320.270 165.280 324.970 220.110 ;
        RECT 320.140 150.850 325.090 165.280 ;
        RECT 320.510 138.650 322.460 140.190 ;
        RECT 320.930 137.050 321.660 138.650 ;
        RECT 320.880 134.600 321.720 137.050 ;
        RECT 320.770 134.170 321.800 134.600 ;
        RECT 310.660 133.920 322.140 134.170 ;
        RECT 310.660 132.440 310.980 133.920 ;
        RECT 321.760 132.500 322.090 133.920 ;
        RECT 324.280 132.500 324.810 132.530 ;
        RECT 310.660 132.090 311.040 132.440 ;
        RECT 321.760 132.140 324.810 132.500 ;
        RECT 321.760 132.100 322.090 132.140 ;
        RECT 322.350 126.430 322.730 132.140 ;
        RECT 324.280 132.080 324.810 132.140 ;
        RECT 322.350 125.950 322.930 126.430 ;
      LAYER via2 ;
        RECT 320.710 368.450 322.630 369.310 ;
        RECT 320.900 151.370 321.870 152.060 ;
        RECT 321.120 139.290 321.520 139.730 ;
      LAYER met3 ;
        RECT 320.350 368.340 323.090 369.580 ;
        RECT 320.320 150.880 322.550 152.500 ;
        RECT 320.840 141.030 321.660 150.880 ;
        RECT 320.460 139.100 322.500 141.030 ;
    END
  END reset
  PIN v9m
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.389200 ;
    PORT
      LAYER li1 ;
        RECT 27.630 69.060 29.350 69.230 ;
        RECT 27.660 66.530 29.380 66.700 ;
        RECT 27.650 63.940 29.370 64.110 ;
        RECT 27.650 61.390 29.370 61.560 ;
        RECT 27.650 58.840 29.370 59.010 ;
        RECT 21.550 56.940 24.830 57.110 ;
        RECT 27.650 56.290 29.370 56.460 ;
        RECT 27.650 53.740 29.370 53.910 ;
        RECT 27.650 51.190 29.370 51.360 ;
        RECT 27.650 48.640 29.370 48.810 ;
      LAYER mcon ;
        RECT 27.710 69.060 29.270 69.230 ;
        RECT 27.740 66.530 29.300 66.700 ;
        RECT 27.730 63.940 29.290 64.110 ;
        RECT 27.730 61.390 29.290 61.560 ;
        RECT 27.730 58.840 29.290 59.010 ;
        RECT 21.630 56.940 22.380 57.110 ;
        RECT 23.070 56.940 24.750 57.110 ;
        RECT 27.730 56.290 29.290 56.460 ;
        RECT 27.730 53.740 29.290 53.910 ;
        RECT 27.730 51.190 29.290 51.360 ;
        RECT 27.730 48.640 29.290 48.810 ;
      LAYER met1 ;
        RECT 27.670 69.260 29.300 69.290 ;
        RECT 27.650 69.030 29.330 69.260 ;
        RECT 27.670 68.990 29.330 69.030 ;
        RECT 28.990 68.930 29.330 68.990 ;
        RECT 28.990 68.650 31.180 68.930 ;
        RECT 27.680 66.500 29.360 66.730 ;
        RECT 29.060 66.310 29.340 66.500 ;
        RECT 30.790 66.310 31.180 68.650 ;
        RECT 28.900 66.000 31.180 66.310 ;
        RECT 29.100 64.140 29.380 64.180 ;
        RECT 27.670 63.910 29.380 64.140 ;
        RECT 29.100 63.810 29.380 63.910 ;
        RECT 30.790 63.810 31.180 66.000 ;
        RECT 29.100 63.510 31.210 63.810 ;
        RECT 29.110 63.500 31.210 63.510 ;
        RECT 27.670 61.540 29.350 61.590 ;
        RECT 27.670 61.360 29.360 61.540 ;
        RECT 29.080 61.150 29.360 61.360 ;
        RECT 30.790 61.150 31.180 63.500 ;
        RECT 29.060 60.840 31.180 61.150 ;
        RECT 29.800 60.390 30.590 60.480 ;
        RECT 29.800 60.350 30.610 60.390 ;
        RECT 30.790 60.350 31.180 60.840 ;
        RECT 29.800 60.290 31.180 60.350 ;
        RECT 29.790 59.800 31.180 60.290 ;
        RECT 29.790 59.770 30.630 59.800 ;
        RECT 29.800 59.620 30.630 59.770 ;
        RECT 29.800 59.610 30.590 59.620 ;
        RECT 27.670 58.930 29.350 59.040 ;
        RECT 27.670 58.810 29.360 58.930 ;
        RECT 29.050 58.730 29.360 58.810 ;
        RECT 30.790 58.730 31.180 59.800 ;
        RECT 29.050 58.420 31.180 58.730 ;
        RECT 29.050 58.370 29.330 58.420 ;
        RECT 21.600 56.850 24.790 57.200 ;
        RECT 21.600 56.840 24.780 56.850 ;
        RECT 29.010 56.490 29.290 56.500 ;
        RECT 27.670 56.260 29.350 56.490 ;
        RECT 29.010 56.120 29.290 56.260 ;
        RECT 30.790 56.120 31.180 58.420 ;
        RECT 29.010 55.830 31.180 56.120 ;
        RECT 29.080 55.810 31.180 55.830 ;
        RECT 29.090 53.940 29.370 53.970 ;
        RECT 27.670 53.710 29.370 53.940 ;
        RECT 29.090 53.630 29.370 53.710 ;
        RECT 30.790 53.630 31.180 55.810 ;
        RECT 29.090 53.320 31.180 53.630 ;
        RECT 29.090 53.300 29.370 53.320 ;
        RECT 29.100 51.390 29.350 51.410 ;
        RECT 27.670 51.160 29.350 51.390 ;
        RECT 29.100 51.070 29.350 51.160 ;
        RECT 30.790 51.070 31.180 53.320 ;
        RECT 29.100 50.780 31.180 51.070 ;
        RECT 29.120 50.760 31.180 50.780 ;
        RECT 27.670 48.610 29.350 48.840 ;
        RECT 29.060 48.450 29.330 48.610 ;
        RECT 30.790 48.450 31.180 50.760 ;
        RECT 29.060 48.310 31.180 48.450 ;
        RECT 29.060 48.140 31.160 48.310 ;
      LAYER via ;
        RECT 29.900 59.750 30.460 60.370 ;
        RECT 21.630 56.880 24.750 57.160 ;
      LAYER met2 ;
        RECT 29.800 60.390 30.590 60.480 ;
        RECT 29.800 59.980 30.610 60.390 ;
        RECT 29.800 59.620 30.630 59.980 ;
        RECT 29.800 59.610 30.590 59.620 ;
        RECT 21.610 56.820 24.790 57.210 ;
      LAYER via2 ;
        RECT 29.900 59.750 30.460 60.370 ;
        RECT 21.630 56.880 24.750 57.160 ;
      LAYER met3 ;
        RECT 17.890 84.050 22.140 84.230 ;
        RECT -37.770 83.170 22.140 84.050 ;
        RECT -37.770 83.050 22.010 83.170 ;
        RECT 21.350 67.270 22.010 83.050 ;
        RECT 21.400 61.890 22.010 67.270 ;
        RECT 21.370 61.600 22.010 61.890 ;
        RECT 21.370 58.860 21.930 61.600 ;
        RECT 23.930 60.510 24.490 60.550 ;
        RECT 23.930 60.500 29.790 60.510 ;
        RECT 23.930 60.490 30.210 60.500 ;
        RECT 23.850 60.480 30.210 60.490 ;
        RECT 23.850 60.390 30.590 60.480 ;
        RECT 23.850 60.040 30.610 60.390 ;
        RECT 23.850 60.030 26.190 60.040 ;
        RECT 21.360 58.260 21.930 58.860 ;
        RECT 21.360 57.220 21.920 58.260 ;
        RECT 23.930 57.220 24.490 60.030 ;
        RECT 29.790 59.980 30.610 60.040 ;
        RECT 29.790 59.740 30.630 59.980 ;
        RECT 29.800 59.620 30.630 59.740 ;
        RECT 29.800 59.610 30.590 59.620 ;
        RECT 21.360 56.840 24.850 57.220 ;
        RECT 21.570 56.820 24.850 56.840 ;
        RECT 21.570 56.780 24.810 56.820 ;
    END
  END v9m
  PIN Fvco
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.885000 ;
    ANTENNADIFFAREA 0.609000 ;
    PORT
      LAYER li1 ;
        RECT 309.715 131.705 310.095 132.375 ;
        RECT 43.380 50.300 43.550 50.350 ;
        RECT 43.110 50.020 43.550 50.300 ;
        RECT 43.110 49.210 43.280 50.020 ;
        RECT 45.575 49.210 45.745 49.350 ;
        RECT 43.110 49.040 45.750 49.210 ;
        RECT 43.110 49.030 45.745 49.040 ;
        RECT 45.020 48.190 45.200 49.030 ;
        RECT 45.575 49.020 45.745 49.030 ;
        RECT 47.100 48.190 47.710 48.580 ;
        RECT 44.660 48.010 47.860 48.190 ;
        RECT 44.660 47.020 44.830 48.010 ;
        RECT 47.690 47.520 47.860 48.010 ;
        RECT 47.685 47.190 47.860 47.520 ;
        RECT 44.650 46.710 44.830 47.020 ;
        RECT 44.650 46.690 44.820 46.710 ;
        RECT 124.050 14.110 124.220 15.050 ;
        RECT 123.970 10.585 124.140 10.915 ;
      LAYER mcon ;
        RECT 309.740 131.930 309.910 132.100 ;
        RECT 47.190 48.100 47.600 48.510 ;
        RECT 124.050 14.190 124.220 14.970 ;
        RECT 123.970 10.665 124.140 10.835 ;
      LAYER met1 ;
        RECT 303.800 132.850 307.330 133.480 ;
        RECT 303.800 132.120 308.810 132.850 ;
        RECT 309.620 132.120 310.140 132.470 ;
        RECT 303.800 131.880 310.140 132.120 ;
        RECT 303.800 131.770 308.810 131.880 ;
        RECT 309.690 131.850 309.960 131.880 ;
        RECT 303.800 131.410 307.330 131.770 ;
        RECT 47.100 48.020 47.710 48.580 ;
        RECT 124.030 15.030 125.790 15.060 ;
        RECT 124.020 14.170 125.790 15.030 ;
        RECT 124.020 14.130 124.250 14.170 ;
        RECT 125.540 12.680 125.790 14.170 ;
        RECT 126.180 12.680 127.450 12.780 ;
        RECT 125.530 12.210 127.450 12.680 ;
        RECT 125.540 10.930 125.790 12.210 ;
        RECT 123.930 10.910 125.790 10.930 ;
        RECT 123.920 10.620 125.790 10.910 ;
        RECT 123.920 10.590 124.200 10.620 ;
        RECT 125.540 10.590 125.790 10.620 ;
        RECT 126.180 1.270 127.450 12.210 ;
        RECT 126.150 0.200 130.760 1.270 ;
        RECT 126.180 0.170 127.450 0.200 ;
      LAYER via ;
        RECT 304.770 131.900 306.420 132.740 ;
        RECT 47.190 48.100 47.600 48.510 ;
        RECT 129.740 0.320 130.650 1.140 ;
      LAYER met2 ;
        RECT -15.730 -5.540 -10.790 396.040 ;
        RECT 303.800 131.410 307.330 133.480 ;
        RECT 312.680 74.450 313.280 85.750 ;
        RECT 47.100 48.020 47.710 48.580 ;
        RECT 129.610 0.190 130.760 1.270 ;
      LAYER via2 ;
        RECT 304.770 131.900 306.420 132.740 ;
        RECT 312.780 85.250 313.190 85.660 ;
        RECT 312.770 74.550 313.210 74.940 ;
        RECT 47.190 48.100 47.600 48.510 ;
        RECT 129.740 0.320 130.650 1.140 ;
        RECT -14.880 -4.800 -12.420 -3.330 ;
      LAYER met3 ;
        RECT 303.800 131.410 307.330 133.480 ;
        RECT 304.610 122.990 305.610 131.410 ;
        RECT 304.610 122.020 313.390 122.990 ;
        RECT 312.810 106.540 313.170 122.020 ;
        RECT 312.800 106.290 313.170 106.540 ;
        RECT 312.800 93.660 313.160 106.290 ;
        RECT 312.800 89.880 313.170 93.660 ;
        RECT 312.810 85.740 313.170 89.880 ;
        RECT 312.730 85.180 313.250 85.740 ;
        RECT 312.680 74.450 313.280 75.010 ;
        RECT 312.760 61.730 313.180 74.450 ;
        RECT 312.750 61.560 313.180 61.730 ;
        RECT 312.750 55.060 313.170 61.560 ;
        RECT 312.750 54.880 313.180 55.060 ;
        RECT 47.100 48.000 54.590 48.580 ;
        RECT 312.760 48.410 313.180 54.880 ;
        RECT 312.750 48.210 313.180 48.410 ;
        RECT 53.960 34.550 54.570 48.000 ;
        RECT 312.750 42.250 313.170 48.210 ;
        RECT 312.730 41.560 313.170 42.250 ;
        RECT -1.860 -1.730 6.120 -1.240 ;
        RECT 53.090 -1.430 54.950 34.550 ;
        RECT 312.730 28.960 313.150 41.560 ;
        RECT 312.710 28.860 313.150 28.960 ;
        RECT 312.710 22.280 313.130 28.860 ;
        RECT 312.700 22.110 313.130 22.280 ;
        RECT 312.700 9.000 313.120 22.110 ;
        RECT 312.690 8.790 313.120 9.000 ;
        RECT 312.690 2.530 313.110 8.790 ;
        RECT 129.470 0.930 130.780 1.320 ;
        RECT 312.670 0.930 313.130 2.530 ;
        RECT 129.470 0.480 313.130 0.930 ;
        RECT -16.470 -1.860 10.540 -1.730 ;
        RECT 53.090 -1.860 55.330 -1.430 ;
        RECT -16.470 -1.980 62.230 -1.860 ;
        RECT -16.470 -2.270 105.720 -1.980 ;
        RECT 129.470 -2.270 130.780 0.480 ;
        RECT 143.850 0.320 144.150 0.480 ;
        RECT -16.470 -3.150 130.840 -2.270 ;
        RECT -16.470 -3.590 105.720 -3.150 ;
        RECT -16.470 -4.310 62.230 -3.590 ;
        RECT -16.470 -5.910 10.540 -4.310 ;
    END
  END Fvco
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 739.020 243.330 766.490 250.120 ;
        RECT 310.645 131.620 314.395 131.715 ;
        RECT 324.335 131.655 328.085 131.750 ;
        RECT 310.645 131.400 316.180 131.620 ;
        RECT 319.785 131.520 321.155 131.525 ;
        RECT 319.785 131.430 323.070 131.520 ;
        RECT 317.865 131.400 323.070 131.430 ;
        RECT 310.645 131.190 323.070 131.400 ;
        RECT 324.335 131.435 329.870 131.655 ;
        RECT 333.475 131.465 334.845 131.560 ;
        RECT 331.555 131.435 334.845 131.465 ;
        RECT 324.335 131.190 334.845 131.435 ;
        RECT 310.645 131.155 334.845 131.190 ;
        RECT 309.195 130.490 334.845 131.155 ;
        RECT 309.195 130.455 334.880 130.490 ;
        RECT 309.190 130.245 334.880 130.455 ;
        RECT 309.190 130.210 323.070 130.245 ;
        RECT 320.980 130.170 323.070 130.210 ;
        RECT 322.445 125.555 326.195 125.650 ;
        RECT 322.445 125.335 327.980 125.555 ;
        RECT 333.760 125.470 335.270 125.480 ;
        RECT 332.900 125.460 335.270 125.470 ;
        RECT 331.585 125.365 335.270 125.460 ;
        RECT 329.665 125.335 335.270 125.365 ;
        RECT 322.445 125.090 335.270 125.335 ;
        RECT 320.995 124.390 335.270 125.090 ;
        RECT 320.990 124.220 335.270 124.390 ;
        RECT 320.990 124.210 333.860 124.220 ;
        RECT 320.990 124.145 332.990 124.210 ;
        RECT 87.445 110.205 87.505 110.235 ;
        RECT 155.550 110.210 155.610 110.240 ;
        RECT 87.445 18.590 105.695 110.205 ;
        RECT 155.550 18.595 173.800 110.210 ;
        RECT 744.310 0.610 771.780 7.400 ;
      LAYER li1 ;
        RECT 739.200 249.770 766.310 249.940 ;
        RECT 739.200 243.680 739.370 249.770 ;
        RECT 741.060 244.190 741.230 249.400 ;
        RECT 743.640 244.190 743.810 249.400 ;
        RECT 746.220 244.190 746.390 249.400 ;
        RECT 748.800 244.190 748.970 249.400 ;
        RECT 751.380 244.190 751.550 249.400 ;
        RECT 753.960 244.190 754.130 249.400 ;
        RECT 756.540 244.190 756.710 249.400 ;
        RECT 759.120 244.190 759.290 249.400 ;
        RECT 761.700 244.190 761.870 249.400 ;
        RECT 764.280 244.190 764.450 249.400 ;
        RECT 739.765 244.020 765.750 244.190 ;
        RECT 766.140 243.680 766.310 249.770 ;
        RECT 739.200 243.510 766.310 243.680 ;
        RECT 369.540 215.330 378.730 221.480 ;
        RECT 389.540 215.330 398.730 221.480 ;
        RECT 409.540 215.330 418.730 221.480 ;
        RECT 429.540 215.330 438.730 221.480 ;
        RECT 449.540 215.330 458.730 221.480 ;
        RECT 469.540 215.330 478.730 221.480 ;
        RECT 489.540 215.330 498.730 221.480 ;
        RECT 509.540 215.330 518.730 221.480 ;
        RECT 529.540 215.330 538.730 221.480 ;
        RECT 549.540 215.330 558.730 221.480 ;
        RECT 569.540 215.330 578.730 221.480 ;
        RECT 589.540 215.330 598.730 221.480 ;
        RECT 609.540 215.330 618.730 221.480 ;
        RECT 629.540 215.330 638.730 221.480 ;
        RECT 649.540 215.330 658.730 221.480 ;
        RECT 360.860 204.510 370.050 210.660 ;
        RECT 649.750 199.320 658.940 205.510 ;
        RECT 360.860 184.510 370.050 190.660 ;
        RECT 384.360 185.470 384.710 187.630 ;
        RECT 385.950 185.470 386.300 187.630 ;
        RECT 387.540 185.470 387.890 187.630 ;
        RECT 389.130 185.470 389.480 187.630 ;
        RECT 649.750 179.320 658.940 185.510 ;
        RECT 360.860 164.510 370.050 170.660 ;
        RECT 384.360 159.680 384.710 161.840 ;
        RECT 385.950 159.680 386.300 161.840 ;
        RECT 387.540 159.680 387.890 161.840 ;
        RECT 389.130 159.680 389.480 161.840 ;
        RECT 649.750 159.320 658.940 165.510 ;
        RECT 168.470 154.870 171.490 155.280 ;
        RECT 360.860 144.510 370.050 150.660 ;
        RECT 384.620 149.080 384.970 151.240 ;
        RECT 389.980 148.900 390.330 151.060 ;
        RECT 649.750 139.320 658.940 145.510 ;
        RECT 128.400 133.820 128.970 133.830 ;
        RECT 118.670 133.360 128.970 133.820 ;
        RECT 150.300 133.380 150.870 133.390 ;
        RECT 118.690 131.060 119.450 133.360 ;
        RECT 128.400 132.580 128.970 133.360 ;
        RECT 140.570 132.920 150.870 133.380 ;
        RECT 171.090 133.150 171.660 133.160 ;
        RECT 128.400 132.220 129.300 132.580 ;
        RECT 128.470 132.180 129.300 132.220 ;
        RECT 118.690 131.040 121.890 131.060 ;
        RECT 118.660 129.820 121.890 131.040 ;
        RECT 140.590 130.620 141.350 132.920 ;
        RECT 150.300 132.140 150.870 132.920 ;
        RECT 161.360 132.690 171.660 133.150 ;
        RECT 150.300 131.780 151.200 132.140 ;
        RECT 150.370 131.740 151.200 131.780 ;
        RECT 140.590 130.600 143.790 130.620 ;
        RECT 117.290 128.560 121.890 129.820 ;
        RECT 140.560 129.380 143.790 130.600 ;
        RECT 161.380 130.390 162.140 132.690 ;
        RECT 171.090 131.910 171.660 132.690 ;
        RECT 171.090 131.550 171.990 131.910 ;
        RECT 171.160 131.510 171.990 131.550 ;
        RECT 161.380 130.370 164.580 130.390 ;
        RECT 117.460 127.320 121.890 128.560 ;
        RECT 139.190 128.120 143.790 129.380 ;
        RECT 161.350 129.150 164.580 130.370 ;
        RECT 309.760 130.295 310.020 130.965 ;
        RECT 310.765 130.295 311.095 130.910 ;
        RECT 314.435 130.295 314.765 130.760 ;
        RECT 316.645 130.295 316.975 131.225 ;
        RECT 317.955 130.295 318.285 130.860 ;
        RECT 318.815 130.295 319.145 131.320 ;
        RECT 319.850 130.295 320.205 131.335 ;
        RECT 320.770 130.295 321.065 131.415 ;
        RECT 321.400 130.610 322.000 131.140 ;
        RECT 321.560 130.380 321.790 130.610 ;
        RECT 321.560 130.330 323.080 130.380 ;
        RECT 323.450 130.330 323.710 131.000 ;
        RECT 324.455 130.330 324.785 130.945 ;
        RECT 328.125 130.330 328.455 130.795 ;
        RECT 330.335 130.330 330.665 131.260 ;
        RECT 331.645 130.330 331.975 130.895 ;
        RECT 332.505 130.330 332.835 131.355 ;
        RECT 333.540 130.330 333.895 131.370 ;
        RECT 334.460 130.330 334.755 131.450 ;
        RECT 309.190 130.125 321.190 130.295 ;
        RECT 321.560 130.190 334.880 130.330 ;
        RECT 322.880 130.160 334.880 130.190 ;
        RECT 117.460 127.300 121.590 127.320 ;
        RECT 117.460 118.820 120.420 127.300 ;
        RECT 140.560 126.880 143.790 128.120 ;
        RECT 159.980 127.890 164.580 129.150 ;
        RECT 140.560 126.860 143.490 126.880 ;
        RECT 161.350 126.650 164.580 127.890 ;
        RECT 161.350 126.630 164.280 126.650 ;
        RECT 321.560 124.230 321.820 124.900 ;
        RECT 322.565 124.230 322.895 124.845 ;
        RECT 326.235 124.230 326.565 124.695 ;
        RECT 328.445 124.230 328.775 125.160 ;
        RECT 329.755 124.230 330.085 124.795 ;
        RECT 330.615 124.230 330.945 125.255 ;
        RECT 331.650 124.230 332.005 125.270 ;
        RECT 332.570 124.270 332.865 125.350 ;
        RECT 333.830 124.540 334.910 125.240 ;
        RECT 333.830 124.510 334.930 124.540 ;
        RECT 360.860 124.510 370.050 130.660 ;
        RECT 333.820 124.270 334.930 124.510 ;
        RECT 332.570 124.230 334.930 124.270 ;
        RECT 320.990 124.060 334.930 124.230 ;
        RECT 332.700 124.020 334.930 124.060 ;
        RECT 333.820 124.010 334.930 124.020 ;
        RECT 333.820 123.980 334.910 124.010 ;
        RECT 384.620 123.290 384.970 125.450 ;
        RECT 389.980 123.110 390.330 125.270 ;
        RECT 649.750 119.320 658.940 125.510 ;
        RECT 117.420 117.670 121.900 118.820 ;
        RECT 296.400 113.890 302.960 118.430 ;
        RECT 384.580 116.580 384.930 118.740 ;
        RECT 389.710 116.670 390.060 118.830 ;
        RECT 208.020 110.720 210.240 111.180 ;
        RECT 229.470 110.780 231.630 111.130 ;
        RECT 234.170 110.720 236.390 111.180 ;
        RECT 255.620 110.780 257.780 111.130 ;
        RECT 260.320 110.720 262.540 111.180 ;
        RECT 281.770 110.780 283.930 111.130 ;
        RECT 286.470 110.720 288.690 111.180 ;
        RECT 307.920 110.780 310.080 111.130 ;
        RECT 41.650 74.520 45.160 74.530 ;
        RECT 41.650 74.050 45.170 74.520 ;
        RECT 41.650 73.490 45.160 74.050 ;
        RECT 41.650 72.480 42.580 73.490 ;
        RECT 41.660 70.630 42.580 72.480 ;
        RECT 43.660 70.730 44.440 70.900 ;
        RECT 19.400 64.770 20.620 64.820 ;
        RECT 19.340 64.760 20.780 64.770 ;
        RECT 19.340 62.960 26.390 64.760 ;
        RECT 41.670 62.970 42.580 70.630 ;
        RECT 80.510 68.590 81.080 68.600 ;
        RECT 70.780 68.130 81.080 68.590 ;
        RECT 43.750 67.840 44.040 67.900 ;
        RECT 43.700 67.670 44.480 67.840 ;
        RECT 43.750 67.590 44.040 67.670 ;
        RECT 70.800 65.830 71.560 68.130 ;
        RECT 80.510 67.350 81.080 68.130 ;
        RECT 80.510 66.990 81.410 67.350 ;
        RECT 80.580 66.950 81.410 66.990 ;
        RECT 70.800 65.810 74.000 65.830 ;
        RECT 43.680 64.780 44.460 64.950 ;
        RECT 70.770 64.590 74.000 65.810 ;
        RECT 69.400 63.330 74.000 64.590 ;
        RECT 19.340 55.910 20.780 62.960 ;
        RECT 22.710 61.430 23.200 62.960 ;
        RECT 21.550 61.260 24.830 61.430 ;
        RECT 22.710 61.240 23.200 61.260 ;
        RECT 41.710 60.650 42.580 62.970 ;
        RECT 70.770 62.090 74.000 63.330 ;
        RECT 43.720 61.910 44.500 62.080 ;
        RECT 70.770 62.070 73.700 62.090 ;
        RECT 22.530 55.910 22.950 56.100 ;
        RECT 16.750 55.520 18.820 55.840 ;
        RECT 19.340 55.520 26.090 55.910 ;
        RECT 41.670 55.700 42.580 60.650 ;
        RECT 43.720 59.020 44.500 59.190 ;
        RECT 43.720 56.130 44.500 56.300 ;
        RECT 16.750 54.160 26.090 55.520 ;
        RECT 40.960 54.720 42.580 55.700 ;
        RECT 16.750 53.750 18.820 54.160 ;
        RECT 19.290 54.020 26.090 54.160 ;
        RECT 19.290 53.780 20.780 54.020 ;
        RECT 19.290 53.770 19.680 53.780 ;
        RECT 41.710 53.320 42.580 54.720 ;
        RECT 41.710 51.190 42.600 53.320 ;
        RECT 43.740 53.220 44.520 53.390 ;
        RECT 41.710 47.230 42.580 51.190 ;
        RECT 43.720 50.340 44.500 50.510 ;
        RECT 43.700 47.490 44.480 47.660 ;
        RECT 41.720 45.200 42.580 47.230 ;
        RECT 41.720 45.180 44.040 45.200 ;
        RECT 41.730 44.850 44.040 45.180 ;
        RECT 41.730 44.510 45.110 44.850 ;
        RECT 41.730 44.290 45.100 44.510 ;
        RECT 41.730 44.230 45.080 44.290 ;
        RECT 42.970 44.220 44.450 44.230 ;
        RECT 42.970 43.510 43.910 44.220 ;
        RECT 41.760 40.450 44.750 43.510 ;
        RECT 80.900 42.840 81.470 42.850 ;
        RECT 71.170 42.380 81.470 42.840 ;
        RECT 71.190 40.080 71.950 42.380 ;
        RECT 80.900 41.600 81.470 42.380 ;
        RECT 80.900 41.240 81.800 41.600 ;
        RECT 80.970 41.200 81.800 41.240 ;
        RECT 71.190 40.060 74.390 40.080 ;
        RECT 71.160 38.840 74.390 40.060 ;
        RECT 69.790 37.580 74.390 38.840 ;
        RECT 71.160 36.340 74.390 37.580 ;
        RECT 71.160 36.320 74.090 36.340 ;
        RECT 87.620 18.950 87.800 110.215 ;
        RECT 88.195 102.670 88.365 109.710 ;
        RECT 96.400 109.530 96.750 109.740 ;
        RECT 88.195 95.120 88.365 102.160 ;
        RECT 88.195 87.570 88.365 94.610 ;
        RECT 88.195 80.020 88.365 87.060 ;
        RECT 88.195 72.470 88.365 79.510 ;
        RECT 88.195 64.920 88.365 71.960 ;
        RECT 88.195 57.370 88.365 64.410 ;
        RECT 88.195 49.820 88.365 56.860 ;
        RECT 88.195 42.270 88.365 49.310 ;
        RECT 88.195 34.720 88.365 41.760 ;
        RECT 88.195 27.170 88.365 34.210 ;
        RECT 88.195 19.620 88.365 26.660 ;
        RECT 96.440 19.200 96.690 109.530 ;
        RECT 104.775 102.670 104.945 109.710 ;
        RECT 104.775 95.120 104.945 102.160 ;
        RECT 104.775 87.570 104.945 94.610 ;
        RECT 104.775 80.020 104.945 87.060 ;
        RECT 104.775 72.470 104.945 79.510 ;
        RECT 104.775 64.920 104.945 71.960 ;
        RECT 104.775 57.370 104.945 64.410 ;
        RECT 104.775 49.820 104.945 56.860 ;
        RECT 104.775 42.270 104.945 49.310 ;
        RECT 104.775 34.720 104.945 41.760 ;
        RECT 104.775 27.170 104.945 34.210 ;
        RECT 104.775 19.620 104.945 26.660 ;
        RECT 105.340 18.950 105.520 110.210 ;
        RECT 131.490 100.340 132.150 100.820 ;
        RECT 111.885 85.100 112.110 99.785 ;
        RECT 111.760 84.935 112.120 85.100 ;
        RECT 125.235 85.070 125.460 99.785 ;
        RECT 125.090 84.935 125.530 85.070 ;
        RECT 138.550 84.940 138.775 99.790 ;
        RECT 111.760 84.460 112.150 84.935 ;
        RECT 125.090 84.730 125.550 84.935 ;
        RECT 138.550 84.920 138.800 84.940 ;
        RECT 111.760 82.040 112.120 84.460 ;
        RECT 116.285 82.040 116.595 82.280 ;
        RECT 125.090 82.040 125.530 84.730 ;
        RECT 129.630 82.040 129.945 82.280 ;
        RECT 138.390 82.040 138.830 84.920 ;
        RECT 142.950 82.040 143.260 82.280 ;
        RECT 110.375 81.440 150.415 82.040 ;
        RECT 111.760 81.410 112.120 81.440 ;
        RECT 138.390 81.430 138.830 81.440 ;
        RECT 122.650 71.900 123.620 72.510 ;
        RECT 136.160 71.900 136.870 72.530 ;
        RECT 111.885 57.440 112.110 71.070 ;
        RECT 111.880 56.430 112.110 57.440 ;
        RECT 125.235 57.410 125.460 71.070 ;
        RECT 111.880 56.320 112.120 56.430 ;
        RECT 111.760 53.455 112.300 56.320 ;
        RECT 116.285 53.455 116.595 53.560 ;
        RECT 125.010 53.455 125.600 57.410 ;
        RECT 138.550 56.780 138.775 71.070 ;
        RECT 138.520 56.770 138.780 56.780 ;
        RECT 138.390 56.580 139.140 56.770 ;
        RECT 138.380 55.770 139.140 56.580 ;
        RECT 129.630 53.455 129.945 53.560 ;
        RECT 138.410 53.455 139.020 55.770 ;
        RECT 142.950 53.455 143.260 53.560 ;
        RECT 110.465 52.855 150.415 53.455 ;
        RECT 111.760 52.820 112.300 52.855 ;
        RECT 125.010 52.830 125.600 52.855 ;
        RECT 129.630 52.850 129.940 52.855 ;
        RECT 117.890 42.330 118.570 42.970 ;
        RECT 131.140 42.320 132.170 43.060 ;
        RECT 111.885 27.390 112.110 41.680 ;
        RECT 111.790 23.935 112.190 27.390 ;
        RECT 125.235 27.320 125.460 41.680 ;
        RECT 138.550 27.650 138.775 41.685 ;
        RECT 116.285 23.935 116.595 24.170 ;
        RECT 125.190 23.935 125.590 27.320 ;
        RECT 129.630 23.935 129.945 24.170 ;
        RECT 138.440 23.935 138.860 27.650 ;
        RECT 142.950 23.935 143.260 24.170 ;
        RECT 110.465 23.900 150.415 23.935 ;
        RECT 110.450 22.960 150.750 23.900 ;
        RECT 138.440 22.940 138.860 22.960 ;
        RECT 155.725 18.985 155.900 110.215 ;
        RECT 156.300 102.675 156.470 109.715 ;
        RECT 156.300 95.125 156.470 102.165 ;
        RECT 156.300 87.575 156.470 94.615 ;
        RECT 156.300 80.025 156.470 87.065 ;
        RECT 156.300 72.475 156.470 79.515 ;
        RECT 156.300 64.925 156.470 71.965 ;
        RECT 156.300 57.375 156.470 64.415 ;
        RECT 156.300 49.825 156.470 56.865 ;
        RECT 156.300 42.275 156.470 49.315 ;
        RECT 156.300 34.725 156.470 41.765 ;
        RECT 156.300 27.175 156.470 34.215 ;
        RECT 156.300 19.625 156.470 26.665 ;
        RECT 164.560 19.205 164.805 109.720 ;
        RECT 172.880 102.675 173.050 109.715 ;
        RECT 172.880 95.125 173.050 102.165 ;
        RECT 172.880 87.575 173.050 94.615 ;
        RECT 172.880 80.025 173.050 87.065 ;
        RECT 172.880 72.475 173.050 79.515 ;
        RECT 172.880 64.925 173.050 71.965 ;
        RECT 172.880 57.375 173.050 64.415 ;
        RECT 172.880 49.825 173.050 56.865 ;
        RECT 172.880 42.275 173.050 49.315 ;
        RECT 172.880 34.725 173.050 41.765 ;
        RECT 172.880 27.175 173.050 34.215 ;
        RECT 172.880 19.625 173.050 26.665 ;
        RECT 173.445 18.985 173.620 110.215 ;
        RECT 208.020 109.120 210.240 109.580 ;
        RECT 229.470 109.180 231.630 109.530 ;
        RECT 234.170 109.120 236.390 109.580 ;
        RECT 255.620 109.180 257.780 109.530 ;
        RECT 260.320 109.120 262.540 109.580 ;
        RECT 281.770 109.180 283.930 109.530 ;
        RECT 286.470 109.120 288.690 109.580 ;
        RECT 307.920 109.180 310.080 109.530 ;
        RECT 208.020 107.520 210.240 107.980 ;
        RECT 229.470 107.580 231.630 107.930 ;
        RECT 260.260 107.480 262.420 107.830 ;
        RECT 286.470 107.520 288.690 107.980 ;
        RECT 307.920 107.580 310.080 107.930 ;
        RECT 208.020 105.920 210.240 106.380 ;
        RECT 229.470 105.980 231.630 106.330 ;
        RECT 260.260 105.890 262.420 106.240 ;
        RECT 286.470 105.920 288.690 106.380 ;
        RECT 307.920 105.980 310.080 106.330 ;
        RECT 208.020 104.320 210.240 104.780 ;
        RECT 229.470 104.380 231.630 104.730 ;
        RECT 286.470 104.320 288.690 104.780 ;
        RECT 307.920 104.380 310.080 104.730 ;
        RECT 360.860 104.510 370.050 110.660 ;
        RECT 208.020 102.720 210.240 103.180 ;
        RECT 229.470 102.780 231.630 103.130 ;
        RECT 286.470 102.720 288.690 103.180 ;
        RECT 307.920 102.780 310.080 103.130 ;
        RECT 208.020 101.120 210.240 101.580 ;
        RECT 229.470 101.180 231.630 101.530 ;
        RECT 286.470 101.120 288.690 101.580 ;
        RECT 307.920 101.180 310.080 101.530 ;
        RECT 208.020 99.520 210.240 99.980 ;
        RECT 229.470 99.580 231.630 99.930 ;
        RECT 286.470 99.520 288.690 99.980 ;
        RECT 307.920 99.580 310.080 99.930 ;
        RECT 649.750 99.320 658.940 105.510 ;
        RECT 208.020 97.920 210.240 98.380 ;
        RECT 229.470 97.980 231.630 98.330 ;
        RECT 255.690 97.930 257.850 98.280 ;
        RECT 286.470 97.920 288.690 98.380 ;
        RECT 307.920 97.980 310.080 98.330 ;
        RECT 208.020 96.320 210.240 96.780 ;
        RECT 229.470 96.380 231.630 96.730 ;
        RECT 255.690 96.340 257.850 96.690 ;
        RECT 281.670 96.350 283.830 96.700 ;
        RECT 286.470 96.320 288.690 96.780 ;
        RECT 307.920 96.380 310.080 96.730 ;
        RECT 208.020 94.720 210.240 95.180 ;
        RECT 229.470 94.780 231.630 95.130 ;
        RECT 281.670 94.760 283.830 95.110 ;
        RECT 286.470 94.720 288.690 95.180 ;
        RECT 307.920 94.780 310.080 95.130 ;
        RECT 208.020 93.120 210.240 93.580 ;
        RECT 229.470 93.180 231.630 93.530 ;
        RECT 234.340 92.960 236.560 93.420 ;
        RECT 255.790 93.020 257.950 93.370 ;
        RECT 260.320 93.110 262.540 93.570 ;
        RECT 281.770 93.170 283.930 93.520 ;
        RECT 286.470 93.120 288.690 93.580 ;
        RECT 307.920 93.180 310.080 93.530 ;
        RECT 208.020 91.520 210.240 91.980 ;
        RECT 229.470 91.580 231.630 91.930 ;
        RECT 234.340 91.360 236.560 91.820 ;
        RECT 255.790 91.420 257.950 91.770 ;
        RECT 260.320 91.520 262.540 91.980 ;
        RECT 281.770 91.580 283.930 91.930 ;
        RECT 286.470 91.520 288.690 91.980 ;
        RECT 307.920 91.580 310.080 91.930 ;
        RECT 384.580 90.790 384.930 92.950 ;
        RECT 389.710 90.880 390.060 93.040 ;
        RECT 360.860 84.510 370.050 90.660 ;
        RECT 384.690 82.820 385.040 84.980 ;
        RECT 386.280 82.820 386.630 84.980 ;
        RECT 387.870 82.820 388.220 84.980 ;
        RECT 389.460 82.820 389.810 84.980 ;
        RECT 649.750 79.320 658.940 85.510 ;
        RECT 274.470 72.880 275.050 73.050 ;
        RECT 287.460 72.630 288.040 72.800 ;
        RECT 221.010 69.970 221.590 70.140 ;
        RECT 233.680 69.970 234.260 70.140 ;
        RECT 220.570 68.980 220.740 69.580 ;
        RECT 221.860 68.980 222.030 69.580 ;
        RECT 222.950 68.990 223.120 69.590 ;
        RECT 227.810 68.990 227.980 69.590 ;
        RECT 233.240 68.980 233.410 69.580 ;
        RECT 234.530 68.980 234.700 69.580 ;
        RECT 224.020 62.040 230.580 66.580 ;
        RECT 261.130 61.120 267.690 65.660 ;
        RECT 274.030 62.140 274.200 69.240 ;
        RECT 275.320 62.140 275.490 69.240 ;
        RECT 287.020 61.890 287.190 68.990 ;
        RECT 288.310 61.890 288.480 68.990 ;
        RECT 294.290 62.710 300.850 67.250 ;
        RECT 360.860 64.510 370.050 70.660 ;
        RECT 649.750 59.320 658.940 65.510 ;
        RECT 384.690 57.030 385.040 59.190 ;
        RECT 386.280 57.030 386.630 59.190 ;
        RECT 387.870 57.030 388.220 59.190 ;
        RECT 389.460 57.030 389.810 59.190 ;
        RECT 196.700 52.440 197.270 52.450 ;
        RECT 186.970 51.980 197.270 52.440 ;
        RECT 186.990 49.680 187.750 51.980 ;
        RECT 196.700 51.200 197.270 51.980 ;
        RECT 196.700 50.840 197.600 51.200 ;
        RECT 196.770 50.800 197.600 50.840 ;
        RECT 186.990 49.660 190.190 49.680 ;
        RECT 186.960 48.440 190.190 49.660 ;
        RECT 185.590 47.180 190.190 48.440 ;
        RECT 186.960 45.940 190.190 47.180 ;
        RECT 186.960 45.920 189.890 45.940 ;
        RECT 360.860 44.510 370.050 50.660 ;
        RECT 223.740 41.840 225.900 42.190 ;
        RECT 245.150 41.840 247.310 42.190 ;
        RECT 250.560 41.840 252.720 42.190 ;
        RECT 271.970 41.840 274.130 42.190 ;
        RECT 276.260 41.840 278.420 42.190 ;
        RECT 297.670 41.840 299.830 42.190 ;
        RECT 223.740 40.160 225.900 40.510 ;
        RECT 245.150 40.160 247.310 40.510 ;
        RECT 276.260 40.160 278.420 40.510 ;
        RECT 297.670 40.160 299.830 40.510 ;
        RECT 649.750 39.320 658.940 45.510 ;
        RECT 219.040 36.390 221.320 38.750 ;
        RECT 223.740 38.480 225.900 38.830 ;
        RECT 245.150 38.480 247.310 38.830 ;
        RECT 276.260 38.480 278.420 38.830 ;
        RECT 297.670 38.480 299.830 38.830 ;
        RECT 223.930 36.810 226.090 37.160 ;
        RECT 245.340 36.810 247.500 37.160 ;
        RECT 276.450 36.810 278.610 37.160 ;
        RECT 297.860 36.810 300.020 37.160 ;
        RECT 224.030 35.220 226.190 35.570 ;
        RECT 245.440 35.220 247.600 35.570 ;
        RECT 276.550 35.220 278.710 35.570 ;
        RECT 297.960 35.220 300.120 35.570 ;
        RECT 223.880 33.400 226.040 33.750 ;
        RECT 245.290 33.400 247.450 33.750 ;
        RECT 251.000 33.500 253.160 33.850 ;
        RECT 272.410 33.500 274.570 33.850 ;
        RECT 276.690 33.550 278.850 33.900 ;
        RECT 298.100 33.550 300.260 33.900 ;
        RECT 360.860 24.510 370.050 30.660 ;
        RECT 242.710 21.020 244.780 21.720 ;
        RECT 246.440 21.020 248.410 23.180 ;
        RECT 258.150 22.990 258.320 23.070 ;
        RECT 249.300 21.460 249.470 22.780 ;
        RECT 258.140 21.830 258.330 22.990 ;
        RECT 289.300 22.500 289.470 22.580 ;
        RECT 291.880 22.500 292.050 22.580 ;
        RECT 258.150 21.750 258.320 21.830 ;
        RECT 284.080 21.780 284.250 22.240 ;
        RECT 284.080 21.480 284.270 21.780 ;
        RECT 284.080 21.200 284.250 21.480 ;
        RECT 242.710 20.100 248.410 21.020 ;
        RECT 242.710 19.630 244.780 20.100 ;
        RECT 87.580 18.765 105.520 18.950 ;
        RECT 87.580 18.735 105.515 18.765 ;
        RECT 155.720 18.760 173.645 18.985 ;
        RECT 246.440 18.070 248.410 20.100 ;
        RECT 289.290 19.620 289.470 22.500 ;
        RECT 291.870 19.620 292.060 22.500 ;
        RECT 293.800 21.780 293.970 22.840 ;
        RECT 289.300 19.540 289.470 19.620 ;
        RECT 291.880 19.540 292.050 19.620 ;
        RECT 246.420 17.340 248.410 18.070 ;
        RECT 296.350 17.470 298.630 21.540 ;
        RECT 649.750 19.320 658.940 25.510 ;
        RECT 246.400 16.850 248.410 17.340 ;
        RECT 122.890 12.190 123.460 12.200 ;
        RECT 158.270 12.190 158.840 12.200 ;
        RECT 113.160 11.730 123.460 12.190 ;
        RECT 139.800 12.100 140.370 12.110 ;
        RECT 113.180 9.430 113.940 11.730 ;
        RECT 122.890 10.950 123.460 11.730 ;
        RECT 130.070 11.640 140.370 12.100 ;
        RECT 148.540 11.730 158.840 12.190 ;
        RECT 122.890 10.590 123.790 10.950 ;
        RECT 122.960 10.550 123.790 10.590 ;
        RECT 113.180 9.410 116.380 9.430 ;
        RECT 113.150 8.190 116.380 9.410 ;
        RECT 130.090 9.340 130.850 11.640 ;
        RECT 139.800 10.860 140.370 11.640 ;
        RECT 139.800 10.500 140.700 10.860 ;
        RECT 139.870 10.460 140.700 10.500 ;
        RECT 148.560 9.430 149.320 11.730 ;
        RECT 158.270 10.950 158.840 11.730 ;
        RECT 246.400 12.050 248.390 16.850 ;
        RECT 285.010 15.430 298.630 17.470 ;
        RECT 258.230 13.570 258.400 14.180 ;
        RECT 258.170 13.390 258.480 13.570 ;
        RECT 258.230 12.640 258.400 13.390 ;
        RECT 285.030 12.050 287.030 15.430 ;
        RECT 246.400 11.010 287.050 12.050 ;
        RECT 158.270 10.590 159.170 10.950 ;
        RECT 158.340 10.550 159.170 10.590 ;
        RECT 246.420 10.240 287.050 11.010 ;
        RECT 246.420 10.220 283.930 10.240 ;
        RECT 148.560 9.410 151.760 9.430 ;
        RECT 130.090 9.320 133.290 9.340 ;
        RECT 111.780 6.930 116.380 8.190 ;
        RECT 130.060 8.100 133.290 9.320 ;
        RECT 148.530 8.190 151.760 9.410 ;
        RECT 374.170 8.920 383.360 15.150 ;
        RECT 394.170 14.650 395.110 15.130 ;
        RECT 397.810 14.650 403.360 15.130 ;
        RECT 394.170 8.920 403.360 14.650 ;
        RECT 414.170 8.920 423.360 15.130 ;
        RECT 434.170 8.920 443.360 15.130 ;
        RECT 454.170 8.920 463.360 15.130 ;
        RECT 474.170 8.920 483.360 15.130 ;
        RECT 494.170 8.920 503.360 15.130 ;
        RECT 514.170 8.920 523.360 15.130 ;
        RECT 534.170 8.920 543.360 15.130 ;
        RECT 554.170 8.920 563.360 15.130 ;
        RECT 574.170 8.920 583.360 15.130 ;
        RECT 594.170 8.920 603.360 15.130 ;
        RECT 614.170 8.920 623.360 15.130 ;
        RECT 634.170 8.920 643.360 15.130 ;
        RECT 113.150 5.690 116.380 6.930 ;
        RECT 128.690 6.840 133.290 8.100 ;
        RECT 147.160 6.930 151.760 8.190 ;
        RECT 113.150 5.670 116.080 5.690 ;
        RECT 130.060 5.600 133.290 6.840 ;
        RECT 148.530 5.690 151.760 6.930 ;
        RECT 744.490 7.050 771.600 7.220 ;
        RECT 148.530 5.670 151.460 5.690 ;
        RECT 130.060 5.580 132.990 5.600 ;
        RECT 744.490 0.960 744.660 7.050 ;
        RECT 746.350 1.470 746.520 6.680 ;
        RECT 748.930 1.470 749.100 6.680 ;
        RECT 751.510 1.470 751.680 6.680 ;
        RECT 754.090 1.470 754.260 6.680 ;
        RECT 756.670 1.470 756.840 6.680 ;
        RECT 759.250 1.470 759.420 6.680 ;
        RECT 761.830 1.470 762.000 6.680 ;
        RECT 764.410 1.470 764.580 6.680 ;
        RECT 766.990 1.470 767.160 6.680 ;
        RECT 769.570 1.470 769.740 6.680 ;
        RECT 745.055 1.300 771.040 1.470 ;
        RECT 771.430 0.960 771.600 7.050 ;
        RECT 744.490 0.790 771.600 0.960 ;
      LAYER mcon ;
        RECT 739.370 249.770 766.140 249.940 ;
        RECT 739.200 244.290 739.370 249.160 ;
        RECT 741.060 244.440 741.230 249.320 ;
        RECT 743.640 244.440 743.810 249.320 ;
        RECT 746.220 244.440 746.390 249.320 ;
        RECT 748.800 244.440 748.970 249.320 ;
        RECT 751.380 244.440 751.550 249.320 ;
        RECT 753.960 244.440 754.130 249.320 ;
        RECT 756.540 244.440 756.710 249.320 ;
        RECT 759.120 244.440 759.290 249.320 ;
        RECT 761.700 244.440 761.870 249.320 ;
        RECT 764.280 244.440 764.450 249.320 ;
        RECT 766.140 244.290 766.310 249.160 ;
        RECT 740.290 244.020 740.710 244.190 ;
        RECT 741.580 244.020 742.000 244.190 ;
        RECT 742.870 244.020 743.290 244.190 ;
        RECT 744.160 244.020 744.580 244.190 ;
        RECT 745.450 244.020 745.870 244.190 ;
        RECT 746.740 244.020 747.160 244.190 ;
        RECT 748.030 244.020 748.450 244.190 ;
        RECT 749.320 244.020 749.740 244.190 ;
        RECT 750.610 244.020 751.030 244.190 ;
        RECT 751.900 244.020 752.320 244.190 ;
        RECT 753.190 244.020 753.610 244.190 ;
        RECT 754.480 244.020 754.900 244.190 ;
        RECT 755.770 244.020 756.190 244.190 ;
        RECT 757.060 244.020 757.480 244.190 ;
        RECT 758.350 244.020 758.770 244.190 ;
        RECT 759.640 244.020 760.060 244.190 ;
        RECT 760.930 244.020 761.350 244.190 ;
        RECT 762.220 244.020 762.640 244.190 ;
        RECT 763.510 244.020 763.930 244.190 ;
        RECT 764.800 244.020 765.220 244.190 ;
        RECT 370.750 216.540 377.680 220.180 ;
        RECT 390.750 216.540 397.680 220.180 ;
        RECT 410.750 216.540 417.680 220.180 ;
        RECT 430.750 216.540 437.680 220.180 ;
        RECT 450.750 216.540 457.680 220.180 ;
        RECT 470.750 216.540 477.680 220.180 ;
        RECT 490.750 216.540 497.680 220.180 ;
        RECT 510.750 216.540 517.680 220.180 ;
        RECT 530.750 216.540 537.680 220.180 ;
        RECT 550.750 216.540 557.680 220.180 ;
        RECT 570.750 216.540 577.680 220.180 ;
        RECT 590.750 216.540 597.680 220.180 ;
        RECT 610.750 216.540 617.680 220.180 ;
        RECT 630.750 216.540 637.680 220.180 ;
        RECT 650.750 216.540 657.680 220.180 ;
        RECT 362.070 205.720 369.000 209.360 ;
        RECT 650.960 200.530 657.890 204.170 ;
        RECT 362.070 185.720 369.000 189.360 ;
        RECT 384.440 185.555 384.630 187.540 ;
        RECT 386.030 185.555 386.220 187.540 ;
        RECT 387.620 185.555 387.810 187.540 ;
        RECT 389.210 185.555 389.400 187.540 ;
        RECT 650.960 180.530 657.890 184.170 ;
        RECT 362.070 165.720 369.000 169.360 ;
        RECT 384.440 159.770 384.630 161.755 ;
        RECT 386.030 159.770 386.220 161.755 ;
        RECT 387.620 159.770 387.810 161.755 ;
        RECT 389.210 159.770 389.400 161.755 ;
        RECT 650.960 160.530 657.890 164.170 ;
        RECT 168.630 154.940 168.920 155.200 ;
        RECT 170.630 154.940 170.920 155.200 ;
        RECT 362.070 145.720 369.000 149.360 ;
        RECT 384.700 149.165 384.890 151.150 ;
        RECT 390.060 148.985 390.250 150.970 ;
        RECT 650.960 140.530 657.890 144.170 ;
        RECT 129.040 132.295 129.210 132.465 ;
        RECT 150.940 131.855 151.110 132.025 ;
        RECT 117.690 128.810 118.420 129.440 ;
        RECT 171.730 131.625 171.900 131.795 ;
        RECT 309.345 130.125 309.515 130.295 ;
        RECT 309.825 130.125 309.995 130.295 ;
        RECT 310.305 130.125 310.475 130.295 ;
        RECT 310.785 130.125 310.955 130.295 ;
        RECT 311.265 130.125 311.435 130.295 ;
        RECT 311.745 130.125 311.915 130.295 ;
        RECT 312.225 130.125 312.395 130.295 ;
        RECT 312.705 130.125 312.875 130.295 ;
        RECT 313.185 130.125 313.355 130.295 ;
        RECT 313.665 130.125 313.835 130.295 ;
        RECT 314.145 130.125 314.315 130.295 ;
        RECT 314.625 130.125 314.795 130.295 ;
        RECT 315.105 130.125 315.275 130.295 ;
        RECT 315.585 130.125 315.755 130.295 ;
        RECT 316.065 130.125 316.235 130.295 ;
        RECT 316.545 130.125 316.715 130.295 ;
        RECT 317.025 130.125 317.195 130.295 ;
        RECT 317.505 130.125 317.675 130.295 ;
        RECT 317.985 130.125 318.155 130.295 ;
        RECT 318.465 130.125 318.635 130.295 ;
        RECT 318.945 130.125 319.115 130.295 ;
        RECT 319.425 130.125 319.595 130.295 ;
        RECT 319.905 130.125 320.075 130.295 ;
        RECT 320.385 130.125 320.555 130.295 ;
        RECT 320.865 130.125 321.035 130.295 ;
        RECT 323.035 130.160 323.205 130.330 ;
        RECT 323.515 130.160 323.685 130.330 ;
        RECT 323.995 130.160 324.165 130.330 ;
        RECT 324.475 130.160 324.645 130.330 ;
        RECT 324.955 130.160 325.125 130.330 ;
        RECT 325.435 130.160 325.605 130.330 ;
        RECT 325.915 130.160 326.085 130.330 ;
        RECT 326.395 130.160 326.565 130.330 ;
        RECT 326.875 130.160 327.045 130.330 ;
        RECT 327.355 130.160 327.525 130.330 ;
        RECT 327.835 130.160 328.005 130.330 ;
        RECT 328.315 130.160 328.485 130.330 ;
        RECT 328.795 130.160 328.965 130.330 ;
        RECT 329.275 130.160 329.445 130.330 ;
        RECT 329.755 130.160 329.925 130.330 ;
        RECT 330.235 130.160 330.405 130.330 ;
        RECT 330.715 130.160 330.885 130.330 ;
        RECT 331.195 130.160 331.365 130.330 ;
        RECT 331.675 130.160 331.845 130.330 ;
        RECT 332.155 130.160 332.325 130.330 ;
        RECT 332.635 130.160 332.805 130.330 ;
        RECT 333.115 130.160 333.285 130.330 ;
        RECT 333.595 130.160 333.765 130.330 ;
        RECT 334.075 130.160 334.245 130.330 ;
        RECT 334.555 130.160 334.725 130.330 ;
        RECT 139.590 128.370 140.320 129.000 ;
        RECT 160.380 128.140 161.110 128.770 ;
        RECT 362.070 125.720 369.000 129.360 ;
        RECT 321.145 124.060 321.315 124.230 ;
        RECT 321.625 124.060 321.795 124.230 ;
        RECT 322.105 124.060 322.275 124.230 ;
        RECT 322.585 124.060 322.755 124.230 ;
        RECT 323.065 124.060 323.235 124.230 ;
        RECT 323.545 124.060 323.715 124.230 ;
        RECT 324.025 124.060 324.195 124.230 ;
        RECT 324.505 124.060 324.675 124.230 ;
        RECT 324.985 124.060 325.155 124.230 ;
        RECT 325.465 124.060 325.635 124.230 ;
        RECT 325.945 124.060 326.115 124.230 ;
        RECT 326.425 124.060 326.595 124.230 ;
        RECT 326.905 124.060 327.075 124.230 ;
        RECT 327.385 124.060 327.555 124.230 ;
        RECT 327.865 124.060 328.035 124.230 ;
        RECT 328.345 124.060 328.515 124.230 ;
        RECT 328.825 124.060 328.995 124.230 ;
        RECT 329.305 124.060 329.475 124.230 ;
        RECT 329.785 124.060 329.955 124.230 ;
        RECT 330.265 124.060 330.435 124.230 ;
        RECT 330.745 124.060 330.915 124.230 ;
        RECT 331.225 124.060 331.395 124.230 ;
        RECT 331.705 124.060 331.875 124.230 ;
        RECT 332.185 124.060 332.355 124.230 ;
        RECT 332.665 124.060 332.835 124.230 ;
        RECT 384.700 123.380 384.890 125.365 ;
        RECT 390.060 123.200 390.250 125.185 ;
        RECT 650.960 120.530 657.890 124.170 ;
        RECT 297.440 114.990 302.240 117.460 ;
        RECT 384.660 116.665 384.850 118.650 ;
        RECT 389.790 116.755 389.980 118.740 ;
        RECT 208.150 110.860 210.135 111.050 ;
        RECT 229.555 110.860 231.540 111.050 ;
        RECT 234.300 110.860 236.285 111.050 ;
        RECT 255.705 110.860 257.690 111.050 ;
        RECT 260.450 110.860 262.435 111.050 ;
        RECT 281.855 110.860 283.840 111.050 ;
        RECT 286.600 110.860 288.585 111.050 ;
        RECT 308.005 110.860 309.990 111.050 ;
        RECT 43.740 70.730 44.360 70.900 ;
        RECT 43.780 67.670 44.400 67.840 ;
        RECT 81.150 67.065 81.320 67.235 ;
        RECT 43.760 64.780 44.380 64.950 ;
        RECT 69.800 63.580 70.530 64.210 ;
        RECT 43.800 61.910 44.420 62.080 ;
        RECT 17.040 54.000 18.530 55.610 ;
        RECT 43.800 59.020 44.420 59.190 ;
        RECT 43.800 56.130 44.420 56.300 ;
        RECT 43.820 53.220 44.440 53.390 ;
        RECT 43.800 50.340 44.420 50.510 ;
        RECT 43.780 47.490 44.400 47.660 ;
        RECT 42.110 40.810 44.410 43.210 ;
        RECT 81.540 41.315 81.710 41.485 ;
        RECT 70.190 37.830 70.920 38.460 ;
        RECT 88.195 102.750 88.365 109.630 ;
        RECT 96.485 102.750 96.655 109.630 ;
        RECT 88.195 95.200 88.365 102.080 ;
        RECT 104.775 102.750 104.945 109.630 ;
        RECT 96.485 95.200 96.655 102.080 ;
        RECT 88.195 87.650 88.365 94.530 ;
        RECT 104.775 95.200 104.945 102.080 ;
        RECT 96.485 87.650 96.655 94.530 ;
        RECT 88.195 80.100 88.365 86.980 ;
        RECT 104.775 87.650 104.945 94.530 ;
        RECT 96.485 80.100 96.655 86.980 ;
        RECT 88.195 72.550 88.365 79.430 ;
        RECT 104.775 80.100 104.945 86.980 ;
        RECT 96.485 72.550 96.655 79.430 ;
        RECT 88.195 65.000 88.365 71.880 ;
        RECT 104.775 72.550 104.945 79.430 ;
        RECT 96.485 65.000 96.655 71.880 ;
        RECT 88.195 57.450 88.365 64.330 ;
        RECT 104.775 65.000 104.945 71.880 ;
        RECT 96.485 57.450 96.655 64.330 ;
        RECT 88.195 49.900 88.365 56.780 ;
        RECT 104.775 57.450 104.945 64.330 ;
        RECT 96.485 49.900 96.655 56.780 ;
        RECT 88.195 42.350 88.365 49.230 ;
        RECT 104.775 49.900 104.945 56.780 ;
        RECT 96.485 42.350 96.655 49.230 ;
        RECT 88.195 34.800 88.365 41.680 ;
        RECT 104.775 42.350 104.945 49.230 ;
        RECT 96.485 34.800 96.655 41.680 ;
        RECT 88.195 27.250 88.365 34.130 ;
        RECT 104.775 34.800 104.945 41.680 ;
        RECT 96.485 27.250 96.655 34.130 ;
        RECT 88.195 19.700 88.365 26.580 ;
        RECT 104.775 27.250 104.945 34.130 ;
        RECT 96.485 19.700 96.655 26.580 ;
        RECT 104.775 19.700 104.945 26.580 ;
        RECT 116.200 81.470 116.730 82.000 ;
        RECT 129.520 81.470 130.050 82.000 ;
        RECT 142.830 81.470 143.360 82.000 ;
        RECT 116.170 52.875 116.700 53.405 ;
        RECT 129.550 52.910 130.010 53.380 ;
        RECT 142.880 52.910 143.340 53.380 ;
        RECT 116.210 23.430 116.670 23.900 ;
        RECT 129.560 23.430 130.020 23.900 ;
        RECT 142.890 23.430 143.350 23.900 ;
        RECT 156.300 102.755 156.470 109.635 ;
        RECT 164.590 102.755 164.760 109.635 ;
        RECT 156.300 95.205 156.470 102.085 ;
        RECT 172.880 102.755 173.050 109.635 ;
        RECT 164.590 95.205 164.760 102.085 ;
        RECT 156.300 87.655 156.470 94.535 ;
        RECT 172.880 95.205 173.050 102.085 ;
        RECT 164.590 87.655 164.760 94.535 ;
        RECT 156.300 80.105 156.470 86.985 ;
        RECT 172.880 87.655 173.050 94.535 ;
        RECT 164.590 80.105 164.760 86.985 ;
        RECT 156.300 72.555 156.470 79.435 ;
        RECT 172.880 80.105 173.050 86.985 ;
        RECT 164.590 72.555 164.760 79.435 ;
        RECT 156.300 65.005 156.470 71.885 ;
        RECT 172.880 72.555 173.050 79.435 ;
        RECT 164.590 65.005 164.760 71.885 ;
        RECT 156.300 57.455 156.470 64.335 ;
        RECT 172.880 65.005 173.050 71.885 ;
        RECT 164.590 57.455 164.760 64.335 ;
        RECT 156.300 49.905 156.470 56.785 ;
        RECT 172.880 57.455 173.050 64.335 ;
        RECT 164.590 49.905 164.760 56.785 ;
        RECT 156.300 42.355 156.470 49.235 ;
        RECT 172.880 49.905 173.050 56.785 ;
        RECT 164.590 42.355 164.760 49.235 ;
        RECT 156.300 34.805 156.470 41.685 ;
        RECT 172.880 42.355 173.050 49.235 ;
        RECT 164.590 34.805 164.760 41.685 ;
        RECT 156.300 27.255 156.470 34.135 ;
        RECT 172.880 34.805 173.050 41.685 ;
        RECT 164.590 27.255 164.760 34.135 ;
        RECT 156.300 19.705 156.470 26.585 ;
        RECT 172.880 27.255 173.050 34.135 ;
        RECT 164.590 19.705 164.760 26.585 ;
        RECT 172.880 19.705 173.050 26.585 ;
        RECT 208.150 109.260 210.135 109.450 ;
        RECT 229.555 109.260 231.540 109.450 ;
        RECT 234.300 109.260 236.285 109.450 ;
        RECT 255.705 109.260 257.690 109.450 ;
        RECT 260.450 109.260 262.435 109.450 ;
        RECT 281.855 109.260 283.840 109.450 ;
        RECT 286.600 109.260 288.585 109.450 ;
        RECT 308.005 109.260 309.990 109.450 ;
        RECT 208.150 107.660 210.135 107.850 ;
        RECT 229.555 107.660 231.540 107.850 ;
        RECT 260.350 107.560 262.335 107.750 ;
        RECT 286.600 107.660 288.585 107.850 ;
        RECT 308.005 107.660 309.990 107.850 ;
        RECT 208.150 106.060 210.135 106.250 ;
        RECT 229.555 106.060 231.540 106.250 ;
        RECT 260.350 105.970 262.335 106.160 ;
        RECT 286.600 106.060 288.585 106.250 ;
        RECT 308.005 106.060 309.990 106.250 ;
        RECT 362.070 105.720 369.000 109.360 ;
        RECT 208.150 104.460 210.135 104.650 ;
        RECT 229.555 104.460 231.540 104.650 ;
        RECT 286.600 104.460 288.585 104.650 ;
        RECT 308.005 104.460 309.990 104.650 ;
        RECT 208.150 102.860 210.135 103.050 ;
        RECT 229.555 102.860 231.540 103.050 ;
        RECT 286.600 102.860 288.585 103.050 ;
        RECT 308.005 102.860 309.990 103.050 ;
        RECT 208.150 101.260 210.135 101.450 ;
        RECT 229.555 101.260 231.540 101.450 ;
        RECT 286.600 101.260 288.585 101.450 ;
        RECT 308.005 101.260 309.990 101.450 ;
        RECT 650.960 100.530 657.890 104.170 ;
        RECT 208.150 99.660 210.135 99.850 ;
        RECT 229.555 99.660 231.540 99.850 ;
        RECT 286.600 99.660 288.585 99.850 ;
        RECT 308.005 99.660 309.990 99.850 ;
        RECT 208.150 98.060 210.135 98.250 ;
        RECT 229.555 98.060 231.540 98.250 ;
        RECT 255.775 98.010 257.760 98.200 ;
        RECT 286.600 98.060 288.585 98.250 ;
        RECT 308.005 98.060 309.990 98.250 ;
        RECT 208.150 96.460 210.135 96.650 ;
        RECT 229.555 96.460 231.540 96.650 ;
        RECT 255.775 96.420 257.760 96.610 ;
        RECT 281.755 96.430 283.740 96.620 ;
        RECT 286.600 96.460 288.585 96.650 ;
        RECT 308.005 96.460 309.990 96.650 ;
        RECT 208.150 94.860 210.135 95.050 ;
        RECT 229.555 94.860 231.540 95.050 ;
        RECT 281.755 94.840 283.740 95.030 ;
        RECT 286.600 94.860 288.585 95.050 ;
        RECT 308.005 94.860 309.990 95.050 ;
        RECT 208.150 93.260 210.135 93.450 ;
        RECT 229.555 93.260 231.540 93.450 ;
        RECT 234.470 93.100 236.455 93.290 ;
        RECT 255.875 93.100 257.860 93.290 ;
        RECT 260.450 93.250 262.435 93.440 ;
        RECT 281.855 93.250 283.840 93.440 ;
        RECT 286.600 93.260 288.585 93.450 ;
        RECT 308.005 93.260 309.990 93.450 ;
        RECT 208.150 91.660 210.135 91.850 ;
        RECT 229.555 91.660 231.540 91.850 ;
        RECT 234.470 91.500 236.455 91.690 ;
        RECT 255.875 91.500 257.860 91.690 ;
        RECT 260.450 91.660 262.435 91.850 ;
        RECT 281.855 91.660 283.840 91.850 ;
        RECT 286.600 91.660 288.585 91.850 ;
        RECT 308.005 91.660 309.990 91.850 ;
        RECT 384.660 90.880 384.850 92.865 ;
        RECT 389.790 90.970 389.980 92.955 ;
        RECT 362.070 85.720 369.000 89.360 ;
        RECT 384.770 82.905 384.960 84.890 ;
        RECT 386.360 82.905 386.550 84.890 ;
        RECT 387.950 82.905 388.140 84.890 ;
        RECT 389.540 82.905 389.730 84.890 ;
        RECT 650.960 80.530 657.890 84.170 ;
        RECT 274.550 72.880 274.970 73.050 ;
        RECT 287.540 72.630 287.960 72.800 ;
        RECT 221.090 69.970 221.510 70.140 ;
        RECT 233.760 69.970 234.180 70.140 ;
        RECT 220.570 69.060 220.740 69.500 ;
        RECT 221.860 69.060 222.030 69.500 ;
        RECT 222.950 69.070 223.120 69.510 ;
        RECT 227.810 69.070 227.980 69.510 ;
        RECT 233.240 69.060 233.410 69.500 ;
        RECT 234.530 69.060 234.700 69.500 ;
        RECT 225.060 63.140 229.860 65.610 ;
        RECT 262.170 62.220 266.970 64.690 ;
        RECT 274.030 62.220 274.200 69.160 ;
        RECT 275.320 62.220 275.490 69.160 ;
        RECT 287.020 61.970 287.190 68.910 ;
        RECT 288.310 61.970 288.480 68.910 ;
        RECT 295.330 63.810 300.130 66.280 ;
        RECT 362.070 65.720 369.000 69.360 ;
        RECT 650.960 60.530 657.890 64.170 ;
        RECT 384.770 57.120 384.960 59.105 ;
        RECT 386.360 57.120 386.550 59.105 ;
        RECT 387.950 57.120 388.140 59.105 ;
        RECT 389.540 57.120 389.730 59.105 ;
        RECT 197.340 50.915 197.510 51.085 ;
        RECT 185.990 47.430 186.720 48.060 ;
        RECT 362.070 45.720 369.000 49.360 ;
        RECT 223.830 41.920 225.815 42.110 ;
        RECT 245.235 41.920 247.220 42.110 ;
        RECT 250.650 41.920 252.635 42.110 ;
        RECT 272.055 41.920 274.040 42.110 ;
        RECT 276.350 41.920 278.335 42.110 ;
        RECT 297.755 41.920 299.740 42.110 ;
        RECT 650.960 40.530 657.890 44.170 ;
        RECT 223.830 40.240 225.815 40.430 ;
        RECT 245.235 40.240 247.220 40.430 ;
        RECT 276.350 40.240 278.335 40.430 ;
        RECT 297.755 40.240 299.740 40.430 ;
        RECT 219.270 36.590 221.180 38.620 ;
        RECT 223.830 38.560 225.815 38.750 ;
        RECT 245.235 38.560 247.220 38.750 ;
        RECT 276.350 38.560 278.335 38.750 ;
        RECT 297.755 38.560 299.740 38.750 ;
        RECT 224.020 36.890 226.005 37.080 ;
        RECT 245.425 36.890 247.410 37.080 ;
        RECT 276.540 36.890 278.525 37.080 ;
        RECT 297.945 36.890 299.930 37.080 ;
        RECT 224.120 35.300 226.105 35.490 ;
        RECT 245.525 35.300 247.510 35.490 ;
        RECT 276.640 35.300 278.625 35.490 ;
        RECT 298.045 35.300 300.030 35.490 ;
        RECT 223.970 33.480 225.955 33.670 ;
        RECT 245.375 33.480 247.360 33.670 ;
        RECT 251.090 33.580 253.075 33.770 ;
        RECT 272.495 33.580 274.480 33.770 ;
        RECT 276.780 33.630 278.765 33.820 ;
        RECT 298.185 33.630 300.170 33.820 ;
        RECT 362.070 25.720 369.000 29.360 ;
        RECT 242.970 19.940 244.450 21.370 ;
        RECT 249.300 21.540 249.470 22.700 ;
        RECT 258.140 21.830 258.330 22.990 ;
        RECT 284.080 21.280 284.250 22.160 ;
        RECT 289.290 19.620 289.470 22.500 ;
        RECT 291.870 19.620 292.060 22.500 ;
        RECT 293.800 21.860 293.970 22.760 ;
        RECT 650.960 20.530 657.890 24.170 ;
        RECT 123.530 10.665 123.700 10.835 ;
        RECT 140.440 10.575 140.610 10.745 ;
        RECT 258.230 12.720 258.400 14.100 ;
        RECT 158.910 10.665 159.080 10.835 ;
        RECT 375.380 10.130 382.310 13.770 ;
        RECT 395.380 10.130 402.310 13.770 ;
        RECT 415.380 10.130 422.310 13.770 ;
        RECT 435.380 10.130 442.310 13.770 ;
        RECT 455.380 10.130 462.310 13.770 ;
        RECT 475.380 10.130 482.310 13.770 ;
        RECT 495.380 10.130 502.310 13.770 ;
        RECT 515.380 10.130 522.310 13.770 ;
        RECT 535.380 10.130 542.310 13.770 ;
        RECT 555.380 10.130 562.310 13.770 ;
        RECT 575.380 10.130 582.310 13.770 ;
        RECT 595.380 10.130 602.310 13.770 ;
        RECT 615.380 10.130 622.310 13.770 ;
        RECT 635.380 10.130 642.310 13.770 ;
        RECT 112.180 7.180 112.910 7.810 ;
        RECT 129.090 7.090 129.820 7.720 ;
        RECT 147.560 7.180 148.290 7.810 ;
        RECT 744.660 7.050 771.430 7.220 ;
        RECT 744.490 1.570 744.660 6.440 ;
        RECT 746.350 1.720 746.520 6.600 ;
        RECT 748.930 1.720 749.100 6.600 ;
        RECT 751.510 1.720 751.680 6.600 ;
        RECT 754.090 1.720 754.260 6.600 ;
        RECT 756.670 1.720 756.840 6.600 ;
        RECT 759.250 1.720 759.420 6.600 ;
        RECT 761.830 1.720 762.000 6.600 ;
        RECT 764.410 1.720 764.580 6.600 ;
        RECT 766.990 1.720 767.160 6.600 ;
        RECT 769.570 1.720 769.740 6.600 ;
        RECT 771.430 1.570 771.600 6.440 ;
        RECT 745.580 1.300 746.000 1.470 ;
        RECT 746.870 1.300 747.290 1.470 ;
        RECT 748.160 1.300 748.580 1.470 ;
        RECT 749.450 1.300 749.870 1.470 ;
        RECT 750.740 1.300 751.160 1.470 ;
        RECT 752.030 1.300 752.450 1.470 ;
        RECT 753.320 1.300 753.740 1.470 ;
        RECT 754.610 1.300 755.030 1.470 ;
        RECT 755.900 1.300 756.320 1.470 ;
        RECT 757.190 1.300 757.610 1.470 ;
        RECT 758.480 1.300 758.900 1.470 ;
        RECT 759.770 1.300 760.190 1.470 ;
        RECT 761.060 1.300 761.480 1.470 ;
        RECT 762.350 1.300 762.770 1.470 ;
        RECT 763.640 1.300 764.060 1.470 ;
        RECT 764.930 1.300 765.350 1.470 ;
        RECT 766.220 1.300 766.640 1.470 ;
        RECT 767.510 1.300 767.930 1.470 ;
        RECT 768.800 1.300 769.220 1.470 ;
        RECT 770.090 1.300 770.510 1.470 ;
      LAYER met1 ;
        RECT 739.170 249.570 766.340 251.075 ;
        RECT 739.170 244.230 739.400 249.570 ;
        RECT 741.060 249.380 741.230 249.570 ;
        RECT 743.640 249.380 743.810 249.570 ;
        RECT 746.220 249.380 746.390 249.570 ;
        RECT 748.800 249.380 748.970 249.570 ;
        RECT 751.380 249.380 751.550 249.570 ;
        RECT 753.960 249.380 754.130 249.570 ;
        RECT 756.540 249.380 756.710 249.570 ;
        RECT 759.120 249.380 759.290 249.570 ;
        RECT 761.700 249.380 761.870 249.570 ;
        RECT 764.280 249.380 764.450 249.570 ;
        RECT 741.030 244.380 741.260 249.380 ;
        RECT 743.610 244.380 743.840 249.380 ;
        RECT 746.190 244.380 746.420 249.380 ;
        RECT 748.770 244.380 749.000 249.380 ;
        RECT 751.350 244.380 751.580 249.380 ;
        RECT 753.930 244.380 754.160 249.380 ;
        RECT 756.510 244.380 756.740 249.380 ;
        RECT 759.090 244.380 759.320 249.380 ;
        RECT 761.670 244.380 761.900 249.380 ;
        RECT 764.250 244.380 764.480 249.380 ;
        RECT 766.110 244.230 766.340 249.570 ;
        RECT 740.230 243.990 740.770 244.220 ;
        RECT 741.520 243.990 742.060 244.220 ;
        RECT 742.810 243.990 743.350 244.220 ;
        RECT 744.100 243.990 744.640 244.220 ;
        RECT 745.390 243.990 745.930 244.220 ;
        RECT 746.680 243.990 747.220 244.220 ;
        RECT 747.970 243.990 748.510 244.220 ;
        RECT 749.260 243.990 749.800 244.220 ;
        RECT 750.550 243.990 751.090 244.220 ;
        RECT 751.840 243.990 752.380 244.220 ;
        RECT 753.130 243.990 753.670 244.220 ;
        RECT 754.420 243.990 754.960 244.220 ;
        RECT 755.710 243.990 756.250 244.220 ;
        RECT 757.000 243.990 757.540 244.220 ;
        RECT 758.290 243.990 758.830 244.220 ;
        RECT 759.580 243.990 760.120 244.220 ;
        RECT 760.870 243.990 761.410 244.220 ;
        RECT 762.160 243.990 762.700 244.220 ;
        RECT 763.450 243.990 763.990 244.220 ;
        RECT 764.740 243.990 765.280 244.220 ;
        RECT 369.540 215.330 378.730 221.480 ;
        RECT 389.540 215.330 398.730 221.480 ;
        RECT 409.540 215.330 418.730 221.480 ;
        RECT 429.540 215.330 438.730 221.480 ;
        RECT 449.540 215.330 458.730 221.480 ;
        RECT 469.540 215.330 478.730 221.480 ;
        RECT 489.540 215.330 498.730 221.480 ;
        RECT 509.540 215.330 518.730 221.480 ;
        RECT 529.540 215.330 538.730 221.480 ;
        RECT 549.540 215.330 558.730 221.480 ;
        RECT 569.540 215.330 578.730 221.480 ;
        RECT 589.540 215.330 598.730 221.480 ;
        RECT 609.540 215.330 618.730 221.480 ;
        RECT 629.540 215.330 638.730 221.480 ;
        RECT 649.540 215.330 658.730 221.480 ;
        RECT 360.860 204.510 370.050 210.660 ;
        RECT 649.750 199.320 658.940 205.510 ;
        RECT 360.860 184.510 370.050 190.660 ;
        RECT 384.260 185.380 389.600 187.710 ;
        RECT 649.750 179.320 658.940 185.510 ;
        RECT 360.860 164.510 370.050 170.660 ;
        RECT 384.250 159.550 389.590 161.880 ;
        RECT 649.750 159.320 658.940 165.510 ;
        RECT 168.470 154.870 171.490 155.280 ;
        RECT 360.860 144.510 370.050 150.660 ;
        RECT 384.540 149.020 385.070 151.310 ;
        RECT 389.880 148.850 390.410 151.140 ;
        RECT 649.750 139.320 658.940 145.510 ;
        RECT 128.980 132.220 129.260 132.540 ;
        RECT 150.880 131.780 151.160 132.100 ;
        RECT 171.670 131.550 171.950 131.870 ;
        RECT 322.270 130.490 323.390 130.510 ;
        RECT 309.190 130.380 321.190 130.455 ;
        RECT 322.270 130.380 334.880 130.490 ;
        RECT 309.190 130.040 334.880 130.380 ;
        RECT 309.190 129.965 321.190 130.040 ;
        RECT 322.270 130.000 334.880 130.040 ;
        RECT 322.270 129.970 323.390 130.000 ;
        RECT 117.550 128.690 118.530 129.590 ;
        RECT 139.450 128.250 140.430 129.150 ;
        RECT 160.240 128.020 161.220 128.920 ;
        RECT 318.820 124.290 319.140 129.965 ;
        RECT 348.190 126.270 349.790 126.360 ;
        RECT 357.440 126.320 370.220 130.860 ;
        RECT 354.560 126.270 370.220 126.320 ;
        RECT 348.190 125.950 370.220 126.270 ;
        RECT 348.190 125.460 349.790 125.950 ;
        RECT 354.560 125.920 370.220 125.950 ;
        RECT 337.240 124.560 337.890 124.840 ;
        RECT 332.610 124.390 337.910 124.560 ;
        RECT 357.440 124.510 370.220 125.920 ;
        RECT 320.990 124.290 337.910 124.390 ;
        RECT 318.820 124.000 337.910 124.290 ;
        RECT 318.820 123.900 332.990 124.000 ;
        RECT 318.820 123.810 321.330 123.900 ;
        RECT 337.240 123.740 337.890 124.000 ;
        RECT 384.540 123.220 385.070 125.510 ;
        RECT 389.890 123.030 390.420 125.320 ;
        RECT 649.750 119.320 658.940 125.510 ;
        RECT 296.400 113.890 302.960 118.430 ;
        RECT 384.470 116.510 385.030 118.810 ;
        RECT 389.570 116.560 390.180 118.890 ;
        RECT 207.440 111.540 286.570 111.700 ;
        RECT 298.030 111.540 298.330 113.890 ;
        RECT 43.680 70.650 44.420 70.960 ;
        RECT 43.720 67.590 44.460 67.900 ;
        RECT 81.090 66.990 81.370 67.310 ;
        RECT 43.670 64.700 44.450 65.010 ;
        RECT 69.660 63.460 70.640 64.360 ;
        RECT 43.740 61.830 44.480 62.140 ;
        RECT 43.740 58.940 44.480 59.250 ;
        RECT 43.740 56.050 44.480 56.360 ;
        RECT 16.750 53.750 18.820 55.840 ;
        RECT 43.760 53.140 44.500 53.450 ;
        RECT 43.740 50.260 44.480 50.570 ;
        RECT 43.720 47.410 44.460 47.720 ;
        RECT 43.250 43.510 43.700 44.070 ;
        RECT 41.760 40.450 44.750 43.510 ;
        RECT 81.480 41.240 81.760 41.560 ;
        RECT 70.050 37.710 71.030 38.610 ;
        RECT 87.430 18.565 105.710 110.275 ;
        RECT 116.100 81.420 116.820 82.040 ;
        RECT 129.430 81.420 130.150 82.040 ;
        RECT 142.735 81.415 143.465 82.040 ;
        RECT 116.060 52.820 116.830 53.455 ;
        RECT 129.480 52.850 130.105 53.460 ;
        RECT 142.800 52.850 143.425 53.480 ;
        RECT 116.010 23.230 117.180 24.030 ;
        RECT 129.430 23.365 130.165 23.980 ;
        RECT 142.770 23.355 143.505 23.970 ;
        RECT 155.520 18.585 173.805 110.255 ;
        RECT 207.440 108.620 310.590 111.540 ;
        RECT 207.440 94.170 232.460 108.620 ;
        RECT 260.200 105.810 262.450 107.890 ;
        RECT 255.670 96.280 257.900 98.370 ;
        RECT 281.630 94.680 283.910 96.770 ;
        RECT 285.570 94.170 310.590 108.620 ;
        RECT 360.860 104.510 370.050 110.660 ;
        RECT 649.750 99.320 658.940 105.510 ;
        RECT 207.440 91.160 310.590 94.170 ;
        RECT 230.330 91.010 310.590 91.160 ;
        RECT 285.570 91.000 310.590 91.010 ;
        RECT 360.860 84.510 370.050 90.660 ;
        RECT 384.440 90.640 385.070 93.070 ;
        RECT 389.600 90.740 390.230 93.150 ;
        RECT 384.420 82.680 390.040 85.250 ;
        RECT 649.750 79.320 658.940 85.510 ;
        RECT 220.460 68.610 222.120 70.310 ;
        RECT 222.880 69.570 228.050 69.660 ;
        RECT 222.880 68.960 228.110 69.570 ;
        RECT 221.120 68.370 221.370 68.610 ;
        RECT 227.720 68.370 228.110 68.960 ;
        RECT 233.210 68.570 234.870 70.270 ;
        RECT 233.780 68.370 234.030 68.570 ;
        RECT 221.090 68.190 234.030 68.370 ;
        RECT 221.090 68.110 234.000 68.190 ;
        RECT 227.390 66.580 227.600 68.110 ;
        RECT 224.020 62.040 230.580 66.580 ;
        RECT 261.130 61.120 267.690 65.660 ;
        RECT 273.740 61.190 275.800 73.420 ;
        RECT 286.690 65.170 288.750 73.250 ;
        RECT 294.290 65.170 300.850 67.250 ;
        RECT 286.690 63.590 300.850 65.170 ;
        RECT 360.860 64.510 370.050 70.660 ;
        RECT 286.690 61.190 288.750 63.590 ;
        RECT 294.290 62.710 300.850 63.590 ;
        RECT 273.740 60.870 288.750 61.190 ;
        RECT 273.740 58.300 275.800 60.870 ;
        RECT 286.690 58.130 288.750 60.870 ;
        RECT 384.370 56.770 390.440 59.390 ;
        RECT 649.750 59.320 658.940 65.510 ;
        RECT 197.280 50.840 197.560 51.160 ;
        RECT 185.850 47.310 186.830 48.210 ;
        RECT 360.860 44.510 370.050 50.660 ;
        RECT 217.760 43.470 221.670 43.590 ;
        RECT 217.760 43.420 247.840 43.470 ;
        RECT 276.810 43.420 300.930 43.450 ;
        RECT 217.760 42.850 300.930 43.420 ;
        RECT 217.760 41.590 300.880 42.850 ;
        RECT 217.760 40.110 247.840 41.590 ;
        RECT 217.610 35.960 247.840 40.110 ;
        RECT 217.610 35.410 247.940 35.960 ;
        RECT 217.760 34.280 247.940 35.410 ;
        RECT 275.700 34.680 300.880 41.590 ;
        RECT 649.750 39.320 658.940 45.510 ;
        RECT 275.800 34.280 300.880 34.680 ;
        RECT 217.760 33.020 300.880 34.280 ;
        RECT 221.310 33.010 300.880 33.020 ;
        RECT 221.310 33.000 275.660 33.010 ;
        RECT 239.580 21.420 240.710 33.000 ;
        RECT 278.420 32.970 299.590 33.010 ;
        RECT 360.860 24.510 370.050 30.660 ;
        RECT 249.210 22.740 249.530 22.770 ;
        RECT 242.710 21.420 244.780 21.720 ;
        RECT 249.210 21.480 249.570 22.740 ;
        RECT 258.090 21.770 258.380 23.060 ;
        RECT 293.710 22.820 294.020 22.830 ;
        RECT 289.240 22.550 289.520 22.560 ;
        RECT 239.460 19.850 244.780 21.420 ;
        RECT 283.970 21.210 284.320 22.230 ;
        RECT 239.580 19.790 240.710 19.850 ;
        RECT 242.710 19.630 244.780 19.850 ;
        RECT 289.240 19.550 289.530 22.550 ;
        RECT 291.830 19.550 292.100 22.560 ;
        RECT 293.710 21.800 294.030 22.820 ;
        RECT 293.710 21.780 294.020 21.800 ;
        RECT 289.270 18.680 289.460 19.550 ;
        RECT 291.870 19.490 292.070 19.550 ;
        RECT 291.880 18.680 292.060 19.490 ;
        RECT 649.750 19.320 658.940 25.510 ;
        RECT 289.270 18.450 292.070 18.680 ;
        RECT 258.130 12.660 258.460 14.150 ;
        RECT 258.160 12.650 258.460 12.660 ;
        RECT 123.470 10.590 123.750 10.910 ;
        RECT 140.380 10.500 140.660 10.820 ;
        RECT 158.850 10.590 159.130 10.910 ;
        RECT 374.170 8.920 383.360 15.150 ;
        RECT 394.170 14.650 395.110 15.130 ;
        RECT 397.810 14.650 403.360 15.130 ;
        RECT 394.170 8.920 403.360 14.650 ;
        RECT 414.170 8.920 423.360 15.130 ;
        RECT 434.170 8.920 443.360 15.130 ;
        RECT 454.170 8.920 463.360 15.130 ;
        RECT 474.170 8.920 483.360 15.130 ;
        RECT 494.170 8.920 503.360 15.130 ;
        RECT 514.170 8.920 523.360 15.130 ;
        RECT 534.170 8.920 543.360 15.130 ;
        RECT 554.170 8.920 563.360 15.130 ;
        RECT 574.170 8.920 583.360 15.130 ;
        RECT 594.170 8.920 603.360 15.130 ;
        RECT 614.170 8.920 623.360 15.130 ;
        RECT 634.170 8.920 643.360 15.130 ;
        RECT 112.040 7.060 113.020 7.960 ;
        RECT 128.950 6.970 129.930 7.870 ;
        RECT 147.420 7.060 148.400 7.960 ;
        RECT 744.460 6.850 771.630 8.355 ;
        RECT 744.460 1.510 744.690 6.850 ;
        RECT 746.350 6.660 746.520 6.850 ;
        RECT 748.930 6.660 749.100 6.850 ;
        RECT 751.510 6.660 751.680 6.850 ;
        RECT 754.090 6.660 754.260 6.850 ;
        RECT 756.670 6.660 756.840 6.850 ;
        RECT 759.250 6.660 759.420 6.850 ;
        RECT 761.830 6.660 762.000 6.850 ;
        RECT 764.410 6.660 764.580 6.850 ;
        RECT 766.990 6.660 767.160 6.850 ;
        RECT 769.570 6.660 769.740 6.850 ;
        RECT 746.320 1.660 746.550 6.660 ;
        RECT 748.900 1.660 749.130 6.660 ;
        RECT 751.480 1.660 751.710 6.660 ;
        RECT 754.060 1.660 754.290 6.660 ;
        RECT 756.640 1.660 756.870 6.660 ;
        RECT 759.220 1.660 759.450 6.660 ;
        RECT 761.800 1.660 762.030 6.660 ;
        RECT 764.380 1.660 764.610 6.660 ;
        RECT 766.960 1.660 767.190 6.660 ;
        RECT 769.540 1.660 769.770 6.660 ;
        RECT 771.400 1.510 771.630 6.850 ;
        RECT 745.520 1.270 746.060 1.500 ;
        RECT 746.810 1.270 747.350 1.500 ;
        RECT 748.100 1.270 748.640 1.500 ;
        RECT 749.390 1.270 749.930 1.500 ;
        RECT 750.680 1.270 751.220 1.500 ;
        RECT 751.970 1.270 752.510 1.500 ;
        RECT 753.260 1.270 753.800 1.500 ;
        RECT 754.550 1.270 755.090 1.500 ;
        RECT 755.840 1.270 756.380 1.500 ;
        RECT 757.130 1.270 757.670 1.500 ;
        RECT 758.420 1.270 758.960 1.500 ;
        RECT 759.710 1.270 760.250 1.500 ;
        RECT 761.000 1.270 761.540 1.500 ;
        RECT 762.290 1.270 762.830 1.500 ;
        RECT 763.580 1.270 764.120 1.500 ;
        RECT 764.870 1.270 765.410 1.500 ;
        RECT 766.160 1.270 766.700 1.500 ;
        RECT 767.450 1.270 767.990 1.500 ;
        RECT 768.740 1.270 769.280 1.500 ;
        RECT 770.030 1.270 770.570 1.500 ;
      LAYER via ;
        RECT 740.820 250.510 741.220 250.910 ;
        RECT 741.620 250.510 742.020 250.910 ;
        RECT 742.420 250.510 742.820 250.910 ;
        RECT 743.220 250.510 743.620 250.910 ;
        RECT 744.020 250.510 744.420 250.910 ;
        RECT 744.820 250.510 745.220 250.910 ;
        RECT 745.620 250.510 746.020 250.910 ;
        RECT 746.420 250.510 746.820 250.910 ;
        RECT 747.220 250.510 747.620 250.910 ;
        RECT 748.020 250.510 748.420 250.910 ;
        RECT 748.820 250.510 749.220 250.910 ;
        RECT 749.620 250.510 750.020 250.910 ;
        RECT 750.420 250.510 750.820 250.910 ;
        RECT 751.220 250.510 751.620 250.910 ;
        RECT 752.020 250.510 752.420 250.910 ;
        RECT 752.820 250.510 753.220 250.910 ;
        RECT 753.620 250.510 754.020 250.910 ;
        RECT 754.420 250.510 754.820 250.910 ;
        RECT 755.220 250.510 755.620 250.910 ;
        RECT 756.020 250.510 756.420 250.910 ;
        RECT 756.820 250.510 757.220 250.910 ;
        RECT 757.620 250.510 758.020 250.910 ;
        RECT 758.420 250.510 758.820 250.910 ;
        RECT 759.220 250.510 759.620 250.910 ;
        RECT 760.020 250.510 760.420 250.910 ;
        RECT 760.820 250.510 761.220 250.910 ;
        RECT 761.620 250.510 762.020 250.910 ;
        RECT 762.420 250.510 762.820 250.910 ;
        RECT 763.220 250.510 763.620 250.910 ;
        RECT 764.020 250.510 764.420 250.910 ;
        RECT 764.820 250.510 765.220 250.910 ;
        RECT 740.820 249.710 741.220 250.110 ;
        RECT 741.620 249.710 742.020 250.110 ;
        RECT 742.420 249.710 742.820 250.110 ;
        RECT 743.220 249.710 743.620 250.110 ;
        RECT 744.020 249.710 744.420 250.110 ;
        RECT 744.820 249.710 745.220 250.110 ;
        RECT 745.620 249.710 746.020 250.110 ;
        RECT 746.420 249.710 746.820 250.110 ;
        RECT 747.220 249.710 747.620 250.110 ;
        RECT 748.020 249.710 748.420 250.110 ;
        RECT 748.820 249.710 749.220 250.110 ;
        RECT 749.620 249.710 750.020 250.110 ;
        RECT 750.420 249.710 750.820 250.110 ;
        RECT 751.220 249.710 751.620 250.110 ;
        RECT 752.020 249.710 752.420 250.110 ;
        RECT 752.820 249.710 753.220 250.110 ;
        RECT 753.620 249.710 754.020 250.110 ;
        RECT 754.420 249.710 754.820 250.110 ;
        RECT 755.220 249.710 755.620 250.110 ;
        RECT 756.020 249.710 756.420 250.110 ;
        RECT 756.820 249.710 757.220 250.110 ;
        RECT 757.620 249.710 758.020 250.110 ;
        RECT 758.420 249.710 758.820 250.110 ;
        RECT 759.220 249.710 759.620 250.110 ;
        RECT 760.020 249.710 760.420 250.110 ;
        RECT 760.820 249.710 761.220 250.110 ;
        RECT 761.620 249.710 762.020 250.110 ;
        RECT 762.420 249.710 762.820 250.110 ;
        RECT 763.220 249.710 763.620 250.110 ;
        RECT 764.020 249.710 764.420 250.110 ;
        RECT 764.820 249.710 765.220 250.110 ;
        RECT 370.750 216.540 377.680 220.180 ;
        RECT 390.750 216.540 397.680 220.180 ;
        RECT 410.750 216.540 417.680 220.180 ;
        RECT 430.750 216.540 437.680 220.180 ;
        RECT 450.750 216.540 457.680 220.180 ;
        RECT 470.750 216.540 477.680 220.180 ;
        RECT 490.750 216.540 497.680 220.180 ;
        RECT 510.750 216.540 517.680 220.180 ;
        RECT 530.750 216.540 537.680 220.180 ;
        RECT 550.750 216.540 557.680 220.180 ;
        RECT 570.750 216.540 577.680 220.180 ;
        RECT 590.750 216.540 597.680 220.180 ;
        RECT 610.750 216.540 617.680 220.180 ;
        RECT 630.750 216.540 637.680 220.180 ;
        RECT 650.750 216.540 657.680 220.180 ;
        RECT 362.070 205.720 369.000 209.360 ;
        RECT 650.960 200.530 657.890 204.170 ;
        RECT 362.070 185.720 369.000 189.360 ;
        RECT 384.340 185.470 384.720 187.650 ;
        RECT 385.940 185.470 386.320 187.650 ;
        RECT 387.520 185.470 387.900 187.650 ;
        RECT 389.120 185.470 389.500 187.650 ;
        RECT 650.960 180.530 657.890 184.170 ;
        RECT 362.070 165.720 369.000 169.360 ;
        RECT 384.360 159.680 384.720 161.840 ;
        RECT 385.940 159.680 386.300 161.840 ;
        RECT 387.540 159.680 387.900 161.840 ;
        RECT 389.120 159.680 389.480 161.840 ;
        RECT 650.960 160.530 657.890 164.170 ;
        RECT 168.630 154.940 168.920 155.200 ;
        RECT 170.630 154.940 170.920 155.200 ;
        RECT 362.070 145.720 369.000 149.360 ;
        RECT 384.620 149.070 384.980 151.230 ;
        RECT 389.970 148.930 390.330 151.090 ;
        RECT 650.960 140.530 657.890 144.170 ;
        RECT 117.690 128.810 118.420 129.440 ;
        RECT 139.590 128.370 140.320 129.000 ;
        RECT 160.380 128.140 161.110 128.770 ;
        RECT 348.710 125.740 349.300 126.000 ;
        RECT 362.070 125.720 369.000 129.360 ;
        RECT 337.420 124.020 337.770 124.510 ;
        RECT 384.610 123.290 384.980 125.450 ;
        RECT 389.970 123.090 390.340 125.250 ;
        RECT 650.960 120.530 657.890 124.170 ;
        RECT 297.440 114.990 302.240 117.460 ;
        RECT 384.570 116.610 384.940 118.770 ;
        RECT 389.690 116.660 390.060 118.820 ;
        RECT 116.200 81.470 116.730 82.000 ;
        RECT 129.520 81.470 130.050 82.000 ;
        RECT 142.830 81.470 143.360 82.000 ;
        RECT 95.820 78.480 97.480 80.650 ;
        RECT 43.720 70.650 44.390 70.960 ;
        RECT 43.760 67.590 44.430 67.900 ;
        RECT 43.740 64.700 44.410 65.010 ;
        RECT 69.800 63.580 70.530 64.210 ;
        RECT 43.780 61.830 44.450 62.140 ;
        RECT 43.780 58.940 44.450 59.250 ;
        RECT 43.780 56.050 44.450 56.360 ;
        RECT 17.040 54.000 18.530 55.610 ;
        RECT 43.800 53.140 44.470 53.450 ;
        RECT 43.780 50.260 44.450 50.570 ;
        RECT 43.760 47.410 44.430 47.720 ;
        RECT 42.110 40.810 44.410 43.210 ;
        RECT 70.190 37.830 70.920 38.460 ;
        RECT 260.260 107.470 262.430 107.840 ;
        RECT 260.260 105.870 262.430 106.240 ;
        RECT 255.690 97.920 257.850 98.280 ;
        RECT 255.690 96.340 257.850 96.700 ;
        RECT 281.670 96.350 283.850 96.700 ;
        RECT 281.670 94.760 283.850 95.110 ;
        RECT 362.070 105.720 369.000 109.360 ;
        RECT 650.960 100.530 657.890 104.170 ;
        RECT 384.580 90.780 384.930 92.950 ;
        RECT 389.710 90.880 390.060 93.050 ;
        RECT 362.070 85.720 369.000 89.360 ;
        RECT 384.680 82.820 385.040 85.010 ;
        RECT 386.310 82.820 386.670 85.010 ;
        RECT 387.870 82.840 388.230 85.030 ;
        RECT 389.460 82.800 389.820 84.990 ;
        RECT 162.210 77.870 167.210 80.850 ;
        RECT 650.960 80.530 657.890 84.170 ;
        RECT 116.170 52.875 116.700 53.405 ;
        RECT 129.550 52.910 130.010 53.380 ;
        RECT 142.880 52.910 143.340 53.380 ;
        RECT 116.210 23.430 116.670 23.900 ;
        RECT 129.560 23.430 130.020 23.900 ;
        RECT 142.890 23.430 143.350 23.900 ;
        RECT 225.060 63.140 229.860 65.610 ;
        RECT 262.170 62.220 266.970 64.690 ;
        RECT 295.330 63.810 300.130 66.280 ;
        RECT 362.070 65.720 369.000 69.360 ;
        RECT 650.960 60.530 657.890 64.170 ;
        RECT 384.680 57.000 385.040 59.190 ;
        RECT 386.260 57.000 386.620 59.190 ;
        RECT 387.880 57.000 388.240 59.190 ;
        RECT 389.460 57.180 389.820 59.220 ;
        RECT 185.990 47.430 186.720 48.060 ;
        RECT 362.070 45.720 369.000 49.360 ;
        RECT 219.300 36.600 221.140 38.590 ;
        RECT 650.960 40.530 657.890 44.170 ;
        RECT 362.070 25.720 369.000 29.360 ;
        RECT 249.240 21.540 249.520 22.700 ;
        RECT 258.090 21.830 258.370 22.990 ;
        RECT 242.970 19.940 244.450 21.370 ;
        RECT 284.030 21.280 284.310 22.160 ;
        RECT 289.240 19.610 289.510 22.500 ;
        RECT 293.740 21.860 294.020 22.760 ;
        RECT 650.960 20.530 657.890 24.170 ;
        RECT 258.170 12.720 258.460 14.110 ;
        RECT 375.380 10.130 382.310 13.770 ;
        RECT 395.380 10.130 402.310 13.770 ;
        RECT 415.380 10.130 422.310 13.770 ;
        RECT 435.380 10.130 442.310 13.770 ;
        RECT 455.380 10.130 462.310 13.770 ;
        RECT 475.380 10.130 482.310 13.770 ;
        RECT 495.380 10.130 502.310 13.770 ;
        RECT 515.380 10.130 522.310 13.770 ;
        RECT 535.380 10.130 542.310 13.770 ;
        RECT 555.380 10.130 562.310 13.770 ;
        RECT 575.380 10.130 582.310 13.770 ;
        RECT 595.380 10.130 602.310 13.770 ;
        RECT 615.380 10.130 622.310 13.770 ;
        RECT 635.380 10.130 642.310 13.770 ;
        RECT 112.180 7.180 112.910 7.810 ;
        RECT 129.090 7.090 129.820 7.720 ;
        RECT 147.560 7.180 148.290 7.810 ;
        RECT 746.110 7.790 746.510 8.190 ;
        RECT 746.910 7.790 747.310 8.190 ;
        RECT 747.710 7.790 748.110 8.190 ;
        RECT 748.510 7.790 748.910 8.190 ;
        RECT 749.310 7.790 749.710 8.190 ;
        RECT 750.110 7.790 750.510 8.190 ;
        RECT 750.910 7.790 751.310 8.190 ;
        RECT 751.710 7.790 752.110 8.190 ;
        RECT 752.510 7.790 752.910 8.190 ;
        RECT 753.310 7.790 753.710 8.190 ;
        RECT 754.110 7.790 754.510 8.190 ;
        RECT 754.910 7.790 755.310 8.190 ;
        RECT 755.710 7.790 756.110 8.190 ;
        RECT 756.510 7.790 756.910 8.190 ;
        RECT 757.310 7.790 757.710 8.190 ;
        RECT 758.110 7.790 758.510 8.190 ;
        RECT 758.910 7.790 759.310 8.190 ;
        RECT 759.710 7.790 760.110 8.190 ;
        RECT 760.510 7.790 760.910 8.190 ;
        RECT 761.310 7.790 761.710 8.190 ;
        RECT 762.110 7.790 762.510 8.190 ;
        RECT 762.910 7.790 763.310 8.190 ;
        RECT 763.710 7.790 764.110 8.190 ;
        RECT 764.510 7.790 764.910 8.190 ;
        RECT 765.310 7.790 765.710 8.190 ;
        RECT 766.110 7.790 766.510 8.190 ;
        RECT 766.910 7.790 767.310 8.190 ;
        RECT 767.710 7.790 768.110 8.190 ;
        RECT 768.510 7.790 768.910 8.190 ;
        RECT 769.310 7.790 769.710 8.190 ;
        RECT 770.110 7.790 770.510 8.190 ;
        RECT 746.110 6.990 746.510 7.390 ;
        RECT 746.910 6.990 747.310 7.390 ;
        RECT 747.710 6.990 748.110 7.390 ;
        RECT 748.510 6.990 748.910 7.390 ;
        RECT 749.310 6.990 749.710 7.390 ;
        RECT 750.110 6.990 750.510 7.390 ;
        RECT 750.910 6.990 751.310 7.390 ;
        RECT 751.710 6.990 752.110 7.390 ;
        RECT 752.510 6.990 752.910 7.390 ;
        RECT 753.310 6.990 753.710 7.390 ;
        RECT 754.110 6.990 754.510 7.390 ;
        RECT 754.910 6.990 755.310 7.390 ;
        RECT 755.710 6.990 756.110 7.390 ;
        RECT 756.510 6.990 756.910 7.390 ;
        RECT 757.310 6.990 757.710 7.390 ;
        RECT 758.110 6.990 758.510 7.390 ;
        RECT 758.910 6.990 759.310 7.390 ;
        RECT 759.710 6.990 760.110 7.390 ;
        RECT 760.510 6.990 760.910 7.390 ;
        RECT 761.310 6.990 761.710 7.390 ;
        RECT 762.110 6.990 762.510 7.390 ;
        RECT 762.910 6.990 763.310 7.390 ;
        RECT 763.710 6.990 764.110 7.390 ;
        RECT 764.510 6.990 764.910 7.390 ;
        RECT 765.310 6.990 765.710 7.390 ;
        RECT 766.110 6.990 766.510 7.390 ;
        RECT 766.910 6.990 767.310 7.390 ;
        RECT 767.710 6.990 768.110 7.390 ;
        RECT 768.510 6.990 768.910 7.390 ;
        RECT 769.310 6.990 769.710 7.390 ;
        RECT 770.110 6.990 770.510 7.390 ;
      LAYER met2 ;
        RECT 740.320 249.510 765.820 251.310 ;
        RECT 369.540 215.330 378.730 221.480 ;
        RECT 389.540 215.330 398.730 221.480 ;
        RECT 409.540 215.330 418.730 221.480 ;
        RECT 429.540 215.330 438.730 221.480 ;
        RECT 449.540 215.330 458.730 221.480 ;
        RECT 469.540 215.330 478.730 221.480 ;
        RECT 489.540 215.330 498.730 221.480 ;
        RECT 509.540 215.330 518.730 221.480 ;
        RECT 529.540 215.330 538.730 221.480 ;
        RECT 549.540 215.330 558.730 221.480 ;
        RECT 569.540 215.330 578.730 221.480 ;
        RECT 589.540 215.330 598.730 221.480 ;
        RECT 609.540 215.330 618.730 221.480 ;
        RECT 629.540 215.330 638.730 221.480 ;
        RECT 649.540 215.330 658.730 221.480 ;
        RECT 360.860 204.510 370.050 210.660 ;
        RECT 649.750 199.320 658.940 205.510 ;
        RECT 360.860 184.510 370.050 190.660 ;
        RECT 360.860 164.510 370.050 170.660 ;
        RECT 168.470 154.870 171.490 155.280 ;
        RECT 170.590 144.850 170.960 154.870 ;
        RECT 170.550 143.500 171.030 144.850 ;
        RECT 360.860 144.510 370.050 150.660 ;
        RECT 170.550 143.460 175.600 143.500 ;
        RECT 176.180 143.460 231.520 143.480 ;
        RECT 170.550 143.100 231.520 143.460 ;
        RECT 170.550 143.090 223.900 143.100 ;
        RECT 170.550 143.020 175.600 143.090 ;
        RECT 117.550 128.690 118.530 129.590 ;
        RECT 139.450 128.250 140.430 129.150 ;
        RECT 160.240 128.020 161.220 128.920 ;
        RECT 231.120 116.200 231.520 143.100 ;
        RECT 348.190 125.460 349.790 126.360 ;
        RECT 337.240 124.710 337.890 124.840 ;
        RECT 348.200 124.710 349.220 125.460 ;
        RECT 337.240 123.890 349.220 124.710 ;
        RECT 360.860 124.510 370.050 130.660 ;
        RECT 337.240 123.850 349.210 123.890 ;
        RECT 337.240 123.740 337.890 123.850 ;
        RECT 253.940 116.200 254.220 116.220 ;
        RECT 231.070 116.170 255.290 116.200 ;
        RECT 231.070 116.140 281.590 116.170 ;
        RECT 296.400 116.140 302.960 118.430 ;
        RECT 231.070 115.710 302.960 116.140 ;
        RECT 231.070 115.510 255.290 115.710 ;
        RECT 279.870 115.550 302.960 115.710 ;
        RECT 253.940 97.430 254.220 115.510 ;
        RECT 260.200 105.810 262.450 107.890 ;
        RECT 255.670 97.430 257.900 98.370 ;
        RECT 253.940 97.130 257.900 97.430 ;
        RECT 255.670 96.280 257.900 97.130 ;
        RECT 279.870 95.820 280.170 115.550 ;
        RECT 296.400 113.890 302.960 115.550 ;
        RECT 360.860 104.510 370.050 110.660 ;
        RECT 281.630 95.820 283.910 96.770 ;
        RECT 279.870 95.430 283.910 95.820 ;
        RECT 281.630 94.680 283.910 95.430 ;
        RECT 360.860 84.510 370.050 90.660 ;
        RECT 383.330 89.040 391.170 187.730 ;
        RECT 649.750 179.320 658.940 185.510 ;
        RECT 649.750 159.320 658.940 165.510 ;
        RECT 649.750 139.320 658.940 145.510 ;
        RECT 649.750 119.320 658.940 125.510 ;
        RECT 649.750 99.320 658.940 105.510 ;
        RECT 383.330 87.790 391.180 89.040 ;
        RECT 95.520 77.960 98.740 81.430 ;
        RECT 116.100 81.420 116.820 82.040 ;
        RECT 129.430 81.420 130.150 82.040 ;
        RECT 142.735 81.415 143.465 82.040 ;
        RECT 160.650 76.235 169.685 81.980 ;
        RECT 42.870 70.950 44.430 70.970 ;
        RECT 42.870 70.650 44.440 70.950 ;
        RECT 42.870 67.900 43.130 70.650 ;
        RECT 42.870 67.600 44.460 67.900 ;
        RECT 42.870 65.010 43.130 67.600 ;
        RECT 43.720 67.590 44.460 67.600 ;
        RECT 42.870 64.710 44.450 65.010 ;
        RECT 42.870 62.150 43.130 64.710 ;
        RECT 43.670 64.700 44.450 64.710 ;
        RECT 69.660 63.460 70.640 64.360 ;
        RECT 42.870 61.850 44.480 62.150 ;
        RECT 224.020 62.040 230.580 66.580 ;
        RECT 42.870 59.240 43.130 61.850 ;
        RECT 43.730 61.840 44.480 61.850 ;
        RECT 43.740 61.830 44.480 61.840 ;
        RECT 261.130 61.120 267.690 65.660 ;
        RECT 294.290 62.710 300.850 67.250 ;
        RECT 360.290 63.380 371.000 71.710 ;
        RECT 43.690 59.240 44.480 59.250 ;
        RECT 42.870 58.940 44.480 59.240 ;
        RECT 42.870 56.360 43.130 58.940 ;
        RECT 42.870 56.060 44.490 56.360 ;
        RECT 16.750 53.750 18.820 55.840 ;
        RECT 42.870 53.450 43.130 56.060 ;
        RECT 43.740 56.050 44.480 56.060 ;
        RECT 42.870 53.150 44.510 53.450 ;
        RECT 42.870 50.560 43.130 53.150 ;
        RECT 43.760 53.140 44.500 53.150 ;
        RECT 116.060 52.820 116.830 53.455 ;
        RECT 129.480 52.850 130.105 53.460 ;
        RECT 142.800 52.850 143.425 53.480 ;
        RECT 383.330 52.650 391.170 87.790 ;
        RECT 423.690 73.670 431.780 80.110 ;
        RECT 649.750 79.320 658.940 85.510 ;
        RECT 424.320 57.910 424.700 73.670 ;
        RECT 649.750 59.320 658.940 65.510 ;
        RECT 43.720 50.560 44.480 50.570 ;
        RECT 42.870 50.260 44.480 50.560 ;
        RECT 42.870 48.850 43.130 50.260 ;
        RECT 42.860 48.840 43.130 48.850 ;
        RECT 42.860 47.720 43.120 48.840 ;
        RECT 42.860 47.660 44.460 47.720 ;
        RECT 42.860 47.420 44.470 47.660 ;
        RECT 42.860 46.180 43.120 47.420 ;
        RECT 43.720 47.410 44.460 47.420 ;
        RECT 185.850 47.310 186.830 48.210 ;
        RECT 42.850 45.820 43.700 46.180 ;
        RECT 43.230 43.510 43.700 45.820 ;
        RECT 360.860 44.510 370.050 50.660 ;
        RECT 41.760 40.450 44.750 43.510 ;
        RECT 70.050 37.710 71.030 38.610 ;
        RECT 218.960 36.380 221.650 38.730 ;
        RECT 360.860 24.510 370.050 30.660 ;
        RECT 116.060 23.370 116.830 24.005 ;
        RECT 129.430 23.365 130.165 23.980 ;
        RECT 142.770 23.355 143.505 23.970 ;
        RECT 249.210 22.740 249.530 22.770 ;
        RECT 242.710 19.630 244.780 21.720 ;
        RECT 249.210 21.480 249.570 22.740 ;
        RECT 258.090 21.770 258.380 23.060 ;
        RECT 293.710 22.820 294.020 22.830 ;
        RECT 283.970 21.200 284.320 22.230 ;
        RECT 287.910 20.070 288.280 20.710 ;
        RECT 289.200 20.070 289.540 22.550 ;
        RECT 293.710 21.800 294.030 22.820 ;
        RECT 293.710 21.780 294.020 21.800 ;
        RECT 287.910 19.650 289.540 20.070 ;
        RECT 287.910 19.640 288.280 19.650 ;
        RECT 289.200 19.560 289.540 19.650 ;
        RECT 258.160 12.650 258.470 14.160 ;
        RECT 374.170 12.260 383.360 15.150 ;
        RECT 384.070 12.260 384.930 52.650 ;
        RECT 424.320 48.370 424.680 57.910 ;
        RECT 424.320 48.040 424.690 48.370 ;
        RECT 424.330 43.170 424.690 48.040 ;
        RECT 424.330 42.880 424.700 43.170 ;
        RECT 424.340 38.120 424.700 42.880 ;
        RECT 649.750 39.320 658.940 45.510 ;
        RECT 424.340 37.680 424.720 38.120 ;
        RECT 424.360 22.410 424.720 37.680 ;
        RECT 424.350 22.130 424.720 22.410 ;
        RECT 424.350 17.280 424.710 22.130 ;
        RECT 649.750 19.320 658.940 25.510 ;
        RECT 424.350 16.920 424.730 17.280 ;
        RECT 374.170 11.910 384.930 12.260 ;
        RECT 374.170 8.920 383.360 11.910 ;
        RECT 384.070 11.770 384.930 11.910 ;
        RECT 394.170 14.650 395.110 15.130 ;
        RECT 397.810 14.650 403.360 15.130 ;
        RECT 394.170 8.920 403.360 14.650 ;
        RECT 414.170 12.140 423.360 15.130 ;
        RECT 424.370 12.140 424.730 16.920 ;
        RECT 414.170 11.850 424.760 12.140 ;
        RECT 414.170 8.920 423.360 11.850 ;
        RECT 424.370 11.790 424.730 11.850 ;
        RECT 434.170 8.920 443.360 15.130 ;
        RECT 454.170 8.920 463.360 15.130 ;
        RECT 474.170 8.920 483.360 15.130 ;
        RECT 494.170 8.920 503.360 15.130 ;
        RECT 514.170 8.920 523.360 15.130 ;
        RECT 534.170 8.920 543.360 15.130 ;
        RECT 554.170 8.920 563.360 15.130 ;
        RECT 574.170 8.920 583.360 15.130 ;
        RECT 594.170 8.920 603.360 15.130 ;
        RECT 614.170 8.920 623.360 15.130 ;
        RECT 634.170 8.920 643.360 15.130 ;
        RECT 112.040 7.060 113.020 7.960 ;
        RECT 128.950 6.970 129.930 7.870 ;
        RECT 147.420 7.060 148.400 7.960 ;
        RECT 745.610 6.790 771.110 8.590 ;
      LAYER via2 ;
        RECT 740.820 250.510 741.220 250.910 ;
        RECT 741.620 250.510 742.020 250.910 ;
        RECT 742.420 250.510 742.820 250.910 ;
        RECT 743.220 250.510 743.620 250.910 ;
        RECT 744.020 250.510 744.420 250.910 ;
        RECT 744.820 250.510 745.220 250.910 ;
        RECT 745.620 250.510 746.020 250.910 ;
        RECT 746.420 250.510 746.820 250.910 ;
        RECT 747.220 250.510 747.620 250.910 ;
        RECT 748.020 250.510 748.420 250.910 ;
        RECT 748.820 250.510 749.220 250.910 ;
        RECT 749.620 250.510 750.020 250.910 ;
        RECT 750.420 250.510 750.820 250.910 ;
        RECT 751.220 250.510 751.620 250.910 ;
        RECT 752.020 250.510 752.420 250.910 ;
        RECT 752.820 250.510 753.220 250.910 ;
        RECT 753.620 250.510 754.020 250.910 ;
        RECT 754.420 250.510 754.820 250.910 ;
        RECT 755.220 250.510 755.620 250.910 ;
        RECT 756.020 250.510 756.420 250.910 ;
        RECT 756.820 250.510 757.220 250.910 ;
        RECT 757.620 250.510 758.020 250.910 ;
        RECT 758.420 250.510 758.820 250.910 ;
        RECT 759.220 250.510 759.620 250.910 ;
        RECT 760.020 250.510 760.420 250.910 ;
        RECT 760.820 250.510 761.220 250.910 ;
        RECT 761.620 250.510 762.020 250.910 ;
        RECT 762.420 250.510 762.820 250.910 ;
        RECT 763.220 250.510 763.620 250.910 ;
        RECT 764.020 250.510 764.420 250.910 ;
        RECT 764.820 250.510 765.220 250.910 ;
        RECT 740.820 249.710 741.220 250.110 ;
        RECT 741.620 249.710 742.020 250.110 ;
        RECT 742.420 249.710 742.820 250.110 ;
        RECT 743.220 249.710 743.620 250.110 ;
        RECT 744.020 249.710 744.420 250.110 ;
        RECT 744.820 249.710 745.220 250.110 ;
        RECT 745.620 249.710 746.020 250.110 ;
        RECT 746.420 249.710 746.820 250.110 ;
        RECT 747.220 249.710 747.620 250.110 ;
        RECT 748.020 249.710 748.420 250.110 ;
        RECT 748.820 249.710 749.220 250.110 ;
        RECT 749.620 249.710 750.020 250.110 ;
        RECT 750.420 249.710 750.820 250.110 ;
        RECT 751.220 249.710 751.620 250.110 ;
        RECT 752.020 249.710 752.420 250.110 ;
        RECT 752.820 249.710 753.220 250.110 ;
        RECT 753.620 249.710 754.020 250.110 ;
        RECT 754.420 249.710 754.820 250.110 ;
        RECT 755.220 249.710 755.620 250.110 ;
        RECT 756.020 249.710 756.420 250.110 ;
        RECT 756.820 249.710 757.220 250.110 ;
        RECT 757.620 249.710 758.020 250.110 ;
        RECT 758.420 249.710 758.820 250.110 ;
        RECT 759.220 249.710 759.620 250.110 ;
        RECT 760.020 249.710 760.420 250.110 ;
        RECT 760.820 249.710 761.220 250.110 ;
        RECT 761.620 249.710 762.020 250.110 ;
        RECT 762.420 249.710 762.820 250.110 ;
        RECT 763.220 249.710 763.620 250.110 ;
        RECT 764.020 249.710 764.420 250.110 ;
        RECT 764.820 249.710 765.220 250.110 ;
        RECT 370.750 216.540 377.680 220.180 ;
        RECT 390.750 216.540 397.680 220.180 ;
        RECT 410.750 216.540 417.680 220.180 ;
        RECT 430.750 216.540 437.680 220.180 ;
        RECT 450.750 216.540 457.680 220.180 ;
        RECT 470.750 216.540 477.680 220.180 ;
        RECT 490.750 216.540 497.680 220.180 ;
        RECT 510.750 216.540 517.680 220.180 ;
        RECT 530.750 216.540 537.680 220.180 ;
        RECT 550.750 216.540 557.680 220.180 ;
        RECT 570.750 216.540 577.680 220.180 ;
        RECT 590.750 216.540 597.680 220.180 ;
        RECT 610.750 216.540 617.680 220.180 ;
        RECT 630.750 216.540 637.680 220.180 ;
        RECT 650.750 216.540 657.680 220.180 ;
        RECT 362.070 205.720 369.000 209.360 ;
        RECT 650.960 200.530 657.890 204.170 ;
        RECT 362.070 185.720 369.000 189.360 ;
        RECT 362.070 165.720 369.000 169.360 ;
        RECT 168.630 154.940 168.920 155.220 ;
        RECT 170.630 154.940 170.920 155.220 ;
        RECT 362.070 145.720 369.000 149.360 ;
        RECT 117.690 128.810 118.420 129.440 ;
        RECT 139.590 128.370 140.320 129.000 ;
        RECT 160.380 128.140 161.110 128.770 ;
        RECT 362.070 125.720 369.000 129.360 ;
        RECT 260.260 107.480 262.420 107.840 ;
        RECT 260.260 105.880 262.420 106.240 ;
        RECT 297.440 114.990 302.240 117.460 ;
        RECT 362.070 105.720 369.000 109.360 ;
        RECT 362.070 85.720 369.000 89.360 ;
        RECT 650.960 180.530 657.890 184.170 ;
        RECT 650.960 160.530 657.890 164.170 ;
        RECT 650.960 140.530 657.890 144.170 ;
        RECT 650.960 120.530 657.890 124.170 ;
        RECT 650.960 100.530 657.890 104.170 ;
        RECT 116.200 81.470 116.730 82.000 ;
        RECT 129.520 81.470 130.050 82.000 ;
        RECT 142.830 81.470 143.360 82.000 ;
        RECT 95.820 78.480 97.480 80.650 ;
        RECT 161.945 77.485 167.955 80.995 ;
        RECT 69.800 63.580 70.530 64.210 ;
        RECT 225.060 63.140 229.860 65.610 ;
        RECT 262.170 62.220 266.970 64.690 ;
        RECT 295.330 63.810 300.130 66.280 ;
        RECT 362.070 65.720 369.000 69.360 ;
        RECT 17.040 54.000 18.530 55.610 ;
        RECT 116.170 52.875 116.700 53.405 ;
        RECT 129.550 52.910 130.010 53.380 ;
        RECT 142.880 52.910 143.340 53.380 ;
        RECT 650.960 80.530 657.890 84.170 ;
        RECT 424.770 74.750 430.720 78.740 ;
        RECT 650.960 60.530 657.890 64.170 ;
        RECT 185.990 47.430 186.720 48.060 ;
        RECT 362.070 45.720 369.000 49.360 ;
        RECT 42.110 40.810 44.410 43.210 ;
        RECT 70.190 37.830 70.920 38.460 ;
        RECT 219.300 36.600 221.140 38.590 ;
        RECT 362.070 25.720 369.000 29.360 ;
        RECT 116.210 23.430 116.670 23.900 ;
        RECT 129.560 23.430 130.020 23.900 ;
        RECT 142.890 23.430 143.350 23.900 ;
        RECT 249.240 21.540 249.520 22.700 ;
        RECT 258.090 21.830 258.370 22.990 ;
        RECT 242.970 19.940 244.450 21.370 ;
        RECT 284.030 21.280 284.310 22.160 ;
        RECT 287.960 20.250 288.280 20.660 ;
        RECT 293.740 21.860 294.020 22.760 ;
        RECT 258.170 12.720 258.460 14.110 ;
        RECT 375.380 10.130 382.310 13.770 ;
        RECT 650.960 40.530 657.890 44.170 ;
        RECT 650.960 20.530 657.890 24.170 ;
        RECT 395.380 10.130 402.310 13.770 ;
        RECT 415.380 10.130 422.310 13.770 ;
        RECT 435.380 10.130 442.310 13.770 ;
        RECT 455.380 10.130 462.310 13.770 ;
        RECT 475.380 10.130 482.310 13.770 ;
        RECT 495.380 10.130 502.310 13.770 ;
        RECT 515.380 10.130 522.310 13.770 ;
        RECT 535.380 10.130 542.310 13.770 ;
        RECT 555.380 10.130 562.310 13.770 ;
        RECT 575.380 10.130 582.310 13.770 ;
        RECT 595.380 10.130 602.310 13.770 ;
        RECT 615.380 10.130 622.310 13.770 ;
        RECT 635.380 10.130 642.310 13.770 ;
        RECT 112.180 7.180 112.910 7.810 ;
        RECT 129.090 7.090 129.820 7.720 ;
        RECT 147.560 7.180 148.290 7.810 ;
        RECT 746.110 7.790 746.510 8.190 ;
        RECT 746.910 7.790 747.310 8.190 ;
        RECT 747.710 7.790 748.110 8.190 ;
        RECT 748.510 7.790 748.910 8.190 ;
        RECT 749.310 7.790 749.710 8.190 ;
        RECT 750.110 7.790 750.510 8.190 ;
        RECT 750.910 7.790 751.310 8.190 ;
        RECT 751.710 7.790 752.110 8.190 ;
        RECT 752.510 7.790 752.910 8.190 ;
        RECT 753.310 7.790 753.710 8.190 ;
        RECT 754.110 7.790 754.510 8.190 ;
        RECT 754.910 7.790 755.310 8.190 ;
        RECT 755.710 7.790 756.110 8.190 ;
        RECT 756.510 7.790 756.910 8.190 ;
        RECT 757.310 7.790 757.710 8.190 ;
        RECT 758.110 7.790 758.510 8.190 ;
        RECT 758.910 7.790 759.310 8.190 ;
        RECT 759.710 7.790 760.110 8.190 ;
        RECT 760.510 7.790 760.910 8.190 ;
        RECT 761.310 7.790 761.710 8.190 ;
        RECT 762.110 7.790 762.510 8.190 ;
        RECT 762.910 7.790 763.310 8.190 ;
        RECT 763.710 7.790 764.110 8.190 ;
        RECT 764.510 7.790 764.910 8.190 ;
        RECT 765.310 7.790 765.710 8.190 ;
        RECT 766.110 7.790 766.510 8.190 ;
        RECT 766.910 7.790 767.310 8.190 ;
        RECT 767.710 7.790 768.110 8.190 ;
        RECT 768.510 7.790 768.910 8.190 ;
        RECT 769.310 7.790 769.710 8.190 ;
        RECT 770.110 7.790 770.510 8.190 ;
        RECT 746.110 6.990 746.510 7.390 ;
        RECT 746.910 6.990 747.310 7.390 ;
        RECT 747.710 6.990 748.110 7.390 ;
        RECT 748.510 6.990 748.910 7.390 ;
        RECT 749.310 6.990 749.710 7.390 ;
        RECT 750.110 6.990 750.510 7.390 ;
        RECT 750.910 6.990 751.310 7.390 ;
        RECT 751.710 6.990 752.110 7.390 ;
        RECT 752.510 6.990 752.910 7.390 ;
        RECT 753.310 6.990 753.710 7.390 ;
        RECT 754.110 6.990 754.510 7.390 ;
        RECT 754.910 6.990 755.310 7.390 ;
        RECT 755.710 6.990 756.110 7.390 ;
        RECT 756.510 6.990 756.910 7.390 ;
        RECT 757.310 6.990 757.710 7.390 ;
        RECT 758.110 6.990 758.510 7.390 ;
        RECT 758.910 6.990 759.310 7.390 ;
        RECT 759.710 6.990 760.110 7.390 ;
        RECT 760.510 6.990 760.910 7.390 ;
        RECT 761.310 6.990 761.710 7.390 ;
        RECT 762.110 6.990 762.510 7.390 ;
        RECT 762.910 6.990 763.310 7.390 ;
        RECT 763.710 6.990 764.110 7.390 ;
        RECT 764.510 6.990 764.910 7.390 ;
        RECT 765.310 6.990 765.710 7.390 ;
        RECT 766.110 6.990 766.510 7.390 ;
        RECT 766.910 6.990 767.310 7.390 ;
        RECT 767.710 6.990 768.110 7.390 ;
        RECT 768.510 6.990 768.910 7.390 ;
        RECT 769.310 6.990 769.710 7.390 ;
        RECT 770.110 6.990 770.510 7.390 ;
      LAYER met3 ;
        RECT 740.320 249.510 765.820 251.310 ;
        RECT 369.540 215.330 378.730 221.480 ;
        RECT 389.540 215.330 398.730 221.480 ;
        RECT 409.540 215.330 418.730 221.480 ;
        RECT 429.540 215.330 438.730 221.480 ;
        RECT 449.540 215.330 458.730 221.480 ;
        RECT 469.540 215.330 478.730 221.480 ;
        RECT 489.540 215.330 498.730 221.480 ;
        RECT 509.540 215.330 518.730 221.480 ;
        RECT 529.540 215.330 538.730 221.480 ;
        RECT 549.540 215.330 558.730 221.480 ;
        RECT 569.540 215.330 578.730 221.480 ;
        RECT 589.540 215.330 598.730 221.480 ;
        RECT 609.540 215.330 618.730 221.480 ;
        RECT 629.540 215.330 638.730 221.480 ;
        RECT 649.540 215.330 658.730 221.480 ;
        RECT 360.860 204.510 370.050 210.660 ;
        RECT 649.750 199.320 658.940 205.510 ;
        RECT 360.860 184.510 370.050 190.660 ;
        RECT 360.860 164.510 370.050 170.660 ;
        RECT 421.465 165.720 612.570 191.310 ;
        RECT 649.750 179.320 658.940 185.510 ;
        RECT 421.465 165.710 548.400 165.720 ;
        RECT 421.465 165.560 495.430 165.710 ;
        RECT 421.465 164.950 465.840 165.560 ;
        RECT 470.290 164.950 495.430 165.560 ;
        RECT 499.940 164.950 548.400 165.710 ;
        RECT 556.570 165.460 612.570 165.720 ;
        RECT 556.570 164.950 576.410 165.460 ;
        RECT 580.970 164.950 612.570 165.460 ;
        RECT 168.470 154.870 171.490 155.280 ;
        RECT 360.860 144.510 370.050 150.660 ;
        RECT 117.550 128.690 118.530 129.590 ;
        RECT 139.450 128.250 140.430 129.150 ;
        RECT 160.240 128.020 161.220 128.920 ;
        RECT 360.860 124.510 370.050 130.660 ;
        RECT 150.230 119.350 155.540 122.500 ;
        RECT 151.020 83.080 154.350 119.350 ;
        RECT 258.980 116.060 259.410 116.290 ;
        RECT 296.400 116.060 302.960 118.430 ;
        RECT 258.980 115.640 302.960 116.060 ;
        RECT 258.980 107.020 259.410 115.640 ;
        RECT 296.400 113.890 302.960 115.640 ;
        RECT 260.190 107.020 262.460 107.910 ;
        RECT 258.980 106.660 262.460 107.020 ;
        RECT 260.190 105.800 262.460 106.660 ;
        RECT 360.860 104.510 370.050 110.660 ;
        RECT 421.630 107.780 447.165 164.950 ;
        RECT 586.375 163.370 611.910 164.950 ;
        RECT 586.375 137.780 612.070 163.370 ;
        RECT 649.750 159.320 658.940 165.510 ;
        RECT 649.750 139.320 658.940 145.510 ;
        RECT 586.375 135.590 611.910 137.780 ;
        RECT 586.375 110.060 612.070 135.590 ;
        RECT 649.750 119.320 658.940 125.510 ;
        RECT 449.150 107.780 474.380 107.870 ;
        RECT 476.770 107.780 502.000 107.870 ;
        RECT 504.295 107.780 529.525 107.870 ;
        RECT 531.715 107.780 547.500 108.070 ;
        RECT 421.135 107.620 547.500 107.780 ;
        RECT 552.120 107.780 556.945 108.070 ;
        RECT 586.375 107.870 611.910 110.060 ;
        RECT 559.340 107.780 584.570 107.870 ;
        RECT 586.375 107.780 612.070 107.870 ;
        RECT 552.120 107.620 612.070 107.780 ;
        RECT 360.860 84.510 370.050 90.660 ;
        RECT 95.520 77.960 98.740 81.430 ;
        RECT 116.100 81.420 116.820 82.040 ;
        RECT 129.430 81.420 130.150 82.040 ;
        RECT 142.735 81.415 143.465 82.040 ;
        RECT 150.640 78.180 154.720 83.080 ;
        RECT 421.135 82.310 612.070 107.620 ;
        RECT 649.750 99.320 658.940 105.510 ;
        RECT 160.795 76.570 169.515 81.785 ;
        RECT 421.135 81.585 611.910 82.310 ;
        RECT 423.630 73.680 431.910 81.585 ;
        RECT 649.750 79.320 658.940 85.510 ;
        RECT 423.690 73.670 431.780 73.680 ;
        RECT 69.660 63.460 70.640 64.360 ;
        RECT 224.020 62.040 230.580 66.580 ;
        RECT 261.130 61.120 267.690 65.660 ;
        RECT 294.290 62.710 300.850 67.250 ;
        RECT 360.290 63.380 371.000 71.710 ;
        RECT 649.750 59.320 658.940 65.510 ;
        RECT 16.750 53.750 18.820 55.840 ;
        RECT 116.060 52.820 116.830 53.455 ;
        RECT 129.480 52.850 130.105 53.460 ;
        RECT 142.800 52.850 143.425 53.480 ;
        RECT 185.850 47.310 186.830 48.210 ;
        RECT 360.860 44.510 370.050 50.660 ;
        RECT 41.760 40.450 44.750 43.510 ;
        RECT 649.750 39.320 658.940 45.510 ;
        RECT 70.050 37.710 71.030 38.610 ;
        RECT 218.960 36.380 221.650 38.730 ;
        RECT 360.860 24.510 370.050 30.660 ;
        RECT 116.060 23.370 116.830 24.005 ;
        RECT 129.430 23.365 130.165 23.980 ;
        RECT 142.770 23.355 143.505 23.970 ;
        RECT 249.210 21.910 249.570 22.770 ;
        RECT 242.710 21.070 244.780 21.720 ;
        RECT 248.680 21.480 249.570 21.910 ;
        RECT 258.040 22.370 258.430 23.060 ;
        RECT 258.040 21.760 258.490 22.370 ;
        RECT 248.680 21.470 249.560 21.480 ;
        RECT 248.710 21.070 249.100 21.470 ;
        RECT 242.710 20.260 249.100 21.070 ;
        RECT 242.710 19.630 244.780 20.260 ;
        RECT 248.710 13.180 249.100 20.260 ;
        RECT 258.130 15.330 258.490 21.760 ;
        RECT 283.940 22.230 284.340 22.240 ;
        RECT 283.940 22.180 284.360 22.230 ;
        RECT 293.710 22.180 294.050 22.840 ;
        RECT 283.940 21.750 294.050 22.180 ;
        RECT 283.940 21.220 284.360 21.750 ;
        RECT 293.750 21.740 294.050 21.750 ;
        RECT 283.960 21.210 284.360 21.220 ;
        RECT 283.970 20.700 284.270 21.210 ;
        RECT 287.910 20.700 288.320 20.710 ;
        RECT 283.950 20.200 288.320 20.700 ;
        RECT 258.130 14.050 258.510 15.330 ;
        RECT 248.710 13.170 256.120 13.180 ;
        RECT 258.130 13.170 258.490 14.050 ;
        RECT 248.710 12.720 258.490 13.170 ;
        RECT 248.710 12.660 249.100 12.720 ;
        RECT 251.600 12.710 258.490 12.720 ;
        RECT 258.130 12.660 258.490 12.710 ;
        RECT 258.140 12.540 258.490 12.660 ;
        RECT 258.140 12.520 260.740 12.540 ;
        RECT 283.970 12.520 284.270 20.200 ;
        RECT 287.910 20.190 288.320 20.200 ;
        RECT 649.750 19.320 658.940 25.510 ;
        RECT 258.140 12.220 284.300 12.520 ;
        RECT 260.550 12.210 284.300 12.220 ;
        RECT 374.170 8.920 383.360 15.150 ;
        RECT 394.170 14.650 395.110 15.130 ;
        RECT 397.810 14.650 403.360 15.130 ;
        RECT 394.170 8.920 403.360 14.650 ;
        RECT 414.170 8.920 423.360 15.130 ;
        RECT 434.170 8.920 443.360 15.130 ;
        RECT 454.170 8.920 463.360 15.130 ;
        RECT 474.170 8.920 483.360 15.130 ;
        RECT 494.170 8.920 503.360 15.130 ;
        RECT 514.170 8.920 523.360 15.130 ;
        RECT 534.170 8.920 543.360 15.130 ;
        RECT 554.170 8.920 563.360 15.130 ;
        RECT 574.170 8.920 583.360 15.130 ;
        RECT 594.170 8.920 603.360 15.130 ;
        RECT 614.170 8.920 623.360 15.130 ;
        RECT 634.170 8.920 643.360 15.130 ;
        RECT 112.040 7.060 113.020 7.960 ;
        RECT 128.950 6.970 129.930 7.870 ;
        RECT 147.420 7.060 148.400 7.960 ;
        RECT 745.610 6.790 771.110 8.590 ;
      LAYER via3 ;
        RECT 740.820 250.510 741.220 250.910 ;
        RECT 741.620 250.510 742.020 250.910 ;
        RECT 742.420 250.510 742.820 250.910 ;
        RECT 743.220 250.510 743.620 250.910 ;
        RECT 744.020 250.510 744.420 250.910 ;
        RECT 744.820 250.510 745.220 250.910 ;
        RECT 745.620 250.510 746.020 250.910 ;
        RECT 746.420 250.510 746.820 250.910 ;
        RECT 747.220 250.510 747.620 250.910 ;
        RECT 748.020 250.510 748.420 250.910 ;
        RECT 748.820 250.510 749.220 250.910 ;
        RECT 749.620 250.510 750.020 250.910 ;
        RECT 750.420 250.510 750.820 250.910 ;
        RECT 751.220 250.510 751.620 250.910 ;
        RECT 752.020 250.510 752.420 250.910 ;
        RECT 752.820 250.510 753.220 250.910 ;
        RECT 753.620 250.510 754.020 250.910 ;
        RECT 754.420 250.510 754.820 250.910 ;
        RECT 755.220 250.510 755.620 250.910 ;
        RECT 756.020 250.510 756.420 250.910 ;
        RECT 756.820 250.510 757.220 250.910 ;
        RECT 757.620 250.510 758.020 250.910 ;
        RECT 758.420 250.510 758.820 250.910 ;
        RECT 759.220 250.510 759.620 250.910 ;
        RECT 760.020 250.510 760.420 250.910 ;
        RECT 760.820 250.510 761.220 250.910 ;
        RECT 761.620 250.510 762.020 250.910 ;
        RECT 762.420 250.510 762.820 250.910 ;
        RECT 763.220 250.510 763.620 250.910 ;
        RECT 764.020 250.510 764.420 250.910 ;
        RECT 764.820 250.510 765.220 250.910 ;
        RECT 740.820 249.710 741.220 250.110 ;
        RECT 741.620 249.710 742.020 250.110 ;
        RECT 742.420 249.710 742.820 250.110 ;
        RECT 743.220 249.710 743.620 250.110 ;
        RECT 744.020 249.710 744.420 250.110 ;
        RECT 744.820 249.710 745.220 250.110 ;
        RECT 745.620 249.710 746.020 250.110 ;
        RECT 746.420 249.710 746.820 250.110 ;
        RECT 747.220 249.710 747.620 250.110 ;
        RECT 748.020 249.710 748.420 250.110 ;
        RECT 748.820 249.710 749.220 250.110 ;
        RECT 749.620 249.710 750.020 250.110 ;
        RECT 750.420 249.710 750.820 250.110 ;
        RECT 751.220 249.710 751.620 250.110 ;
        RECT 752.020 249.710 752.420 250.110 ;
        RECT 752.820 249.710 753.220 250.110 ;
        RECT 753.620 249.710 754.020 250.110 ;
        RECT 754.420 249.710 754.820 250.110 ;
        RECT 755.220 249.710 755.620 250.110 ;
        RECT 756.020 249.710 756.420 250.110 ;
        RECT 756.820 249.710 757.220 250.110 ;
        RECT 757.620 249.710 758.020 250.110 ;
        RECT 758.420 249.710 758.820 250.110 ;
        RECT 759.220 249.710 759.620 250.110 ;
        RECT 760.020 249.710 760.420 250.110 ;
        RECT 760.820 249.710 761.220 250.110 ;
        RECT 761.620 249.710 762.020 250.110 ;
        RECT 762.420 249.710 762.820 250.110 ;
        RECT 763.220 249.710 763.620 250.110 ;
        RECT 764.020 249.710 764.420 250.110 ;
        RECT 764.820 249.710 765.220 250.110 ;
        RECT 370.750 216.540 377.680 220.180 ;
        RECT 390.750 216.540 397.680 220.180 ;
        RECT 410.750 216.540 417.680 220.180 ;
        RECT 430.750 216.540 437.680 220.180 ;
        RECT 450.750 216.540 457.680 220.180 ;
        RECT 470.750 216.540 477.680 220.180 ;
        RECT 490.750 216.540 497.680 220.180 ;
        RECT 510.750 216.540 517.680 220.180 ;
        RECT 530.750 216.540 537.680 220.180 ;
        RECT 550.750 216.540 557.680 220.180 ;
        RECT 570.750 216.540 577.680 220.180 ;
        RECT 590.750 216.540 597.680 220.180 ;
        RECT 610.750 216.540 617.680 220.180 ;
        RECT 630.750 216.540 637.680 220.180 ;
        RECT 650.750 216.540 657.680 220.180 ;
        RECT 362.070 205.720 369.000 209.360 ;
        RECT 650.960 200.530 657.890 204.170 ;
        RECT 362.070 185.720 369.000 189.360 ;
        RECT 362.070 165.720 369.000 169.360 ;
        RECT 650.960 180.530 657.890 184.170 ;
        RECT 168.630 154.940 168.950 155.260 ;
        RECT 170.630 154.940 170.950 155.260 ;
        RECT 362.070 145.720 369.000 149.360 ;
        RECT 117.690 128.810 118.420 129.440 ;
        RECT 139.590 128.370 140.320 129.000 ;
        RECT 160.380 128.140 161.110 128.770 ;
        RECT 361.850 125.520 369.110 129.450 ;
        RECT 151.650 120.060 153.190 121.220 ;
        RECT 297.440 114.990 302.240 117.460 ;
        RECT 362.070 105.720 369.000 109.360 ;
        RECT 650.960 160.530 657.890 164.170 ;
        RECT 650.960 140.530 657.890 144.170 ;
        RECT 650.960 120.530 657.890 124.170 ;
        RECT 362.070 85.720 369.000 89.360 ;
        RECT 116.200 81.470 116.730 82.000 ;
        RECT 129.520 81.470 130.050 82.000 ;
        RECT 142.830 81.470 143.360 82.000 ;
        RECT 95.820 78.480 97.480 80.650 ;
        RECT 650.960 100.530 657.890 104.170 ;
        RECT 152.030 79.080 154.160 80.580 ;
        RECT 161.345 77.315 168.340 81.280 ;
        RECT 650.960 80.530 657.890 84.170 ;
        RECT 424.770 74.750 430.720 78.740 ;
        RECT 69.800 63.580 70.530 64.210 ;
        RECT 225.060 63.140 229.860 65.610 ;
        RECT 262.170 62.220 266.970 64.690 ;
        RECT 295.330 63.810 300.130 66.280 ;
        RECT 360.700 63.900 370.600 71.350 ;
        RECT 650.960 60.530 657.890 64.170 ;
        RECT 17.040 54.000 18.530 55.610 ;
        RECT 116.170 52.875 116.700 53.405 ;
        RECT 129.550 52.910 130.010 53.380 ;
        RECT 142.880 52.910 143.340 53.380 ;
        RECT 185.990 47.430 186.720 48.060 ;
        RECT 362.070 45.720 369.000 49.360 ;
        RECT 42.110 40.810 44.410 43.210 ;
        RECT 650.960 40.530 657.890 44.170 ;
        RECT 70.190 37.830 70.920 38.460 ;
        RECT 219.300 36.600 221.140 38.590 ;
        RECT 362.070 25.720 369.000 29.360 ;
        RECT 116.210 23.430 116.670 23.900 ;
        RECT 129.560 23.430 130.020 23.900 ;
        RECT 142.890 23.430 143.350 23.900 ;
        RECT 249.220 21.540 249.540 22.710 ;
        RECT 242.970 19.940 244.450 21.370 ;
        RECT 650.960 20.530 657.890 24.170 ;
        RECT 375.380 10.130 382.310 13.770 ;
        RECT 395.380 10.130 402.310 13.770 ;
        RECT 415.380 10.130 422.310 13.770 ;
        RECT 435.380 10.130 442.310 13.770 ;
        RECT 455.380 10.130 462.310 13.770 ;
        RECT 475.380 10.130 482.310 13.770 ;
        RECT 495.380 10.130 502.310 13.770 ;
        RECT 515.380 10.130 522.310 13.770 ;
        RECT 535.380 10.130 542.310 13.770 ;
        RECT 555.380 10.130 562.310 13.770 ;
        RECT 575.380 10.130 582.310 13.770 ;
        RECT 595.380 10.130 602.310 13.770 ;
        RECT 615.380 10.130 622.310 13.770 ;
        RECT 635.380 10.130 642.310 13.770 ;
        RECT 112.180 7.180 112.910 7.810 ;
        RECT 129.090 7.090 129.820 7.720 ;
        RECT 147.560 7.180 148.290 7.810 ;
        RECT 746.110 7.790 746.510 8.190 ;
        RECT 746.910 7.790 747.310 8.190 ;
        RECT 747.710 7.790 748.110 8.190 ;
        RECT 748.510 7.790 748.910 8.190 ;
        RECT 749.310 7.790 749.710 8.190 ;
        RECT 750.110 7.790 750.510 8.190 ;
        RECT 750.910 7.790 751.310 8.190 ;
        RECT 751.710 7.790 752.110 8.190 ;
        RECT 752.510 7.790 752.910 8.190 ;
        RECT 753.310 7.790 753.710 8.190 ;
        RECT 754.110 7.790 754.510 8.190 ;
        RECT 754.910 7.790 755.310 8.190 ;
        RECT 755.710 7.790 756.110 8.190 ;
        RECT 756.510 7.790 756.910 8.190 ;
        RECT 757.310 7.790 757.710 8.190 ;
        RECT 758.110 7.790 758.510 8.190 ;
        RECT 758.910 7.790 759.310 8.190 ;
        RECT 759.710 7.790 760.110 8.190 ;
        RECT 760.510 7.790 760.910 8.190 ;
        RECT 761.310 7.790 761.710 8.190 ;
        RECT 762.110 7.790 762.510 8.190 ;
        RECT 762.910 7.790 763.310 8.190 ;
        RECT 763.710 7.790 764.110 8.190 ;
        RECT 764.510 7.790 764.910 8.190 ;
        RECT 765.310 7.790 765.710 8.190 ;
        RECT 766.110 7.790 766.510 8.190 ;
        RECT 766.910 7.790 767.310 8.190 ;
        RECT 767.710 7.790 768.110 8.190 ;
        RECT 768.510 7.790 768.910 8.190 ;
        RECT 769.310 7.790 769.710 8.190 ;
        RECT 770.110 7.790 770.510 8.190 ;
        RECT 746.110 6.990 746.510 7.390 ;
        RECT 746.910 6.990 747.310 7.390 ;
        RECT 747.710 6.990 748.110 7.390 ;
        RECT 748.510 6.990 748.910 7.390 ;
        RECT 749.310 6.990 749.710 7.390 ;
        RECT 750.110 6.990 750.510 7.390 ;
        RECT 750.910 6.990 751.310 7.390 ;
        RECT 751.710 6.990 752.110 7.390 ;
        RECT 752.510 6.990 752.910 7.390 ;
        RECT 753.310 6.990 753.710 7.390 ;
        RECT 754.110 6.990 754.510 7.390 ;
        RECT 754.910 6.990 755.310 7.390 ;
        RECT 755.710 6.990 756.110 7.390 ;
        RECT 756.510 6.990 756.910 7.390 ;
        RECT 757.310 6.990 757.710 7.390 ;
        RECT 758.110 6.990 758.510 7.390 ;
        RECT 758.910 6.990 759.310 7.390 ;
        RECT 759.710 6.990 760.110 7.390 ;
        RECT 760.510 6.990 760.910 7.390 ;
        RECT 761.310 6.990 761.710 7.390 ;
        RECT 762.110 6.990 762.510 7.390 ;
        RECT 762.910 6.990 763.310 7.390 ;
        RECT 763.710 6.990 764.110 7.390 ;
        RECT 764.510 6.990 764.910 7.390 ;
        RECT 765.310 6.990 765.710 7.390 ;
        RECT 766.110 6.990 766.510 7.390 ;
        RECT 766.910 6.990 767.310 7.390 ;
        RECT 767.710 6.990 768.110 7.390 ;
        RECT 768.510 6.990 768.910 7.390 ;
        RECT 769.310 6.990 769.710 7.390 ;
        RECT 770.110 6.990 770.510 7.390 ;
      LAYER met4 ;
        RECT -7.880 -28.090 8.410 357.670 ;
        RECT 369.540 215.330 378.730 221.480 ;
        RECT 389.540 215.330 398.730 221.480 ;
        RECT 409.540 215.330 418.730 221.480 ;
        RECT 429.540 215.330 438.730 221.480 ;
        RECT 449.540 215.330 458.730 221.480 ;
        RECT 469.540 215.330 478.730 221.480 ;
        RECT 489.540 215.330 498.730 221.480 ;
        RECT 509.540 215.330 518.730 221.480 ;
        RECT 529.540 215.330 538.730 221.480 ;
        RECT 549.540 215.330 558.730 221.480 ;
        RECT 569.540 215.330 578.730 221.480 ;
        RECT 589.540 215.330 598.730 221.480 ;
        RECT 609.540 215.330 618.730 221.480 ;
        RECT 629.540 215.330 638.730 221.480 ;
        RECT 649.540 215.330 658.730 221.480 ;
        RECT 360.860 204.510 370.050 210.660 ;
        RECT 649.750 199.320 658.940 205.510 ;
        RECT 360.860 184.510 370.050 190.660 ;
        RECT 423.960 183.260 432.240 183.425 ;
        RECT 423.960 183.095 597.655 183.260 ;
        RECT 423.960 172.000 597.985 183.095 ;
        RECT 649.750 179.320 658.940 185.510 ;
        RECT 360.860 164.510 370.050 170.660 ;
        RECT 168.470 154.870 171.490 155.280 ;
        RECT 360.860 144.510 370.050 150.660 ;
        RECT 117.450 130.600 118.600 139.740 ;
        RECT 139.350 130.600 140.500 139.300 ;
        RECT 117.180 129.890 140.570 130.600 ;
        RECT 151.200 129.890 153.950 130.030 ;
        RECT 160.140 129.890 161.290 139.070 ;
        RECT 360.860 130.630 370.050 130.660 ;
        RECT 117.180 127.860 161.490 129.890 ;
        RECT 151.200 122.500 153.950 127.860 ;
        RECT 150.230 119.350 155.540 122.500 ;
        RECT 296.400 116.260 302.960 118.430 ;
        RECT 296.370 114.790 302.960 116.260 ;
        RECT 296.400 113.890 302.960 114.790 ;
        RECT 87.290 84.155 103.830 84.210 ;
        RECT 106.530 84.155 109.040 84.180 ;
        RECT 111.120 84.155 113.000 84.330 ;
        RECT 87.290 84.150 113.770 84.155 ;
        RECT 115.510 84.150 118.610 84.180 ;
        RECT 87.290 83.650 118.610 84.150 ;
        RECT 87.290 82.105 118.660 83.650 ;
        RECT 150.640 82.125 154.720 83.080 ;
        RECT 167.240 82.125 179.080 82.230 ;
        RECT 87.290 82.080 137.810 82.105 ;
        RECT 142.760 82.080 147.920 82.125 ;
        RECT 87.290 82.070 147.920 82.080 ;
        RECT 149.850 82.070 179.080 82.125 ;
        RECT 87.290 81.170 179.080 82.070 ;
        RECT 87.290 81.140 118.610 81.170 ;
        RECT 87.290 78.430 116.970 81.140 ;
        RECT 129.430 80.045 130.150 81.170 ;
        RECT 87.290 78.405 116.995 78.430 ;
        RECT 87.290 77.850 103.830 78.405 ;
        RECT 87.290 77.840 96.300 77.850 ;
        RECT 69.560 66.890 70.710 74.510 ;
        RECT 106.290 71.120 109.740 78.405 ;
        RECT 115.870 78.240 116.995 78.405 ;
        RECT 129.405 78.270 130.175 80.045 ;
        RECT 142.025 79.370 179.080 81.170 ;
        RECT 142.020 78.310 179.080 79.370 ;
        RECT 115.870 78.010 117.010 78.240 ;
        RECT 129.330 78.080 130.340 78.270 ;
        RECT 115.870 74.410 117.190 78.010 ;
        RECT 129.180 74.480 130.500 78.080 ;
        RECT 141.990 77.760 179.080 78.310 ;
        RECT 141.990 77.380 147.730 77.760 ;
        RECT 141.990 77.370 147.280 77.380 ;
        RECT 141.990 75.510 146.380 77.370 ;
        RECT 156.060 76.070 179.080 77.760 ;
        RECT 156.060 75.970 170.310 76.070 ;
        RECT 116.000 74.250 117.010 74.410 ;
        RECT 129.330 74.280 130.340 74.480 ;
        RECT 141.990 74.410 146.280 75.510 ;
        RECT 116.060 72.605 116.995 74.250 ;
        RECT 129.405 72.705 130.175 74.280 ;
        RECT 142.035 72.725 146.280 74.410 ;
        RECT 69.070 65.880 71.330 66.890 ;
        RECT 106.530 65.880 109.040 71.120 ;
        RECT 69.070 62.500 109.080 65.880 ;
        RECT 16.750 53.750 18.820 55.840 ;
        RECT 17.090 41.830 18.630 53.750 ;
        RECT 69.070 43.830 71.330 62.500 ;
        RECT 106.530 62.380 109.040 62.500 ;
        RECT 116.060 56.450 116.830 72.605 ;
        RECT 115.820 53.545 117.060 56.450 ;
        RECT 129.430 56.180 130.150 72.705 ;
        RECT 142.775 60.955 143.495 72.725 ;
        RECT 175.870 62.440 178.910 76.070 ;
        RECT 299.050 67.320 300.790 113.890 ;
        RECT 360.560 71.710 370.220 130.630 ;
        RECT 423.960 100.635 432.240 172.000 ;
        RECT 588.880 100.635 597.985 172.000 ;
        RECT 649.750 159.320 658.940 165.510 ;
        RECT 649.750 139.320 658.940 145.510 ;
        RECT 649.750 119.320 658.940 125.510 ;
        RECT 423.630 88.880 598.810 100.635 ;
        RECT 649.750 99.320 658.940 105.510 ;
        RECT 423.630 73.680 431.910 88.880 ;
        RECT 588.880 88.380 597.985 88.880 ;
        RECT 649.750 79.320 658.940 85.510 ;
        RECT 360.290 71.660 371.000 71.710 ;
        RECT 360.290 67.360 371.180 71.660 ;
        RECT 352.930 67.320 371.180 67.360 ;
        RECT 294.910 67.250 371.180 67.320 ;
        RECT 224.020 65.080 230.580 66.580 ;
        RECT 261.130 65.080 267.690 65.660 ;
        RECT 294.290 65.080 371.180 67.250 ;
        RECT 224.020 63.610 371.180 65.080 ;
        RECT 142.775 59.715 143.500 60.955 ;
        RECT 142.775 56.220 143.495 59.715 ;
        RECT 129.240 53.545 130.480 56.180 ;
        RECT 142.570 53.545 143.810 56.220 ;
        RECT 115.730 52.890 143.810 53.545 ;
        RECT 115.730 52.610 143.570 52.890 ;
        RECT 115.930 50.750 116.910 52.610 ;
        RECT 115.930 48.470 116.940 50.750 ;
        RECT 116.010 45.370 116.940 48.470 ;
        RECT 129.240 48.380 130.220 52.610 ;
        RECT 129.240 48.330 130.230 48.380 ;
        RECT 115.950 45.040 117.040 45.370 ;
        RECT 129.240 45.100 130.330 48.330 ;
        RECT 142.590 48.200 143.570 52.610 ;
        RECT 175.830 48.810 178.960 62.440 ;
        RECT 224.020 62.040 230.580 63.610 ;
        RECT 185.750 48.810 186.900 55.110 ;
        RECT 175.830 48.450 187.180 48.810 ;
        RECT 212.910 48.450 214.640 48.780 ;
        RECT 226.150 48.450 227.670 62.040 ;
        RECT 261.130 61.120 267.690 63.610 ;
        RECT 294.290 63.420 371.180 63.610 ;
        RECT 294.290 62.710 300.850 63.420 ;
        RECT 142.510 45.910 143.580 48.200 ;
        RECT 175.830 47.190 227.670 48.450 ;
        RECT 175.830 47.030 187.180 47.190 ;
        RECT 142.510 45.870 147.770 45.910 ;
        RECT 142.510 45.205 148.840 45.870 ;
        RECT 115.990 44.940 116.950 45.040 ;
        RECT 116.010 44.640 116.940 44.940 ;
        RECT 129.270 44.700 130.230 45.100 ;
        RECT 142.510 44.840 147.770 45.205 ;
        RECT 142.570 44.830 146.720 44.840 ;
        RECT 42.840 43.690 71.590 43.830 ;
        RECT 17.090 41.760 22.670 41.830 ;
        RECT 40.430 41.820 71.590 43.690 ;
        RECT 17.090 41.650 28.130 41.760 ;
        RECT 33.980 41.720 71.590 41.820 ;
        RECT 31.260 41.650 71.590 41.720 ;
        RECT 17.090 40.360 71.590 41.650 ;
        RECT 17.090 40.290 32.130 40.360 ;
        RECT 33.980 40.330 71.590 40.360 ;
        RECT 17.090 40.210 18.630 40.290 ;
        RECT 40.430 40.270 71.590 40.330 ;
        RECT 42.840 40.120 71.590 40.270 ;
        RECT 69.070 36.940 71.330 40.120 ;
        RECT 116.060 27.070 116.830 44.640 ;
        RECT 129.430 27.250 130.150 44.700 ;
        RECT 142.660 44.320 143.510 44.830 ;
        RECT 115.840 25.790 116.840 27.070 ;
        RECT 111.940 24.190 113.090 24.220 ;
        RECT 115.790 24.190 116.880 25.790 ;
        RECT 129.200 25.380 130.510 27.250 ;
        RECT 142.775 27.120 143.495 44.320 ;
        RECT 212.910 40.570 214.640 47.190 ;
        RECT 226.150 47.140 227.670 47.190 ;
        RECT 212.880 38.900 215.100 40.570 ;
        RECT 212.880 38.410 221.820 38.900 ;
        RECT 212.910 36.190 221.820 38.410 ;
        RECT 129.140 24.690 130.510 25.380 ;
        RECT 142.730 25.320 143.730 27.120 ;
        RECT 212.910 26.730 214.640 36.190 ;
        RECT 111.940 24.085 116.910 24.190 ;
        RECT 129.140 24.170 130.470 24.690 ;
        RECT 129.140 24.085 130.510 24.170 ;
        RECT 142.480 24.085 143.810 25.320 ;
        RECT 111.940 23.950 143.810 24.085 ;
        RECT 111.940 23.150 143.565 23.950 ;
        RECT 111.940 23.040 116.910 23.150 ;
        RECT 111.940 17.550 113.090 23.040 ;
        RECT 212.890 21.640 214.910 26.730 ;
        RECT 212.890 21.450 218.170 21.640 ;
        RECT 242.710 21.450 244.780 21.720 ;
        RECT 249.210 21.480 249.570 22.770 ;
        RECT 212.890 20.000 245.570 21.450 ;
        RECT 213.370 19.810 245.570 20.000 ;
        RECT 242.710 19.630 244.780 19.810 ;
        RECT 128.850 17.550 130.000 18.020 ;
        RECT 147.320 17.550 148.470 18.110 ;
        RECT 111.940 14.230 148.520 17.550 ;
        RECT 111.940 6.990 113.090 14.230 ;
        RECT 128.850 6.900 130.000 14.230 ;
        RECT 147.320 6.990 148.470 14.230 ;
        RECT 323.230 -28.090 336.720 63.420 ;
        RECT 352.930 63.350 371.180 63.420 ;
        RECT 360.450 63.330 371.180 63.350 ;
        RECT 360.450 63.300 370.760 63.330 ;
        RECT 649.750 59.320 658.940 65.510 ;
        RECT 360.860 44.510 370.050 50.660 ;
        RECT 649.750 39.320 658.940 45.510 ;
        RECT 360.860 24.510 370.050 30.660 ;
        RECT 649.750 19.320 658.940 25.510 ;
        RECT 374.170 8.920 383.360 15.150 ;
        RECT 394.170 14.650 395.110 15.130 ;
        RECT 397.810 14.650 403.360 15.130 ;
        RECT 394.170 8.920 403.360 14.650 ;
        RECT 414.170 8.920 423.360 15.130 ;
        RECT 434.170 8.920 443.360 15.130 ;
        RECT 454.170 8.920 463.360 15.130 ;
        RECT 474.170 8.920 483.360 15.130 ;
        RECT 494.170 8.920 503.360 15.130 ;
        RECT 514.170 8.920 523.360 15.130 ;
        RECT 534.170 8.920 543.360 15.130 ;
        RECT 554.170 8.920 563.360 15.130 ;
        RECT 574.170 8.920 583.360 15.130 ;
        RECT 594.170 8.920 603.360 15.130 ;
        RECT 614.170 8.920 623.360 15.130 ;
        RECT 634.170 8.920 643.360 15.130 ;
        RECT 668.840 -24.760 676.720 -24.690 ;
        RECT 738.260 -24.760 771.230 275.290 ;
        RECT 668.840 -28.090 772.700 -24.760 ;
        RECT -7.880 -40.590 772.700 -28.090 ;
        RECT -7.880 -43.920 676.720 -40.590 ;
        RECT -7.880 -44.270 8.410 -43.920 ;
        RECT 668.840 -43.940 676.720 -43.920 ;
    END
  END vssa1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 32.670 339.550 86.210 339.710 ;
        RECT 32.670 165.240 310.430 339.550 ;
        RECT 688.220 243.110 715.690 249.950 ;
        RECT 32.670 164.580 86.210 165.240 ;
        RECT 166.400 161.130 176.340 165.240 ;
        RECT 166.670 160.710 176.280 161.130 ;
        RECT 167.670 160.560 176.280 160.710 ;
        RECT 167.670 160.390 172.140 160.560 ;
        RECT 168.280 159.600 172.140 160.390 ;
        RECT 173.820 160.260 176.280 160.560 ;
        RECT 168.710 157.710 172.140 159.600 ;
        RECT 171.170 157.700 172.140 157.710 ;
        RECT 116.480 138.430 131.850 139.380 ;
        RECT 116.480 134.340 131.830 138.430 ;
        RECT 138.380 137.990 153.750 138.940 ;
        RECT 116.480 134.170 118.950 134.340 ;
        RECT 138.380 133.900 153.730 137.990 ;
        RECT 159.170 137.760 174.540 138.710 ;
        RECT 138.380 133.730 140.850 133.900 ;
        RECT 159.170 133.670 174.520 137.760 ;
        RECT 321.270 133.765 322.860 133.790 ;
        RECT 321.270 133.730 335.070 133.765 ;
        RECT 159.170 133.500 161.640 133.670 ;
        RECT 309.000 131.960 335.070 133.730 ;
        RECT 309.000 131.925 324.125 131.960 ;
        RECT 328.125 131.945 335.070 131.960 ;
        RECT 309.000 131.865 310.435 131.925 ;
        RECT 314.435 131.910 324.125 131.925 ;
        RECT 316.390 131.900 324.125 131.910 ;
        RECT 330.080 131.900 335.070 131.945 ;
        RECT 316.390 131.865 322.860 131.900 ;
        RECT 316.390 131.670 319.205 131.865 ;
        RECT 321.270 131.850 322.860 131.865 ;
        RECT 330.080 131.705 332.895 131.900 ;
        RECT 319.730 127.665 320.930 127.670 ;
        RECT 319.730 125.860 333.180 127.665 ;
        RECT 319.730 125.800 322.235 125.860 ;
        RECT 326.235 125.845 333.180 125.860 ;
        RECT 328.190 125.800 333.180 125.845 ;
        RECT 319.730 125.710 320.930 125.800 ;
        RECT 328.190 125.605 331.005 125.800 ;
        RECT 110.640 111.730 148.220 111.740 ;
        RECT 110.640 108.495 150.280 111.730 ;
        RECT 110.640 108.380 150.390 108.495 ;
        RECT 110.705 101.465 150.390 108.380 ;
        RECT 110.710 101.150 150.390 101.465 ;
        RECT 146.660 101.140 150.390 101.150 ;
        RECT 211.660 79.730 301.820 88.390 ;
        RECT 211.660 79.710 256.540 79.730 ;
        RECT 258.050 79.710 301.820 79.730 ;
        RECT 26.920 69.700 33.460 72.210 ;
        RECT 45.850 72.160 52.750 75.540 ;
        RECT 45.230 71.050 52.750 72.160 ;
        RECT 26.940 47.180 33.460 69.700 ;
        RECT 45.280 69.600 52.750 71.050 ;
        RECT 45.270 69.550 52.750 69.600 ;
        RECT 45.230 66.210 52.750 69.550 ;
        RECT 68.590 73.200 83.960 74.150 ;
        RECT 68.590 69.110 83.940 73.200 ;
        RECT 110.570 73.100 150.430 79.360 ;
        RECT 273.000 79.180 288.750 79.710 ;
        RECT 292.060 78.850 297.560 79.710 ;
        RECT 68.590 68.940 71.060 69.110 ;
        RECT 45.240 65.030 52.750 66.210 ;
        RECT 45.240 64.690 52.740 65.030 ;
        RECT 45.260 61.450 52.740 64.690 ;
        RECT 45.250 56.570 52.740 61.450 ;
        RECT 45.230 54.250 52.740 56.570 ;
        RECT 45.260 50.920 52.740 54.250 ;
        RECT 184.780 57.050 200.150 58.000 ;
        RECT 184.780 52.960 200.130 57.050 ;
        RECT 184.780 52.790 187.250 52.960 ;
        RECT 45.270 47.640 52.740 50.920 ;
        RECT 26.940 46.350 33.520 47.180 ;
        RECT 26.970 45.360 33.520 46.350 ;
        RECT 45.260 45.710 52.740 47.640 ;
        RECT 26.970 45.290 33.090 45.360 ;
        RECT 45.630 41.820 52.740 45.710 ;
        RECT 68.980 47.450 84.350 48.400 ;
        RECT 68.980 43.360 84.330 47.450 ;
        RECT 109.400 47.280 149.290 50.880 ;
        RECT 109.445 46.900 148.840 47.280 ;
        RECT 109.445 43.660 148.800 46.900 ;
        RECT 110.680 43.645 148.800 43.660 ;
        RECT 68.980 43.190 71.450 43.360 ;
        RECT 45.620 40.770 52.740 41.820 ;
        RECT 297.480 32.370 298.580 32.380 ;
        RECT 281.310 32.360 298.580 32.370 ;
        RECT 246.070 23.480 298.580 32.360 ;
        RECT 246.070 23.450 250.170 23.480 ;
        RECT 249.290 23.440 250.170 23.450 ;
        RECT 280.800 23.430 298.580 23.480 ;
        RECT 282.980 23.420 298.580 23.430 ;
        RECT 292.480 23.410 298.580 23.420 ;
        RECT 110.970 16.800 126.340 17.750 ;
        RECT 110.970 12.710 126.320 16.800 ;
        RECT 127.880 16.710 143.250 17.660 ;
        RECT 146.350 16.800 161.720 17.750 ;
        RECT 110.970 12.540 113.440 12.710 ;
        RECT 127.880 12.620 143.230 16.710 ;
        RECT 146.350 12.710 161.700 16.800 ;
        RECT 127.880 12.450 130.350 12.620 ;
        RECT 146.350 12.540 148.820 12.710 ;
        RECT 693.510 0.390 720.980 7.230 ;
      LAYER li1 ;
        RECT 39.390 322.160 44.790 327.250 ;
        RECT 46.540 323.700 46.710 330.740 ;
        RECT 54.830 323.700 55.000 330.740 ;
        RECT 63.120 323.700 63.290 330.740 ;
        RECT 39.390 312.160 44.790 317.250 ;
        RECT 46.540 315.520 46.710 322.560 ;
        RECT 54.830 315.520 55.000 322.560 ;
        RECT 63.120 315.520 63.290 322.560 ;
        RECT 65.390 322.160 70.790 327.250 ;
        RECT 72.540 323.700 72.710 330.740 ;
        RECT 80.830 323.700 81.000 330.740 ;
        RECT 89.120 323.700 89.290 330.740 ;
        RECT 46.540 307.340 46.710 314.380 ;
        RECT 54.830 307.340 55.000 314.380 ;
        RECT 63.120 307.340 63.290 314.380 ;
        RECT 65.390 312.160 70.790 317.250 ;
        RECT 72.540 315.520 72.710 322.560 ;
        RECT 80.830 315.520 81.000 322.560 ;
        RECT 89.120 315.520 89.290 322.560 ;
        RECT 91.390 322.160 96.790 327.250 ;
        RECT 98.540 323.700 98.710 330.740 ;
        RECT 106.830 323.700 107.000 330.740 ;
        RECT 115.120 323.700 115.290 330.740 ;
        RECT 72.540 307.340 72.710 314.380 ;
        RECT 80.830 307.340 81.000 314.380 ;
        RECT 89.120 307.340 89.290 314.380 ;
        RECT 91.390 312.160 96.790 317.250 ;
        RECT 98.540 315.520 98.710 322.560 ;
        RECT 106.830 315.520 107.000 322.560 ;
        RECT 115.120 315.520 115.290 322.560 ;
        RECT 117.390 322.160 122.790 327.250 ;
        RECT 124.540 323.700 124.710 330.740 ;
        RECT 132.830 323.700 133.000 330.740 ;
        RECT 141.120 323.700 141.290 330.740 ;
        RECT 98.540 307.340 98.710 314.380 ;
        RECT 106.830 307.340 107.000 314.380 ;
        RECT 115.120 307.340 115.290 314.380 ;
        RECT 117.390 312.160 122.790 317.250 ;
        RECT 124.540 315.520 124.710 322.560 ;
        RECT 132.830 315.520 133.000 322.560 ;
        RECT 141.120 315.520 141.290 322.560 ;
        RECT 143.390 322.160 148.790 327.250 ;
        RECT 150.540 323.700 150.710 330.740 ;
        RECT 158.830 323.700 159.000 330.740 ;
        RECT 167.120 323.700 167.290 330.740 ;
        RECT 124.540 307.340 124.710 314.380 ;
        RECT 132.830 307.340 133.000 314.380 ;
        RECT 141.120 307.340 141.290 314.380 ;
        RECT 143.390 312.160 148.790 317.250 ;
        RECT 150.540 315.520 150.710 322.560 ;
        RECT 158.830 315.520 159.000 322.560 ;
        RECT 167.120 315.520 167.290 322.560 ;
        RECT 169.390 322.160 174.790 327.250 ;
        RECT 176.540 323.700 176.710 330.740 ;
        RECT 184.830 323.700 185.000 330.740 ;
        RECT 193.120 323.700 193.290 330.740 ;
        RECT 150.540 307.340 150.710 314.380 ;
        RECT 158.830 307.340 159.000 314.380 ;
        RECT 167.120 307.340 167.290 314.380 ;
        RECT 169.390 312.160 174.790 317.250 ;
        RECT 176.540 315.520 176.710 322.560 ;
        RECT 184.830 315.520 185.000 322.560 ;
        RECT 193.120 315.520 193.290 322.560 ;
        RECT 195.390 322.160 200.790 327.250 ;
        RECT 202.540 323.700 202.710 330.740 ;
        RECT 210.830 323.700 211.000 330.740 ;
        RECT 219.120 323.700 219.290 330.740 ;
        RECT 176.540 307.340 176.710 314.380 ;
        RECT 184.830 307.340 185.000 314.380 ;
        RECT 193.120 307.340 193.290 314.380 ;
        RECT 195.390 312.160 200.790 317.250 ;
        RECT 202.540 315.520 202.710 322.560 ;
        RECT 210.830 315.520 211.000 322.560 ;
        RECT 219.120 315.520 219.290 322.560 ;
        RECT 221.390 322.160 226.790 327.250 ;
        RECT 228.540 323.700 228.710 330.740 ;
        RECT 236.830 323.700 237.000 330.740 ;
        RECT 245.120 323.700 245.290 330.740 ;
        RECT 202.540 307.340 202.710 314.380 ;
        RECT 210.830 307.340 211.000 314.380 ;
        RECT 219.120 307.340 219.290 314.380 ;
        RECT 221.390 312.160 226.790 317.250 ;
        RECT 228.540 315.520 228.710 322.560 ;
        RECT 236.830 315.520 237.000 322.560 ;
        RECT 245.120 315.520 245.290 322.560 ;
        RECT 247.390 322.160 252.790 327.250 ;
        RECT 254.540 323.700 254.710 330.740 ;
        RECT 262.830 323.700 263.000 330.740 ;
        RECT 271.120 323.700 271.290 330.740 ;
        RECT 228.540 307.340 228.710 314.380 ;
        RECT 236.830 307.340 237.000 314.380 ;
        RECT 245.120 307.340 245.290 314.380 ;
        RECT 247.390 312.160 252.790 317.250 ;
        RECT 254.540 315.520 254.710 322.560 ;
        RECT 262.830 315.520 263.000 322.560 ;
        RECT 271.120 315.520 271.290 322.560 ;
        RECT 273.390 322.160 278.790 327.250 ;
        RECT 280.540 323.700 280.710 330.740 ;
        RECT 288.830 323.700 289.000 330.740 ;
        RECT 297.120 323.700 297.290 330.740 ;
        RECT 254.540 307.340 254.710 314.380 ;
        RECT 262.830 307.340 263.000 314.380 ;
        RECT 271.120 307.340 271.290 314.380 ;
        RECT 273.390 312.160 278.790 317.250 ;
        RECT 280.540 315.520 280.710 322.560 ;
        RECT 288.830 315.520 289.000 322.560 ;
        RECT 297.120 315.520 297.290 322.560 ;
        RECT 299.390 322.160 304.790 327.250 ;
        RECT 280.540 307.340 280.710 314.380 ;
        RECT 288.830 307.340 289.000 314.380 ;
        RECT 297.120 307.340 297.290 314.380 ;
        RECT 299.390 312.160 304.790 317.250 ;
        RECT 39.390 302.160 44.790 307.250 ;
        RECT 46.540 299.160 46.710 306.200 ;
        RECT 54.830 299.160 55.000 306.200 ;
        RECT 63.120 299.160 63.290 306.200 ;
        RECT 65.390 302.160 70.790 307.250 ;
        RECT 72.540 299.160 72.710 306.200 ;
        RECT 80.830 299.160 81.000 306.200 ;
        RECT 89.120 299.160 89.290 306.200 ;
        RECT 91.390 302.160 96.790 307.250 ;
        RECT 98.540 299.160 98.710 306.200 ;
        RECT 106.830 299.160 107.000 306.200 ;
        RECT 115.120 299.160 115.290 306.200 ;
        RECT 117.390 302.160 122.790 307.250 ;
        RECT 124.540 299.160 124.710 306.200 ;
        RECT 132.830 299.160 133.000 306.200 ;
        RECT 141.120 299.160 141.290 306.200 ;
        RECT 143.390 302.160 148.790 307.250 ;
        RECT 150.540 299.160 150.710 306.200 ;
        RECT 158.830 299.160 159.000 306.200 ;
        RECT 167.120 299.160 167.290 306.200 ;
        RECT 169.390 302.160 174.790 307.250 ;
        RECT 176.540 299.160 176.710 306.200 ;
        RECT 184.830 299.160 185.000 306.200 ;
        RECT 193.120 299.160 193.290 306.200 ;
        RECT 195.390 302.160 200.790 307.250 ;
        RECT 202.540 299.160 202.710 306.200 ;
        RECT 210.830 299.160 211.000 306.200 ;
        RECT 219.120 299.160 219.290 306.200 ;
        RECT 221.390 302.160 226.790 307.250 ;
        RECT 228.540 299.160 228.710 306.200 ;
        RECT 236.830 299.160 237.000 306.200 ;
        RECT 245.120 299.160 245.290 306.200 ;
        RECT 247.390 302.160 252.790 307.250 ;
        RECT 254.540 299.160 254.710 306.200 ;
        RECT 262.830 299.160 263.000 306.200 ;
        RECT 271.120 299.160 271.290 306.200 ;
        RECT 273.390 302.160 278.790 307.250 ;
        RECT 280.540 299.160 280.710 306.200 ;
        RECT 288.830 299.160 289.000 306.200 ;
        RECT 297.120 299.160 297.290 306.200 ;
        RECT 299.390 302.160 304.790 307.250 ;
        RECT 39.390 292.160 44.790 297.250 ;
        RECT 46.540 290.980 46.710 298.020 ;
        RECT 54.830 290.980 55.000 298.020 ;
        RECT 63.120 290.980 63.290 298.020 ;
        RECT 65.390 292.160 70.790 297.250 ;
        RECT 72.540 290.980 72.710 298.020 ;
        RECT 80.830 290.980 81.000 298.020 ;
        RECT 89.120 290.980 89.290 298.020 ;
        RECT 91.390 292.160 96.790 297.250 ;
        RECT 98.540 290.980 98.710 298.020 ;
        RECT 106.830 290.980 107.000 298.020 ;
        RECT 115.120 290.980 115.290 298.020 ;
        RECT 117.390 292.160 122.790 297.250 ;
        RECT 124.540 290.980 124.710 298.020 ;
        RECT 132.830 290.980 133.000 298.020 ;
        RECT 141.120 290.980 141.290 298.020 ;
        RECT 143.390 292.160 148.790 297.250 ;
        RECT 150.540 290.980 150.710 298.020 ;
        RECT 158.830 290.980 159.000 298.020 ;
        RECT 167.120 290.980 167.290 298.020 ;
        RECT 169.390 292.160 174.790 297.250 ;
        RECT 176.540 290.980 176.710 298.020 ;
        RECT 184.830 290.980 185.000 298.020 ;
        RECT 193.120 290.980 193.290 298.020 ;
        RECT 195.390 292.160 200.790 297.250 ;
        RECT 202.540 290.980 202.710 298.020 ;
        RECT 210.830 290.980 211.000 298.020 ;
        RECT 219.120 290.980 219.290 298.020 ;
        RECT 221.390 292.160 226.790 297.250 ;
        RECT 228.540 290.980 228.710 298.020 ;
        RECT 236.830 290.980 237.000 298.020 ;
        RECT 245.120 290.980 245.290 298.020 ;
        RECT 247.390 292.160 252.790 297.250 ;
        RECT 254.540 290.980 254.710 298.020 ;
        RECT 262.830 290.980 263.000 298.020 ;
        RECT 271.120 290.980 271.290 298.020 ;
        RECT 273.390 292.160 278.790 297.250 ;
        RECT 280.540 290.980 280.710 298.020 ;
        RECT 288.830 290.980 289.000 298.020 ;
        RECT 297.120 290.980 297.290 298.020 ;
        RECT 299.390 292.160 304.790 297.250 ;
        RECT 39.390 282.160 44.790 287.250 ;
        RECT 46.540 282.800 46.710 289.840 ;
        RECT 54.830 282.800 55.000 289.840 ;
        RECT 63.120 282.800 63.290 289.840 ;
        RECT 65.390 282.160 70.790 287.250 ;
        RECT 72.540 282.800 72.710 289.840 ;
        RECT 80.830 282.800 81.000 289.840 ;
        RECT 89.120 282.800 89.290 289.840 ;
        RECT 91.390 282.160 96.790 287.250 ;
        RECT 98.540 282.800 98.710 289.840 ;
        RECT 106.830 282.800 107.000 289.840 ;
        RECT 115.120 282.800 115.290 289.840 ;
        RECT 117.390 282.160 122.790 287.250 ;
        RECT 124.540 282.800 124.710 289.840 ;
        RECT 132.830 282.800 133.000 289.840 ;
        RECT 141.120 282.800 141.290 289.840 ;
        RECT 143.390 282.160 148.790 287.250 ;
        RECT 150.540 282.800 150.710 289.840 ;
        RECT 158.830 282.800 159.000 289.840 ;
        RECT 167.120 282.800 167.290 289.840 ;
        RECT 169.390 282.160 174.790 287.250 ;
        RECT 176.540 282.800 176.710 289.840 ;
        RECT 184.830 282.800 185.000 289.840 ;
        RECT 193.120 282.800 193.290 289.840 ;
        RECT 195.390 282.160 200.790 287.250 ;
        RECT 202.540 282.800 202.710 289.840 ;
        RECT 210.830 282.800 211.000 289.840 ;
        RECT 219.120 282.800 219.290 289.840 ;
        RECT 221.390 282.160 226.790 287.250 ;
        RECT 228.540 282.800 228.710 289.840 ;
        RECT 236.830 282.800 237.000 289.840 ;
        RECT 245.120 282.800 245.290 289.840 ;
        RECT 247.390 282.160 252.790 287.250 ;
        RECT 254.540 282.800 254.710 289.840 ;
        RECT 262.830 282.800 263.000 289.840 ;
        RECT 271.120 282.800 271.290 289.840 ;
        RECT 273.390 282.160 278.790 287.250 ;
        RECT 280.540 282.800 280.710 289.840 ;
        RECT 288.830 282.800 289.000 289.840 ;
        RECT 297.120 282.800 297.290 289.840 ;
        RECT 299.390 282.160 304.790 287.250 ;
        RECT 39.390 272.160 44.790 277.250 ;
        RECT 46.540 274.620 46.710 281.660 ;
        RECT 54.830 274.620 55.000 281.660 ;
        RECT 63.120 274.620 63.290 281.660 ;
        RECT 39.390 262.160 44.790 267.250 ;
        RECT 46.540 266.440 46.710 273.480 ;
        RECT 54.830 266.440 55.000 273.480 ;
        RECT 63.120 266.440 63.290 273.480 ;
        RECT 65.390 272.160 70.790 277.250 ;
        RECT 72.540 274.620 72.710 281.660 ;
        RECT 80.830 274.620 81.000 281.660 ;
        RECT 89.120 274.620 89.290 281.660 ;
        RECT 46.540 258.260 46.710 265.300 ;
        RECT 54.830 258.260 55.000 265.300 ;
        RECT 63.120 258.260 63.290 265.300 ;
        RECT 65.390 262.160 70.790 267.250 ;
        RECT 72.540 266.440 72.710 273.480 ;
        RECT 80.830 266.440 81.000 273.480 ;
        RECT 89.120 266.440 89.290 273.480 ;
        RECT 91.390 272.160 96.790 277.250 ;
        RECT 98.540 274.620 98.710 281.660 ;
        RECT 106.830 274.620 107.000 281.660 ;
        RECT 115.120 274.620 115.290 281.660 ;
        RECT 72.540 258.260 72.710 265.300 ;
        RECT 80.830 258.260 81.000 265.300 ;
        RECT 89.120 258.260 89.290 265.300 ;
        RECT 91.390 262.160 96.790 267.250 ;
        RECT 98.540 266.440 98.710 273.480 ;
        RECT 106.830 266.440 107.000 273.480 ;
        RECT 115.120 266.440 115.290 273.480 ;
        RECT 117.390 272.160 122.790 277.250 ;
        RECT 124.540 274.620 124.710 281.660 ;
        RECT 132.830 274.620 133.000 281.660 ;
        RECT 141.120 274.620 141.290 281.660 ;
        RECT 98.540 258.260 98.710 265.300 ;
        RECT 106.830 258.260 107.000 265.300 ;
        RECT 115.120 258.260 115.290 265.300 ;
        RECT 117.390 262.160 122.790 267.250 ;
        RECT 124.540 266.440 124.710 273.480 ;
        RECT 132.830 266.440 133.000 273.480 ;
        RECT 141.120 266.440 141.290 273.480 ;
        RECT 143.390 272.160 148.790 277.250 ;
        RECT 150.540 274.620 150.710 281.660 ;
        RECT 158.830 274.620 159.000 281.660 ;
        RECT 167.120 274.620 167.290 281.660 ;
        RECT 124.540 258.260 124.710 265.300 ;
        RECT 132.830 258.260 133.000 265.300 ;
        RECT 141.120 258.260 141.290 265.300 ;
        RECT 143.390 262.160 148.790 267.250 ;
        RECT 150.540 266.440 150.710 273.480 ;
        RECT 158.830 266.440 159.000 273.480 ;
        RECT 167.120 266.440 167.290 273.480 ;
        RECT 169.390 272.160 174.790 277.250 ;
        RECT 176.540 274.620 176.710 281.660 ;
        RECT 184.830 274.620 185.000 281.660 ;
        RECT 193.120 274.620 193.290 281.660 ;
        RECT 150.540 258.260 150.710 265.300 ;
        RECT 158.830 258.260 159.000 265.300 ;
        RECT 167.120 258.260 167.290 265.300 ;
        RECT 169.390 262.160 174.790 267.250 ;
        RECT 176.540 266.440 176.710 273.480 ;
        RECT 184.830 266.440 185.000 273.480 ;
        RECT 193.120 266.440 193.290 273.480 ;
        RECT 195.390 272.160 200.790 277.250 ;
        RECT 202.540 274.620 202.710 281.660 ;
        RECT 210.830 274.620 211.000 281.660 ;
        RECT 219.120 274.620 219.290 281.660 ;
        RECT 176.540 258.260 176.710 265.300 ;
        RECT 184.830 258.260 185.000 265.300 ;
        RECT 193.120 258.260 193.290 265.300 ;
        RECT 195.390 262.160 200.790 267.250 ;
        RECT 202.540 266.440 202.710 273.480 ;
        RECT 210.830 266.440 211.000 273.480 ;
        RECT 219.120 266.440 219.290 273.480 ;
        RECT 221.390 272.160 226.790 277.250 ;
        RECT 228.540 274.620 228.710 281.660 ;
        RECT 236.830 274.620 237.000 281.660 ;
        RECT 245.120 274.620 245.290 281.660 ;
        RECT 202.540 258.260 202.710 265.300 ;
        RECT 210.830 258.260 211.000 265.300 ;
        RECT 219.120 258.260 219.290 265.300 ;
        RECT 221.390 262.160 226.790 267.250 ;
        RECT 228.540 266.440 228.710 273.480 ;
        RECT 236.830 266.440 237.000 273.480 ;
        RECT 245.120 266.440 245.290 273.480 ;
        RECT 247.390 272.160 252.790 277.250 ;
        RECT 254.540 274.620 254.710 281.660 ;
        RECT 262.830 274.620 263.000 281.660 ;
        RECT 271.120 274.620 271.290 281.660 ;
        RECT 228.540 258.260 228.710 265.300 ;
        RECT 236.830 258.260 237.000 265.300 ;
        RECT 245.120 258.260 245.290 265.300 ;
        RECT 247.390 262.160 252.790 267.250 ;
        RECT 254.540 266.440 254.710 273.480 ;
        RECT 262.830 266.440 263.000 273.480 ;
        RECT 271.120 266.440 271.290 273.480 ;
        RECT 273.390 272.160 278.790 277.250 ;
        RECT 280.540 274.620 280.710 281.660 ;
        RECT 288.830 274.620 289.000 281.660 ;
        RECT 297.120 274.620 297.290 281.660 ;
        RECT 254.540 258.260 254.710 265.300 ;
        RECT 262.830 258.260 263.000 265.300 ;
        RECT 271.120 258.260 271.290 265.300 ;
        RECT 273.390 262.160 278.790 267.250 ;
        RECT 280.540 266.440 280.710 273.480 ;
        RECT 288.830 266.440 289.000 273.480 ;
        RECT 297.120 266.440 297.290 273.480 ;
        RECT 299.390 272.160 304.790 277.250 ;
        RECT 280.540 258.260 280.710 265.300 ;
        RECT 288.830 258.260 289.000 265.300 ;
        RECT 297.120 258.260 297.290 265.300 ;
        RECT 299.390 262.160 304.790 267.250 ;
        RECT 39.390 252.160 44.790 257.250 ;
        RECT 46.540 250.080 46.710 257.120 ;
        RECT 54.830 250.080 55.000 257.120 ;
        RECT 63.120 250.080 63.290 257.120 ;
        RECT 65.390 252.160 70.790 257.250 ;
        RECT 72.540 250.080 72.710 257.120 ;
        RECT 80.830 250.080 81.000 257.120 ;
        RECT 89.120 250.080 89.290 257.120 ;
        RECT 91.390 252.160 96.790 257.250 ;
        RECT 98.540 250.080 98.710 257.120 ;
        RECT 106.830 250.080 107.000 257.120 ;
        RECT 115.120 250.080 115.290 257.120 ;
        RECT 117.390 252.160 122.790 257.250 ;
        RECT 124.540 250.080 124.710 257.120 ;
        RECT 132.830 250.080 133.000 257.120 ;
        RECT 141.120 250.080 141.290 257.120 ;
        RECT 143.390 252.160 148.790 257.250 ;
        RECT 150.540 250.080 150.710 257.120 ;
        RECT 158.830 250.080 159.000 257.120 ;
        RECT 167.120 250.080 167.290 257.120 ;
        RECT 169.390 252.160 174.790 257.250 ;
        RECT 176.540 250.080 176.710 257.120 ;
        RECT 184.830 250.080 185.000 257.120 ;
        RECT 193.120 250.080 193.290 257.120 ;
        RECT 195.390 252.160 200.790 257.250 ;
        RECT 202.540 250.080 202.710 257.120 ;
        RECT 210.830 250.080 211.000 257.120 ;
        RECT 219.120 250.080 219.290 257.120 ;
        RECT 221.390 252.160 226.790 257.250 ;
        RECT 228.540 250.080 228.710 257.120 ;
        RECT 236.830 250.080 237.000 257.120 ;
        RECT 245.120 250.080 245.290 257.120 ;
        RECT 247.390 252.160 252.790 257.250 ;
        RECT 254.540 250.080 254.710 257.120 ;
        RECT 262.830 250.080 263.000 257.120 ;
        RECT 271.120 250.080 271.290 257.120 ;
        RECT 273.390 252.160 278.790 257.250 ;
        RECT 280.540 250.080 280.710 257.120 ;
        RECT 288.830 250.080 289.000 257.120 ;
        RECT 297.120 250.080 297.290 257.120 ;
        RECT 299.390 252.160 304.790 257.250 ;
        RECT 688.400 249.600 715.510 249.770 ;
        RECT 39.390 240.160 44.790 245.250 ;
        RECT 46.540 241.900 46.710 248.940 ;
        RECT 54.830 241.900 55.000 248.940 ;
        RECT 63.120 241.900 63.290 248.940 ;
        RECT 39.390 230.160 44.790 235.250 ;
        RECT 46.540 233.720 46.710 240.760 ;
        RECT 54.830 233.720 55.000 240.760 ;
        RECT 63.120 233.720 63.290 240.760 ;
        RECT 65.390 240.160 70.790 245.250 ;
        RECT 72.540 241.900 72.710 248.940 ;
        RECT 80.830 241.900 81.000 248.940 ;
        RECT 89.120 241.900 89.290 248.940 ;
        RECT 46.540 225.540 46.710 232.580 ;
        RECT 54.830 225.540 55.000 232.580 ;
        RECT 63.120 225.540 63.290 232.580 ;
        RECT 65.390 230.160 70.790 235.250 ;
        RECT 72.540 233.720 72.710 240.760 ;
        RECT 80.830 233.720 81.000 240.760 ;
        RECT 89.120 233.720 89.290 240.760 ;
        RECT 91.390 240.160 96.790 245.250 ;
        RECT 98.540 241.900 98.710 248.940 ;
        RECT 106.830 241.900 107.000 248.940 ;
        RECT 115.120 241.900 115.290 248.940 ;
        RECT 72.540 225.540 72.710 232.580 ;
        RECT 80.830 225.540 81.000 232.580 ;
        RECT 89.120 225.540 89.290 232.580 ;
        RECT 91.390 230.160 96.790 235.250 ;
        RECT 98.540 233.720 98.710 240.760 ;
        RECT 106.830 233.720 107.000 240.760 ;
        RECT 115.120 233.720 115.290 240.760 ;
        RECT 117.390 240.160 122.790 245.250 ;
        RECT 124.540 241.900 124.710 248.940 ;
        RECT 132.830 241.900 133.000 248.940 ;
        RECT 141.120 241.900 141.290 248.940 ;
        RECT 98.540 225.540 98.710 232.580 ;
        RECT 106.830 225.540 107.000 232.580 ;
        RECT 115.120 225.540 115.290 232.580 ;
        RECT 117.390 230.160 122.790 235.250 ;
        RECT 124.540 233.720 124.710 240.760 ;
        RECT 132.830 233.720 133.000 240.760 ;
        RECT 141.120 233.720 141.290 240.760 ;
        RECT 143.390 240.160 148.790 245.250 ;
        RECT 150.540 241.900 150.710 248.940 ;
        RECT 158.830 241.900 159.000 248.940 ;
        RECT 167.120 241.900 167.290 248.940 ;
        RECT 124.540 225.540 124.710 232.580 ;
        RECT 132.830 225.540 133.000 232.580 ;
        RECT 141.120 225.540 141.290 232.580 ;
        RECT 143.390 230.160 148.790 235.250 ;
        RECT 150.540 233.720 150.710 240.760 ;
        RECT 158.830 233.720 159.000 240.760 ;
        RECT 167.120 233.720 167.290 240.760 ;
        RECT 169.390 240.160 174.790 245.250 ;
        RECT 176.540 241.900 176.710 248.940 ;
        RECT 184.830 241.900 185.000 248.940 ;
        RECT 193.120 241.900 193.290 248.940 ;
        RECT 150.540 225.540 150.710 232.580 ;
        RECT 158.830 225.540 159.000 232.580 ;
        RECT 167.120 225.540 167.290 232.580 ;
        RECT 169.390 230.160 174.790 235.250 ;
        RECT 176.540 233.720 176.710 240.760 ;
        RECT 184.830 233.720 185.000 240.760 ;
        RECT 193.120 233.720 193.290 240.760 ;
        RECT 195.390 240.160 200.790 245.250 ;
        RECT 202.540 241.900 202.710 248.940 ;
        RECT 210.830 241.900 211.000 248.940 ;
        RECT 219.120 241.900 219.290 248.940 ;
        RECT 176.540 225.540 176.710 232.580 ;
        RECT 184.830 225.540 185.000 232.580 ;
        RECT 193.120 225.540 193.290 232.580 ;
        RECT 195.390 230.160 200.790 235.250 ;
        RECT 202.540 233.720 202.710 240.760 ;
        RECT 210.830 233.720 211.000 240.760 ;
        RECT 219.120 233.720 219.290 240.760 ;
        RECT 221.390 240.160 226.790 245.250 ;
        RECT 228.540 241.900 228.710 248.940 ;
        RECT 236.830 241.900 237.000 248.940 ;
        RECT 245.120 241.900 245.290 248.940 ;
        RECT 202.540 225.540 202.710 232.580 ;
        RECT 210.830 225.540 211.000 232.580 ;
        RECT 219.120 225.540 219.290 232.580 ;
        RECT 221.390 230.160 226.790 235.250 ;
        RECT 228.540 233.720 228.710 240.760 ;
        RECT 236.830 233.720 237.000 240.760 ;
        RECT 245.120 233.720 245.290 240.760 ;
        RECT 247.390 240.160 252.790 245.250 ;
        RECT 254.540 241.900 254.710 248.940 ;
        RECT 262.830 241.900 263.000 248.940 ;
        RECT 271.120 241.900 271.290 248.940 ;
        RECT 228.540 225.540 228.710 232.580 ;
        RECT 236.830 225.540 237.000 232.580 ;
        RECT 245.120 225.540 245.290 232.580 ;
        RECT 247.390 230.160 252.790 235.250 ;
        RECT 254.540 233.720 254.710 240.760 ;
        RECT 262.830 233.720 263.000 240.760 ;
        RECT 271.120 233.720 271.290 240.760 ;
        RECT 273.390 240.160 278.790 245.250 ;
        RECT 280.540 241.900 280.710 248.940 ;
        RECT 288.830 241.900 289.000 248.940 ;
        RECT 297.120 241.900 297.290 248.940 ;
        RECT 254.540 225.540 254.710 232.580 ;
        RECT 262.830 225.540 263.000 232.580 ;
        RECT 271.120 225.540 271.290 232.580 ;
        RECT 273.390 230.160 278.790 235.250 ;
        RECT 280.540 233.720 280.710 240.760 ;
        RECT 288.830 233.720 289.000 240.760 ;
        RECT 297.120 233.720 297.290 240.760 ;
        RECT 299.390 240.160 304.790 245.250 ;
        RECT 688.400 243.460 688.570 249.600 ;
        RECT 690.260 243.975 690.430 249.230 ;
        RECT 692.840 243.975 693.010 249.230 ;
        RECT 695.420 243.975 695.590 249.230 ;
        RECT 698.000 243.975 698.170 249.230 ;
        RECT 700.580 243.975 700.750 249.230 ;
        RECT 703.160 243.975 703.330 249.230 ;
        RECT 705.740 243.975 705.910 249.230 ;
        RECT 708.320 243.975 708.490 249.230 ;
        RECT 710.900 243.975 711.070 249.230 ;
        RECT 713.480 243.975 713.650 249.230 ;
        RECT 688.970 243.805 714.940 243.975 ;
        RECT 715.340 243.460 715.510 249.600 ;
        RECT 688.400 243.290 715.510 243.460 ;
        RECT 280.540 225.540 280.710 232.580 ;
        RECT 288.830 225.540 289.000 232.580 ;
        RECT 297.120 225.540 297.290 232.580 ;
        RECT 299.390 230.160 304.790 235.250 ;
        RECT 39.390 220.160 44.790 225.250 ;
        RECT 46.540 217.360 46.710 224.400 ;
        RECT 54.830 217.360 55.000 224.400 ;
        RECT 63.120 217.360 63.290 224.400 ;
        RECT 65.390 220.160 70.790 225.250 ;
        RECT 72.540 217.360 72.710 224.400 ;
        RECT 80.830 217.360 81.000 224.400 ;
        RECT 89.120 217.360 89.290 224.400 ;
        RECT 91.390 220.160 96.790 225.250 ;
        RECT 98.540 217.360 98.710 224.400 ;
        RECT 106.830 217.360 107.000 224.400 ;
        RECT 115.120 217.360 115.290 224.400 ;
        RECT 117.390 220.160 122.790 225.250 ;
        RECT 124.540 217.360 124.710 224.400 ;
        RECT 132.830 217.360 133.000 224.400 ;
        RECT 141.120 217.360 141.290 224.400 ;
        RECT 143.390 220.160 148.790 225.250 ;
        RECT 150.540 217.360 150.710 224.400 ;
        RECT 158.830 217.360 159.000 224.400 ;
        RECT 167.120 217.360 167.290 224.400 ;
        RECT 169.390 220.160 174.790 225.250 ;
        RECT 176.540 217.360 176.710 224.400 ;
        RECT 184.830 217.360 185.000 224.400 ;
        RECT 193.120 217.360 193.290 224.400 ;
        RECT 195.390 220.160 200.790 225.250 ;
        RECT 202.540 217.360 202.710 224.400 ;
        RECT 210.830 217.360 211.000 224.400 ;
        RECT 219.120 217.360 219.290 224.400 ;
        RECT 221.390 220.160 226.790 225.250 ;
        RECT 228.540 217.360 228.710 224.400 ;
        RECT 236.830 217.360 237.000 224.400 ;
        RECT 245.120 217.360 245.290 224.400 ;
        RECT 247.390 220.160 252.790 225.250 ;
        RECT 254.540 217.360 254.710 224.400 ;
        RECT 262.830 217.360 263.000 224.400 ;
        RECT 271.120 217.360 271.290 224.400 ;
        RECT 273.390 220.160 278.790 225.250 ;
        RECT 280.540 217.360 280.710 224.400 ;
        RECT 288.830 217.360 289.000 224.400 ;
        RECT 297.120 217.360 297.290 224.400 ;
        RECT 299.390 220.160 304.790 225.250 ;
        RECT 39.390 210.160 44.790 215.250 ;
        RECT 46.540 209.180 46.710 216.220 ;
        RECT 54.830 209.180 55.000 216.220 ;
        RECT 63.120 209.180 63.290 216.220 ;
        RECT 65.390 210.160 70.790 215.250 ;
        RECT 72.540 209.180 72.710 216.220 ;
        RECT 80.830 209.180 81.000 216.220 ;
        RECT 89.120 209.180 89.290 216.220 ;
        RECT 91.390 210.160 96.790 215.250 ;
        RECT 98.540 209.180 98.710 216.220 ;
        RECT 106.830 209.180 107.000 216.220 ;
        RECT 115.120 209.180 115.290 216.220 ;
        RECT 117.390 210.160 122.790 215.250 ;
        RECT 124.540 209.180 124.710 216.220 ;
        RECT 132.830 209.180 133.000 216.220 ;
        RECT 141.120 209.180 141.290 216.220 ;
        RECT 143.390 210.160 148.790 215.250 ;
        RECT 150.540 209.180 150.710 216.220 ;
        RECT 158.830 209.180 159.000 216.220 ;
        RECT 167.120 209.180 167.290 216.220 ;
        RECT 169.390 210.160 174.790 215.250 ;
        RECT 176.540 209.180 176.710 216.220 ;
        RECT 184.830 209.180 185.000 216.220 ;
        RECT 193.120 209.180 193.290 216.220 ;
        RECT 195.390 210.160 200.790 215.250 ;
        RECT 202.540 209.180 202.710 216.220 ;
        RECT 210.830 209.180 211.000 216.220 ;
        RECT 219.120 209.180 219.290 216.220 ;
        RECT 221.390 210.160 226.790 215.250 ;
        RECT 228.540 209.180 228.710 216.220 ;
        RECT 236.830 209.180 237.000 216.220 ;
        RECT 245.120 209.180 245.290 216.220 ;
        RECT 247.390 210.160 252.790 215.250 ;
        RECT 254.540 209.180 254.710 216.220 ;
        RECT 262.830 209.180 263.000 216.220 ;
        RECT 271.120 209.180 271.290 216.220 ;
        RECT 273.390 210.160 278.790 215.250 ;
        RECT 280.540 209.180 280.710 216.220 ;
        RECT 288.830 209.180 289.000 216.220 ;
        RECT 297.120 209.180 297.290 216.220 ;
        RECT 299.390 210.160 304.790 215.250 ;
        RECT 39.390 200.160 44.790 205.250 ;
        RECT 46.540 201.000 46.710 208.040 ;
        RECT 54.830 201.000 55.000 208.040 ;
        RECT 63.120 201.000 63.290 208.040 ;
        RECT 65.390 200.160 70.790 205.250 ;
        RECT 72.540 201.000 72.710 208.040 ;
        RECT 80.830 201.000 81.000 208.040 ;
        RECT 89.120 201.000 89.290 208.040 ;
        RECT 91.390 200.160 96.790 205.250 ;
        RECT 98.540 201.000 98.710 208.040 ;
        RECT 106.830 201.000 107.000 208.040 ;
        RECT 115.120 201.000 115.290 208.040 ;
        RECT 117.390 200.160 122.790 205.250 ;
        RECT 124.540 201.000 124.710 208.040 ;
        RECT 132.830 201.000 133.000 208.040 ;
        RECT 141.120 201.000 141.290 208.040 ;
        RECT 143.390 200.160 148.790 205.250 ;
        RECT 150.540 201.000 150.710 208.040 ;
        RECT 158.830 201.000 159.000 208.040 ;
        RECT 167.120 201.000 167.290 208.040 ;
        RECT 169.390 200.160 174.790 205.250 ;
        RECT 176.540 201.000 176.710 208.040 ;
        RECT 184.830 201.000 185.000 208.040 ;
        RECT 193.120 201.000 193.290 208.040 ;
        RECT 195.390 200.160 200.790 205.250 ;
        RECT 202.540 201.000 202.710 208.040 ;
        RECT 210.830 201.000 211.000 208.040 ;
        RECT 219.120 201.000 219.290 208.040 ;
        RECT 221.390 200.160 226.790 205.250 ;
        RECT 228.540 201.000 228.710 208.040 ;
        RECT 236.830 201.000 237.000 208.040 ;
        RECT 245.120 201.000 245.290 208.040 ;
        RECT 247.390 200.160 252.790 205.250 ;
        RECT 254.540 201.000 254.710 208.040 ;
        RECT 262.830 201.000 263.000 208.040 ;
        RECT 271.120 201.000 271.290 208.040 ;
        RECT 273.390 200.160 278.790 205.250 ;
        RECT 280.540 201.000 280.710 208.040 ;
        RECT 288.830 201.000 289.000 208.040 ;
        RECT 297.120 201.000 297.290 208.040 ;
        RECT 299.390 200.160 304.790 205.250 ;
        RECT 39.390 190.160 44.790 195.250 ;
        RECT 46.540 192.820 46.710 199.860 ;
        RECT 54.830 192.820 55.000 199.860 ;
        RECT 63.120 192.820 63.290 199.860 ;
        RECT 39.390 180.160 44.790 185.250 ;
        RECT 46.540 184.640 46.710 191.680 ;
        RECT 54.830 184.640 55.000 191.680 ;
        RECT 63.120 184.640 63.290 191.680 ;
        RECT 65.390 190.160 70.790 195.250 ;
        RECT 72.540 192.820 72.710 199.860 ;
        RECT 80.830 192.820 81.000 199.860 ;
        RECT 89.120 192.820 89.290 199.860 ;
        RECT 46.540 176.460 46.710 183.500 ;
        RECT 54.830 176.460 55.000 183.500 ;
        RECT 63.120 176.460 63.290 183.500 ;
        RECT 65.390 180.160 70.790 185.250 ;
        RECT 72.540 184.640 72.710 191.680 ;
        RECT 80.830 184.640 81.000 191.680 ;
        RECT 89.120 184.640 89.290 191.680 ;
        RECT 91.390 190.160 96.790 195.250 ;
        RECT 98.540 192.820 98.710 199.860 ;
        RECT 106.830 192.820 107.000 199.860 ;
        RECT 115.120 192.820 115.290 199.860 ;
        RECT 72.540 176.460 72.710 183.500 ;
        RECT 80.830 176.460 81.000 183.500 ;
        RECT 89.120 176.460 89.290 183.500 ;
        RECT 91.390 180.160 96.790 185.250 ;
        RECT 98.540 184.640 98.710 191.680 ;
        RECT 106.830 184.640 107.000 191.680 ;
        RECT 115.120 184.640 115.290 191.680 ;
        RECT 117.390 190.160 122.790 195.250 ;
        RECT 124.540 192.820 124.710 199.860 ;
        RECT 132.830 192.820 133.000 199.860 ;
        RECT 141.120 192.820 141.290 199.860 ;
        RECT 98.540 176.460 98.710 183.500 ;
        RECT 106.830 176.460 107.000 183.500 ;
        RECT 115.120 176.460 115.290 183.500 ;
        RECT 117.390 180.160 122.790 185.250 ;
        RECT 124.540 184.640 124.710 191.680 ;
        RECT 132.830 184.640 133.000 191.680 ;
        RECT 141.120 184.640 141.290 191.680 ;
        RECT 143.390 190.160 148.790 195.250 ;
        RECT 150.540 192.820 150.710 199.860 ;
        RECT 158.830 192.820 159.000 199.860 ;
        RECT 167.120 192.820 167.290 199.860 ;
        RECT 124.540 176.460 124.710 183.500 ;
        RECT 132.830 176.460 133.000 183.500 ;
        RECT 141.120 176.460 141.290 183.500 ;
        RECT 143.390 180.160 148.790 185.250 ;
        RECT 150.540 184.640 150.710 191.680 ;
        RECT 158.830 184.640 159.000 191.680 ;
        RECT 167.120 184.640 167.290 191.680 ;
        RECT 169.390 190.160 174.790 195.250 ;
        RECT 176.540 192.820 176.710 199.860 ;
        RECT 184.830 192.820 185.000 199.860 ;
        RECT 193.120 192.820 193.290 199.860 ;
        RECT 150.540 176.460 150.710 183.500 ;
        RECT 158.830 176.460 159.000 183.500 ;
        RECT 167.120 176.460 167.290 183.500 ;
        RECT 169.390 180.160 174.790 185.250 ;
        RECT 176.540 184.640 176.710 191.680 ;
        RECT 184.830 184.640 185.000 191.680 ;
        RECT 193.120 184.640 193.290 191.680 ;
        RECT 195.390 190.160 200.790 195.250 ;
        RECT 202.540 192.820 202.710 199.860 ;
        RECT 210.830 192.820 211.000 199.860 ;
        RECT 219.120 192.820 219.290 199.860 ;
        RECT 176.540 176.460 176.710 183.500 ;
        RECT 184.830 176.460 185.000 183.500 ;
        RECT 193.120 176.460 193.290 183.500 ;
        RECT 195.390 180.160 200.790 185.250 ;
        RECT 202.540 184.640 202.710 191.680 ;
        RECT 210.830 184.640 211.000 191.680 ;
        RECT 219.120 184.640 219.290 191.680 ;
        RECT 221.390 190.160 226.790 195.250 ;
        RECT 228.540 192.820 228.710 199.860 ;
        RECT 236.830 192.820 237.000 199.860 ;
        RECT 245.120 192.820 245.290 199.860 ;
        RECT 202.540 176.460 202.710 183.500 ;
        RECT 210.830 176.460 211.000 183.500 ;
        RECT 219.120 176.460 219.290 183.500 ;
        RECT 221.390 180.160 226.790 185.250 ;
        RECT 228.540 184.640 228.710 191.680 ;
        RECT 236.830 184.640 237.000 191.680 ;
        RECT 245.120 184.640 245.290 191.680 ;
        RECT 247.390 190.160 252.790 195.250 ;
        RECT 254.540 192.820 254.710 199.860 ;
        RECT 262.830 192.820 263.000 199.860 ;
        RECT 271.120 192.820 271.290 199.860 ;
        RECT 228.540 176.460 228.710 183.500 ;
        RECT 236.830 176.460 237.000 183.500 ;
        RECT 245.120 176.460 245.290 183.500 ;
        RECT 247.390 180.160 252.790 185.250 ;
        RECT 254.540 184.640 254.710 191.680 ;
        RECT 262.830 184.640 263.000 191.680 ;
        RECT 271.120 184.640 271.290 191.680 ;
        RECT 273.390 190.160 278.790 195.250 ;
        RECT 280.540 192.820 280.710 199.860 ;
        RECT 288.830 192.820 289.000 199.860 ;
        RECT 297.120 192.820 297.290 199.860 ;
        RECT 254.540 176.460 254.710 183.500 ;
        RECT 262.830 176.460 263.000 183.500 ;
        RECT 271.120 176.460 271.290 183.500 ;
        RECT 273.390 180.160 278.790 185.250 ;
        RECT 280.540 184.640 280.710 191.680 ;
        RECT 288.830 184.640 289.000 191.680 ;
        RECT 297.120 184.640 297.290 191.680 ;
        RECT 299.390 190.160 304.790 195.250 ;
        RECT 280.540 176.460 280.710 183.500 ;
        RECT 288.830 176.460 289.000 183.500 ;
        RECT 297.120 176.460 297.290 183.500 ;
        RECT 299.390 180.160 304.790 185.250 ;
        RECT 39.390 170.160 44.790 175.250 ;
        RECT 46.540 168.280 46.710 175.320 ;
        RECT 54.830 168.280 55.000 175.320 ;
        RECT 63.120 168.280 63.290 175.320 ;
        RECT 65.390 170.160 70.790 175.250 ;
        RECT 72.540 168.280 72.710 175.320 ;
        RECT 80.830 168.280 81.000 175.320 ;
        RECT 89.120 168.280 89.290 175.320 ;
        RECT 91.390 170.160 96.790 175.250 ;
        RECT 98.540 168.280 98.710 175.320 ;
        RECT 106.830 168.280 107.000 175.320 ;
        RECT 115.120 168.280 115.290 175.320 ;
        RECT 117.390 170.160 122.790 175.250 ;
        RECT 124.540 168.280 124.710 175.320 ;
        RECT 132.830 168.280 133.000 175.320 ;
        RECT 141.120 168.280 141.290 175.320 ;
        RECT 143.390 170.160 148.790 175.250 ;
        RECT 150.540 168.280 150.710 175.320 ;
        RECT 158.830 168.280 159.000 175.320 ;
        RECT 167.120 168.280 167.290 175.320 ;
        RECT 169.390 170.160 174.790 175.250 ;
        RECT 176.540 168.280 176.710 175.320 ;
        RECT 184.830 168.280 185.000 175.320 ;
        RECT 193.120 168.280 193.290 175.320 ;
        RECT 195.390 170.160 200.790 175.250 ;
        RECT 202.540 168.280 202.710 175.320 ;
        RECT 210.830 168.280 211.000 175.320 ;
        RECT 219.120 168.280 219.290 175.320 ;
        RECT 221.390 170.160 226.790 175.250 ;
        RECT 228.540 168.280 228.710 175.320 ;
        RECT 236.830 168.280 237.000 175.320 ;
        RECT 245.120 168.280 245.290 175.320 ;
        RECT 247.390 170.160 252.790 175.250 ;
        RECT 254.540 168.280 254.710 175.320 ;
        RECT 262.830 168.280 263.000 175.320 ;
        RECT 271.120 168.280 271.290 175.320 ;
        RECT 273.390 170.160 278.790 175.250 ;
        RECT 280.540 168.280 280.710 175.320 ;
        RECT 288.830 168.280 289.000 175.320 ;
        RECT 297.120 168.280 297.290 175.320 ;
        RECT 299.390 170.160 304.790 175.250 ;
        RECT 124.440 139.130 126.160 139.740 ;
        RECT 147.800 139.590 168.440 139.650 ;
        RECT 127.960 139.130 168.440 139.590 ;
        RECT 118.370 139.080 168.440 139.130 ;
        RECT 118.350 139.070 168.440 139.080 ;
        RECT 118.350 138.580 168.850 139.070 ;
        RECT 118.350 138.130 118.890 138.580 ;
        RECT 127.960 138.460 168.850 138.580 ;
        RECT 118.350 135.460 118.910 138.130 ;
        RECT 127.960 138.060 171.980 138.460 ;
        RECT 127.960 138.000 148.180 138.060 ;
        RECT 128.680 136.670 128.900 138.000 ;
        RECT 129.120 136.670 129.290 136.680 ;
        RECT 128.680 135.790 129.340 136.670 ;
        RECT 129.120 135.740 129.290 135.790 ;
        RECT 132.860 117.000 134.640 138.000 ;
        RECT 140.250 137.690 140.790 138.000 ;
        RECT 140.250 135.020 140.810 137.690 ;
        RECT 150.580 136.230 150.800 138.060 ;
        RECT 158.570 137.910 171.980 138.060 ;
        RECT 158.570 137.470 168.440 137.910 ;
        RECT 171.180 137.900 171.970 137.910 ;
        RECT 161.040 136.840 162.270 137.470 ;
        RECT 151.020 136.230 151.190 136.240 ;
        RECT 150.580 135.350 151.240 136.230 ;
        RECT 151.020 135.300 151.190 135.350 ;
        RECT 161.040 134.790 161.600 136.840 ;
        RECT 171.370 136.000 171.590 137.900 ;
        RECT 171.810 136.000 171.980 136.010 ;
        RECT 171.370 135.120 172.030 136.000 ;
        RECT 171.810 135.070 171.980 135.120 ;
        RECT 309.190 133.455 321.190 133.625 ;
        RECT 322.170 133.490 334.880 133.660 ;
        RECT 309.740 132.545 310.070 133.455 ;
        RECT 311.180 132.875 311.530 133.455 ;
        RECT 313.550 132.860 313.880 133.455 ;
        RECT 314.560 132.450 314.890 133.455 ;
        RECT 316.535 132.735 317.215 133.455 ;
        RECT 317.875 132.150 318.205 133.455 ;
        RECT 318.815 131.830 319.065 133.455 ;
        RECT 319.790 132.025 320.145 133.455 ;
        RECT 320.770 132.025 321.065 133.455 ;
        RECT 322.170 133.150 322.520 133.490 ;
        RECT 322.030 132.670 322.600 133.150 ;
        RECT 323.430 132.580 323.760 133.490 ;
        RECT 324.870 132.910 325.220 133.490 ;
        RECT 327.240 132.895 327.570 133.490 ;
        RECT 328.250 132.485 328.580 133.490 ;
        RECT 330.225 132.770 330.905 133.490 ;
        RECT 331.565 132.185 331.895 133.490 ;
        RECT 332.505 131.865 332.755 133.490 ;
        RECT 333.480 132.060 333.835 133.490 ;
        RECT 334.460 132.060 334.755 133.490 ;
        RECT 320.060 127.560 320.730 127.580 ;
        RECT 320.060 127.390 332.990 127.560 ;
        RECT 320.060 127.370 321.200 127.390 ;
        RECT 320.060 126.390 320.730 127.370 ;
        RECT 321.540 126.480 321.870 127.390 ;
        RECT 322.980 126.810 323.330 127.390 ;
        RECT 325.350 126.795 325.680 127.390 ;
        RECT 326.360 126.385 326.690 127.390 ;
        RECT 328.335 126.670 329.015 127.390 ;
        RECT 329.675 126.085 330.005 127.390 ;
        RECT 330.615 125.765 330.865 127.390 ;
        RECT 331.590 125.960 331.945 127.390 ;
        RECT 332.570 125.960 332.865 127.390 ;
        RECT 123.460 116.150 134.640 117.000 ;
        RECT 132.860 116.070 134.640 116.150 ;
        RECT 120.850 114.790 123.010 115.140 ;
        RECT 148.320 111.000 149.620 111.130 ;
        RECT 132.710 110.955 149.620 111.000 ;
        RECT 116.900 110.410 149.620 110.955 ;
        RECT 116.900 110.270 136.400 110.410 ;
        RECT 117.180 110.170 136.400 110.270 ;
        RECT 117.180 110.105 130.100 110.170 ;
        RECT 117.180 110.100 127.325 110.105 ;
        RECT 117.180 110.095 121.855 110.100 ;
        RECT 131.740 108.600 132.130 110.170 ;
        RECT 148.320 109.920 149.620 110.410 ;
        RECT 111.530 103.010 112.395 104.520 ;
        RECT 148.530 102.860 149.605 104.455 ;
        RECT 234.280 104.290 236.440 104.640 ;
        RECT 234.280 102.700 236.440 103.050 ;
        RECT 234.280 101.110 236.440 101.460 ;
        RECT 260.260 99.530 262.420 99.880 ;
        RECT 281.670 97.940 283.830 98.290 ;
        RECT 234.280 94.750 236.440 95.100 ;
        RECT 213.840 85.510 216.410 87.680 ;
        RECT 220.980 86.935 221.560 87.105 ;
        RECT 233.790 86.995 234.370 87.165 ;
        RECT 238.280 85.900 240.850 88.070 ;
        RECT 220.540 82.900 220.710 85.500 ;
        RECT 221.830 82.900 222.000 85.500 ;
        RECT 233.350 82.960 233.520 85.560 ;
        RECT 234.640 82.960 234.810 85.560 ;
        RECT 264.840 84.840 267.410 87.010 ;
        RECT 277.030 84.995 277.610 85.165 ;
        RECT 284.970 85.055 285.550 85.225 ;
        RECT 292.020 84.550 294.590 86.720 ;
        RECT 276.590 80.960 276.760 83.560 ;
        RECT 277.880 80.960 278.050 83.560 ;
        RECT 284.530 81.020 284.700 83.620 ;
        RECT 285.820 81.020 285.990 83.620 ;
        RECT 121.190 77.780 122.190 78.750 ;
        RECT 32.140 76.110 33.230 76.130 ;
        RECT 34.220 76.110 41.030 76.120 ;
        RECT 32.140 76.060 41.290 76.110 ;
        RECT 32.140 75.980 51.230 76.060 ;
        RECT 32.140 75.130 51.280 75.980 ;
        RECT 27.710 71.650 28.370 72.820 ;
        RECT 32.140 71.650 33.230 75.130 ;
        RECT 34.220 75.080 51.280 75.130 ;
        RECT 34.220 75.060 41.030 75.080 ;
        RECT 48.940 74.990 51.280 75.080 ;
        RECT 48.940 74.500 64.830 74.990 ;
        RECT 49.390 72.290 64.830 74.500 ;
        RECT 76.550 73.900 78.270 74.510 ;
        RECT 85.050 74.000 87.000 75.190 ;
        RECT 111.305 75.180 112.220 76.705 ;
        RECT 148.385 76.580 149.255 76.670 ;
        RECT 148.320 74.990 149.330 76.580 ;
        RECT 80.320 73.900 87.000 74.000 ;
        RECT 70.480 73.850 87.000 73.900 ;
        RECT 49.860 72.250 51.280 72.290 ;
        RECT 27.290 70.170 33.230 71.650 ;
        RECT 45.710 70.730 47.430 70.900 ;
        RECT 27.630 69.500 29.350 69.670 ;
        RECT 27.660 66.970 29.380 67.140 ;
        RECT 27.650 64.380 29.370 64.550 ;
        RECT 27.650 61.830 29.370 62.000 ;
        RECT 27.650 59.280 29.370 59.450 ;
        RECT 27.650 56.730 29.370 56.900 ;
        RECT 27.650 54.180 29.370 54.350 ;
        RECT 27.650 51.630 29.370 51.800 ;
        RECT 27.650 49.080 29.370 49.250 ;
        RECT 31.680 47.200 33.230 70.170 ;
        RECT 49.880 70.560 51.280 72.250 ;
        RECT 45.900 69.710 47.620 69.880 ;
        RECT 45.750 67.670 47.470 67.840 ;
        RECT 45.940 66.650 47.660 66.820 ;
        RECT 45.730 64.780 47.450 64.950 ;
        RECT 45.920 63.760 47.640 63.930 ;
        RECT 45.770 61.910 47.490 62.080 ;
        RECT 45.960 60.890 47.680 61.060 ;
        RECT 45.770 59.020 47.490 59.190 ;
        RECT 45.960 58.000 47.680 58.170 ;
        RECT 45.770 56.130 47.490 56.300 ;
        RECT 45.960 55.110 47.680 55.280 ;
        RECT 45.790 53.220 47.510 53.390 ;
        RECT 45.980 52.200 47.700 52.370 ;
        RECT 45.770 50.340 47.490 50.510 ;
        RECT 45.960 49.320 47.680 49.490 ;
        RECT 45.750 47.490 47.470 47.660 ;
        RECT 49.880 47.330 51.240 70.560 ;
        RECT 60.840 48.710 64.830 72.290 ;
        RECT 70.460 73.400 87.000 73.850 ;
        RECT 70.460 73.350 81.400 73.400 ;
        RECT 70.460 72.900 71.000 73.350 ;
        RECT 80.600 73.340 81.390 73.350 ;
        RECT 70.460 70.230 71.020 72.900 ;
        RECT 80.790 71.440 81.010 73.340 ;
        RECT 85.050 73.030 87.000 73.400 ;
        RECT 85.050 72.880 86.920 73.030 ;
        RECT 81.230 71.440 81.400 71.450 ;
        RECT 80.790 70.560 81.450 71.440 ;
        RECT 81.230 70.510 81.400 70.560 ;
        RECT 192.180 57.750 195.500 62.350 ;
        RECT 186.670 57.700 197.590 57.750 ;
        RECT 186.650 57.200 197.590 57.700 ;
        RECT 186.650 56.750 187.190 57.200 ;
        RECT 186.650 54.080 187.210 56.750 ;
        RECT 192.180 55.880 195.500 57.200 ;
        RECT 196.790 57.190 197.580 57.200 ;
        RECT 196.980 55.290 197.200 57.190 ;
        RECT 197.420 55.290 197.590 55.300 ;
        RECT 196.980 54.410 197.640 55.290 ;
        RECT 197.420 54.360 197.590 54.410 ;
        RECT 147.515 49.155 148.685 49.990 ;
        RECT 76.940 48.710 78.660 48.760 ;
        RECT 60.560 48.150 79.200 48.710 ;
        RECT 147.515 48.655 148.840 49.155 ;
        RECT 84.770 48.330 86.630 48.370 ;
        RECT 84.690 48.270 86.640 48.330 ;
        RECT 81.030 48.150 86.660 48.270 ;
        RECT 147.515 48.255 148.685 48.655 ;
        RECT 60.560 47.600 86.660 48.150 ;
        RECT 27.530 45.790 33.230 47.200 ;
        RECT 45.940 46.470 47.660 46.640 ;
        RECT 32.800 45.690 33.230 45.790 ;
        RECT 49.860 45.400 51.250 47.330 ;
        RECT 60.560 46.870 79.200 47.600 ;
        RECT 80.990 47.590 86.660 47.600 ;
        RECT 81.030 47.540 86.660 47.590 ;
        RECT 46.610 44.330 46.800 44.350 ;
        RECT 46.610 44.300 48.670 44.330 ;
        RECT 49.850 44.300 51.250 45.400 ;
        RECT 70.850 44.480 71.410 46.870 ;
        RECT 81.180 45.690 81.400 47.540 ;
        RECT 84.690 46.170 86.640 47.540 ;
        RECT 84.760 46.130 86.630 46.170 ;
        RECT 111.105 45.705 112.025 47.285 ;
        RECT 81.620 45.690 81.790 45.700 ;
        RECT 81.180 44.810 81.840 45.690 ;
        RECT 81.620 44.760 81.790 44.810 ;
        RECT 46.610 44.100 51.250 44.300 ;
        RECT 127.100 44.100 128.280 44.930 ;
        RECT 46.610 43.140 51.260 44.100 ;
        RECT 46.610 42.950 51.270 43.140 ;
        RECT 46.630 42.910 51.270 42.950 ;
        RECT 46.630 42.850 51.260 42.910 ;
        RECT 48.630 42.840 51.260 42.850 ;
        RECT 48.630 42.810 51.250 42.840 ;
        RECT 250.560 40.160 252.720 40.510 ;
        RECT 250.850 35.220 253.010 35.570 ;
        RECT 246.630 31.720 248.470 31.730 ;
        RECT 246.630 31.650 297.740 31.720 ;
        RECT 246.630 30.100 297.950 31.650 ;
        RECT 246.630 26.540 248.470 30.100 ;
        RECT 284.320 27.720 284.490 28.370 ;
        RECT 284.320 27.240 284.540 27.720 ;
        RECT 284.320 26.610 284.490 27.240 ;
        RECT 243.010 25.330 248.470 26.540 ;
        RECT 270.440 25.430 270.610 25.510 ;
        RECT 243.010 24.740 244.430 25.330 ;
        RECT 242.670 22.670 244.760 24.740 ;
        RECT 246.630 23.770 248.470 25.330 ;
        RECT 270.430 25.070 270.620 25.430 ;
        RECT 249.580 24.760 249.750 24.860 ;
        RECT 249.570 24.580 249.760 24.760 ;
        RECT 270.420 24.590 270.630 25.070 ;
        RECT 275.360 24.860 275.530 25.500 ;
        RECT 283.850 25.100 284.020 25.140 ;
        RECT 249.580 23.820 249.750 24.580 ;
        RECT 270.430 23.890 270.620 24.590 ;
        RECT 275.350 24.380 275.560 24.860 ;
        RECT 283.830 24.620 284.040 25.100 ;
        RECT 283.850 24.560 284.020 24.620 ;
        RECT 270.440 23.810 270.610 23.890 ;
        RECT 275.360 23.800 275.530 24.380 ;
        RECT 295.910 23.710 297.950 30.100 ;
        RECT 118.930 17.500 120.650 19.620 ;
        RECT 112.860 17.450 123.780 17.500 ;
        RECT 112.840 17.380 123.780 17.450 ;
        RECT 135.840 17.410 137.560 18.020 ;
        RECT 154.310 17.500 156.030 18.110 ;
        RECT 148.240 17.490 159.160 17.500 ;
        RECT 140.170 17.410 159.160 17.490 ;
        RECT 129.770 17.380 159.160 17.410 ;
        RECT 112.840 16.950 159.160 17.380 ;
        RECT 112.840 16.500 113.380 16.950 ;
        RECT 122.070 16.910 150.210 16.950 ;
        RECT 158.360 16.940 159.150 16.950 ;
        RECT 122.070 16.880 140.690 16.910 ;
        RECT 112.840 13.830 113.400 16.500 ;
        RECT 123.170 15.040 123.390 16.880 ;
        RECT 129.750 16.860 140.690 16.880 ;
        RECT 129.750 16.410 130.290 16.860 ;
        RECT 139.890 16.850 140.680 16.860 ;
        RECT 123.610 15.040 123.780 15.050 ;
        RECT 123.170 14.160 123.830 15.040 ;
        RECT 123.610 14.110 123.780 14.160 ;
        RECT 129.750 13.740 130.310 16.410 ;
        RECT 140.080 14.950 140.300 16.850 ;
        RECT 148.220 16.500 148.760 16.910 ;
        RECT 140.520 14.950 140.690 14.960 ;
        RECT 140.080 14.070 140.740 14.950 ;
        RECT 140.520 14.020 140.690 14.070 ;
        RECT 148.220 13.830 148.780 16.500 ;
        RECT 158.550 15.040 158.770 16.940 ;
        RECT 158.990 15.040 159.160 15.050 ;
        RECT 158.550 14.160 159.210 15.040 ;
        RECT 158.990 14.110 159.160 14.160 ;
        RECT 693.690 6.880 720.800 7.050 ;
        RECT 693.690 0.740 693.860 6.880 ;
        RECT 695.550 1.255 695.720 6.510 ;
        RECT 698.130 1.255 698.300 6.510 ;
        RECT 700.710 1.255 700.880 6.510 ;
        RECT 703.290 1.255 703.460 6.510 ;
        RECT 705.870 1.255 706.040 6.510 ;
        RECT 708.450 1.255 708.620 6.510 ;
        RECT 711.030 1.255 711.200 6.510 ;
        RECT 713.610 1.255 713.780 6.510 ;
        RECT 716.190 1.255 716.360 6.510 ;
        RECT 718.770 1.255 718.940 6.510 ;
        RECT 694.260 1.085 720.230 1.255 ;
        RECT 720.630 0.740 720.800 6.880 ;
        RECT 693.690 0.570 720.800 0.740 ;
      LAYER mcon ;
        RECT 40.380 323.190 43.810 326.180 ;
        RECT 46.540 323.780 46.710 330.660 ;
        RECT 54.830 323.780 55.000 330.660 ;
        RECT 63.120 323.780 63.290 330.660 ;
        RECT 66.380 323.190 69.810 326.180 ;
        RECT 72.540 323.780 72.710 330.660 ;
        RECT 80.830 323.780 81.000 330.660 ;
        RECT 89.120 323.780 89.290 330.660 ;
        RECT 40.380 313.190 43.810 316.180 ;
        RECT 46.540 315.600 46.710 322.480 ;
        RECT 54.830 315.600 55.000 322.480 ;
        RECT 63.120 315.600 63.290 322.480 ;
        RECT 92.380 323.190 95.810 326.180 ;
        RECT 98.540 323.780 98.710 330.660 ;
        RECT 106.830 323.780 107.000 330.660 ;
        RECT 115.120 323.780 115.290 330.660 ;
        RECT 46.540 307.420 46.710 314.300 ;
        RECT 54.830 307.420 55.000 314.300 ;
        RECT 63.120 307.420 63.290 314.300 ;
        RECT 66.380 313.190 69.810 316.180 ;
        RECT 72.540 315.600 72.710 322.480 ;
        RECT 80.830 315.600 81.000 322.480 ;
        RECT 89.120 315.600 89.290 322.480 ;
        RECT 118.380 323.190 121.810 326.180 ;
        RECT 124.540 323.780 124.710 330.660 ;
        RECT 132.830 323.780 133.000 330.660 ;
        RECT 141.120 323.780 141.290 330.660 ;
        RECT 72.540 307.420 72.710 314.300 ;
        RECT 80.830 307.420 81.000 314.300 ;
        RECT 89.120 307.420 89.290 314.300 ;
        RECT 92.380 313.190 95.810 316.180 ;
        RECT 98.540 315.600 98.710 322.480 ;
        RECT 106.830 315.600 107.000 322.480 ;
        RECT 115.120 315.600 115.290 322.480 ;
        RECT 144.380 323.190 147.810 326.180 ;
        RECT 150.540 323.780 150.710 330.660 ;
        RECT 158.830 323.780 159.000 330.660 ;
        RECT 167.120 323.780 167.290 330.660 ;
        RECT 98.540 307.420 98.710 314.300 ;
        RECT 106.830 307.420 107.000 314.300 ;
        RECT 115.120 307.420 115.290 314.300 ;
        RECT 118.380 313.190 121.810 316.180 ;
        RECT 124.540 315.600 124.710 322.480 ;
        RECT 132.830 315.600 133.000 322.480 ;
        RECT 141.120 315.600 141.290 322.480 ;
        RECT 170.380 323.190 173.810 326.180 ;
        RECT 176.540 323.780 176.710 330.660 ;
        RECT 184.830 323.780 185.000 330.660 ;
        RECT 193.120 323.780 193.290 330.660 ;
        RECT 124.540 307.420 124.710 314.300 ;
        RECT 132.830 307.420 133.000 314.300 ;
        RECT 141.120 307.420 141.290 314.300 ;
        RECT 144.380 313.190 147.810 316.180 ;
        RECT 150.540 315.600 150.710 322.480 ;
        RECT 158.830 315.600 159.000 322.480 ;
        RECT 167.120 315.600 167.290 322.480 ;
        RECT 196.380 323.190 199.810 326.180 ;
        RECT 202.540 323.780 202.710 330.660 ;
        RECT 210.830 323.780 211.000 330.660 ;
        RECT 219.120 323.780 219.290 330.660 ;
        RECT 150.540 307.420 150.710 314.300 ;
        RECT 158.830 307.420 159.000 314.300 ;
        RECT 167.120 307.420 167.290 314.300 ;
        RECT 170.380 313.190 173.810 316.180 ;
        RECT 176.540 315.600 176.710 322.480 ;
        RECT 184.830 315.600 185.000 322.480 ;
        RECT 193.120 315.600 193.290 322.480 ;
        RECT 222.380 323.190 225.810 326.180 ;
        RECT 228.540 323.780 228.710 330.660 ;
        RECT 236.830 323.780 237.000 330.660 ;
        RECT 245.120 323.780 245.290 330.660 ;
        RECT 176.540 307.420 176.710 314.300 ;
        RECT 184.830 307.420 185.000 314.300 ;
        RECT 193.120 307.420 193.290 314.300 ;
        RECT 196.380 313.190 199.810 316.180 ;
        RECT 202.540 315.600 202.710 322.480 ;
        RECT 210.830 315.600 211.000 322.480 ;
        RECT 219.120 315.600 219.290 322.480 ;
        RECT 248.380 323.190 251.810 326.180 ;
        RECT 254.540 323.780 254.710 330.660 ;
        RECT 262.830 323.780 263.000 330.660 ;
        RECT 271.120 323.780 271.290 330.660 ;
        RECT 202.540 307.420 202.710 314.300 ;
        RECT 210.830 307.420 211.000 314.300 ;
        RECT 219.120 307.420 219.290 314.300 ;
        RECT 222.380 313.190 225.810 316.180 ;
        RECT 228.540 315.600 228.710 322.480 ;
        RECT 236.830 315.600 237.000 322.480 ;
        RECT 245.120 315.600 245.290 322.480 ;
        RECT 274.380 323.190 277.810 326.180 ;
        RECT 280.540 323.780 280.710 330.660 ;
        RECT 288.830 323.780 289.000 330.660 ;
        RECT 297.120 323.780 297.290 330.660 ;
        RECT 228.540 307.420 228.710 314.300 ;
        RECT 236.830 307.420 237.000 314.300 ;
        RECT 245.120 307.420 245.290 314.300 ;
        RECT 248.380 313.190 251.810 316.180 ;
        RECT 254.540 315.600 254.710 322.480 ;
        RECT 262.830 315.600 263.000 322.480 ;
        RECT 271.120 315.600 271.290 322.480 ;
        RECT 300.380 323.190 303.810 326.180 ;
        RECT 254.540 307.420 254.710 314.300 ;
        RECT 262.830 307.420 263.000 314.300 ;
        RECT 271.120 307.420 271.290 314.300 ;
        RECT 274.380 313.190 277.810 316.180 ;
        RECT 280.540 315.600 280.710 322.480 ;
        RECT 288.830 315.600 289.000 322.480 ;
        RECT 297.120 315.600 297.290 322.480 ;
        RECT 280.540 307.420 280.710 314.300 ;
        RECT 288.830 307.420 289.000 314.300 ;
        RECT 297.120 307.420 297.290 314.300 ;
        RECT 300.380 313.190 303.810 316.180 ;
        RECT 40.380 303.190 43.810 306.180 ;
        RECT 46.540 299.240 46.710 306.120 ;
        RECT 54.830 299.240 55.000 306.120 ;
        RECT 63.120 299.240 63.290 306.120 ;
        RECT 66.380 303.190 69.810 306.180 ;
        RECT 72.540 299.240 72.710 306.120 ;
        RECT 80.830 299.240 81.000 306.120 ;
        RECT 89.120 299.240 89.290 306.120 ;
        RECT 92.380 303.190 95.810 306.180 ;
        RECT 98.540 299.240 98.710 306.120 ;
        RECT 106.830 299.240 107.000 306.120 ;
        RECT 115.120 299.240 115.290 306.120 ;
        RECT 118.380 303.190 121.810 306.180 ;
        RECT 124.540 299.240 124.710 306.120 ;
        RECT 132.830 299.240 133.000 306.120 ;
        RECT 141.120 299.240 141.290 306.120 ;
        RECT 144.380 303.190 147.810 306.180 ;
        RECT 150.540 299.240 150.710 306.120 ;
        RECT 158.830 299.240 159.000 306.120 ;
        RECT 167.120 299.240 167.290 306.120 ;
        RECT 170.380 303.190 173.810 306.180 ;
        RECT 176.540 299.240 176.710 306.120 ;
        RECT 184.830 299.240 185.000 306.120 ;
        RECT 193.120 299.240 193.290 306.120 ;
        RECT 196.380 303.190 199.810 306.180 ;
        RECT 202.540 299.240 202.710 306.120 ;
        RECT 210.830 299.240 211.000 306.120 ;
        RECT 219.120 299.240 219.290 306.120 ;
        RECT 222.380 303.190 225.810 306.180 ;
        RECT 228.540 299.240 228.710 306.120 ;
        RECT 236.830 299.240 237.000 306.120 ;
        RECT 245.120 299.240 245.290 306.120 ;
        RECT 248.380 303.190 251.810 306.180 ;
        RECT 254.540 299.240 254.710 306.120 ;
        RECT 262.830 299.240 263.000 306.120 ;
        RECT 271.120 299.240 271.290 306.120 ;
        RECT 274.380 303.190 277.810 306.180 ;
        RECT 280.540 299.240 280.710 306.120 ;
        RECT 288.830 299.240 289.000 306.120 ;
        RECT 297.120 299.240 297.290 306.120 ;
        RECT 300.380 303.190 303.810 306.180 ;
        RECT 40.380 293.190 43.810 296.180 ;
        RECT 46.540 291.060 46.710 297.940 ;
        RECT 54.830 291.060 55.000 297.940 ;
        RECT 63.120 291.060 63.290 297.940 ;
        RECT 66.380 293.190 69.810 296.180 ;
        RECT 72.540 291.060 72.710 297.940 ;
        RECT 80.830 291.060 81.000 297.940 ;
        RECT 89.120 291.060 89.290 297.940 ;
        RECT 92.380 293.190 95.810 296.180 ;
        RECT 98.540 291.060 98.710 297.940 ;
        RECT 106.830 291.060 107.000 297.940 ;
        RECT 115.120 291.060 115.290 297.940 ;
        RECT 118.380 293.190 121.810 296.180 ;
        RECT 124.540 291.060 124.710 297.940 ;
        RECT 132.830 291.060 133.000 297.940 ;
        RECT 141.120 291.060 141.290 297.940 ;
        RECT 144.380 293.190 147.810 296.180 ;
        RECT 150.540 291.060 150.710 297.940 ;
        RECT 158.830 291.060 159.000 297.940 ;
        RECT 167.120 291.060 167.290 297.940 ;
        RECT 170.380 293.190 173.810 296.180 ;
        RECT 176.540 291.060 176.710 297.940 ;
        RECT 184.830 291.060 185.000 297.940 ;
        RECT 193.120 291.060 193.290 297.940 ;
        RECT 196.380 293.190 199.810 296.180 ;
        RECT 202.540 291.060 202.710 297.940 ;
        RECT 210.830 291.060 211.000 297.940 ;
        RECT 219.120 291.060 219.290 297.940 ;
        RECT 222.380 293.190 225.810 296.180 ;
        RECT 228.540 291.060 228.710 297.940 ;
        RECT 236.830 291.060 237.000 297.940 ;
        RECT 245.120 291.060 245.290 297.940 ;
        RECT 248.380 293.190 251.810 296.180 ;
        RECT 254.540 291.060 254.710 297.940 ;
        RECT 262.830 291.060 263.000 297.940 ;
        RECT 271.120 291.060 271.290 297.940 ;
        RECT 274.380 293.190 277.810 296.180 ;
        RECT 280.540 291.060 280.710 297.940 ;
        RECT 288.830 291.060 289.000 297.940 ;
        RECT 297.120 291.060 297.290 297.940 ;
        RECT 300.380 293.190 303.810 296.180 ;
        RECT 40.380 283.190 43.810 286.180 ;
        RECT 46.540 282.880 46.710 289.760 ;
        RECT 54.830 282.880 55.000 289.760 ;
        RECT 63.120 282.880 63.290 289.760 ;
        RECT 66.380 283.190 69.810 286.180 ;
        RECT 72.540 282.880 72.710 289.760 ;
        RECT 80.830 282.880 81.000 289.760 ;
        RECT 89.120 282.880 89.290 289.760 ;
        RECT 92.380 283.190 95.810 286.180 ;
        RECT 98.540 282.880 98.710 289.760 ;
        RECT 106.830 282.880 107.000 289.760 ;
        RECT 115.120 282.880 115.290 289.760 ;
        RECT 118.380 283.190 121.810 286.180 ;
        RECT 124.540 282.880 124.710 289.760 ;
        RECT 132.830 282.880 133.000 289.760 ;
        RECT 141.120 282.880 141.290 289.760 ;
        RECT 144.380 283.190 147.810 286.180 ;
        RECT 150.540 282.880 150.710 289.760 ;
        RECT 158.830 282.880 159.000 289.760 ;
        RECT 167.120 282.880 167.290 289.760 ;
        RECT 170.380 283.190 173.810 286.180 ;
        RECT 176.540 282.880 176.710 289.760 ;
        RECT 184.830 282.880 185.000 289.760 ;
        RECT 193.120 282.880 193.290 289.760 ;
        RECT 196.380 283.190 199.810 286.180 ;
        RECT 202.540 282.880 202.710 289.760 ;
        RECT 210.830 282.880 211.000 289.760 ;
        RECT 219.120 282.880 219.290 289.760 ;
        RECT 222.380 283.190 225.810 286.180 ;
        RECT 228.540 282.880 228.710 289.760 ;
        RECT 236.830 282.880 237.000 289.760 ;
        RECT 245.120 282.880 245.290 289.760 ;
        RECT 248.380 283.190 251.810 286.180 ;
        RECT 254.540 282.880 254.710 289.760 ;
        RECT 262.830 282.880 263.000 289.760 ;
        RECT 271.120 282.880 271.290 289.760 ;
        RECT 274.380 283.190 277.810 286.180 ;
        RECT 280.540 282.880 280.710 289.760 ;
        RECT 288.830 282.880 289.000 289.760 ;
        RECT 297.120 282.880 297.290 289.760 ;
        RECT 300.380 283.190 303.810 286.180 ;
        RECT 40.380 273.190 43.810 276.180 ;
        RECT 46.540 274.700 46.710 281.580 ;
        RECT 54.830 274.700 55.000 281.580 ;
        RECT 63.120 274.700 63.290 281.580 ;
        RECT 46.540 266.520 46.710 273.400 ;
        RECT 54.830 266.520 55.000 273.400 ;
        RECT 63.120 266.520 63.290 273.400 ;
        RECT 66.380 273.190 69.810 276.180 ;
        RECT 72.540 274.700 72.710 281.580 ;
        RECT 80.830 274.700 81.000 281.580 ;
        RECT 89.120 274.700 89.290 281.580 ;
        RECT 40.380 263.190 43.810 266.180 ;
        RECT 72.540 266.520 72.710 273.400 ;
        RECT 80.830 266.520 81.000 273.400 ;
        RECT 89.120 266.520 89.290 273.400 ;
        RECT 92.380 273.190 95.810 276.180 ;
        RECT 98.540 274.700 98.710 281.580 ;
        RECT 106.830 274.700 107.000 281.580 ;
        RECT 115.120 274.700 115.290 281.580 ;
        RECT 46.540 258.340 46.710 265.220 ;
        RECT 54.830 258.340 55.000 265.220 ;
        RECT 63.120 258.340 63.290 265.220 ;
        RECT 66.380 263.190 69.810 266.180 ;
        RECT 98.540 266.520 98.710 273.400 ;
        RECT 106.830 266.520 107.000 273.400 ;
        RECT 115.120 266.520 115.290 273.400 ;
        RECT 118.380 273.190 121.810 276.180 ;
        RECT 124.540 274.700 124.710 281.580 ;
        RECT 132.830 274.700 133.000 281.580 ;
        RECT 141.120 274.700 141.290 281.580 ;
        RECT 72.540 258.340 72.710 265.220 ;
        RECT 80.830 258.340 81.000 265.220 ;
        RECT 89.120 258.340 89.290 265.220 ;
        RECT 92.380 263.190 95.810 266.180 ;
        RECT 124.540 266.520 124.710 273.400 ;
        RECT 132.830 266.520 133.000 273.400 ;
        RECT 141.120 266.520 141.290 273.400 ;
        RECT 144.380 273.190 147.810 276.180 ;
        RECT 150.540 274.700 150.710 281.580 ;
        RECT 158.830 274.700 159.000 281.580 ;
        RECT 167.120 274.700 167.290 281.580 ;
        RECT 98.540 258.340 98.710 265.220 ;
        RECT 106.830 258.340 107.000 265.220 ;
        RECT 115.120 258.340 115.290 265.220 ;
        RECT 118.380 263.190 121.810 266.180 ;
        RECT 150.540 266.520 150.710 273.400 ;
        RECT 158.830 266.520 159.000 273.400 ;
        RECT 167.120 266.520 167.290 273.400 ;
        RECT 170.380 273.190 173.810 276.180 ;
        RECT 176.540 274.700 176.710 281.580 ;
        RECT 184.830 274.700 185.000 281.580 ;
        RECT 193.120 274.700 193.290 281.580 ;
        RECT 124.540 258.340 124.710 265.220 ;
        RECT 132.830 258.340 133.000 265.220 ;
        RECT 141.120 258.340 141.290 265.220 ;
        RECT 144.380 263.190 147.810 266.180 ;
        RECT 176.540 266.520 176.710 273.400 ;
        RECT 184.830 266.520 185.000 273.400 ;
        RECT 193.120 266.520 193.290 273.400 ;
        RECT 196.380 273.190 199.810 276.180 ;
        RECT 202.540 274.700 202.710 281.580 ;
        RECT 210.830 274.700 211.000 281.580 ;
        RECT 219.120 274.700 219.290 281.580 ;
        RECT 150.540 258.340 150.710 265.220 ;
        RECT 158.830 258.340 159.000 265.220 ;
        RECT 167.120 258.340 167.290 265.220 ;
        RECT 170.380 263.190 173.810 266.180 ;
        RECT 202.540 266.520 202.710 273.400 ;
        RECT 210.830 266.520 211.000 273.400 ;
        RECT 219.120 266.520 219.290 273.400 ;
        RECT 222.380 273.190 225.810 276.180 ;
        RECT 228.540 274.700 228.710 281.580 ;
        RECT 236.830 274.700 237.000 281.580 ;
        RECT 245.120 274.700 245.290 281.580 ;
        RECT 176.540 258.340 176.710 265.220 ;
        RECT 184.830 258.340 185.000 265.220 ;
        RECT 193.120 258.340 193.290 265.220 ;
        RECT 196.380 263.190 199.810 266.180 ;
        RECT 228.540 266.520 228.710 273.400 ;
        RECT 236.830 266.520 237.000 273.400 ;
        RECT 245.120 266.520 245.290 273.400 ;
        RECT 248.380 273.190 251.810 276.180 ;
        RECT 254.540 274.700 254.710 281.580 ;
        RECT 262.830 274.700 263.000 281.580 ;
        RECT 271.120 274.700 271.290 281.580 ;
        RECT 202.540 258.340 202.710 265.220 ;
        RECT 210.830 258.340 211.000 265.220 ;
        RECT 219.120 258.340 219.290 265.220 ;
        RECT 222.380 263.190 225.810 266.180 ;
        RECT 254.540 266.520 254.710 273.400 ;
        RECT 262.830 266.520 263.000 273.400 ;
        RECT 271.120 266.520 271.290 273.400 ;
        RECT 274.380 273.190 277.810 276.180 ;
        RECT 280.540 274.700 280.710 281.580 ;
        RECT 288.830 274.700 289.000 281.580 ;
        RECT 297.120 274.700 297.290 281.580 ;
        RECT 228.540 258.340 228.710 265.220 ;
        RECT 236.830 258.340 237.000 265.220 ;
        RECT 245.120 258.340 245.290 265.220 ;
        RECT 248.380 263.190 251.810 266.180 ;
        RECT 280.540 266.520 280.710 273.400 ;
        RECT 288.830 266.520 289.000 273.400 ;
        RECT 297.120 266.520 297.290 273.400 ;
        RECT 300.380 273.190 303.810 276.180 ;
        RECT 254.540 258.340 254.710 265.220 ;
        RECT 262.830 258.340 263.000 265.220 ;
        RECT 271.120 258.340 271.290 265.220 ;
        RECT 274.380 263.190 277.810 266.180 ;
        RECT 280.540 258.340 280.710 265.220 ;
        RECT 288.830 258.340 289.000 265.220 ;
        RECT 297.120 258.340 297.290 265.220 ;
        RECT 300.380 263.190 303.810 266.180 ;
        RECT 40.380 253.190 43.810 256.180 ;
        RECT 46.540 250.160 46.710 257.040 ;
        RECT 54.830 250.160 55.000 257.040 ;
        RECT 63.120 250.160 63.290 257.040 ;
        RECT 66.380 253.190 69.810 256.180 ;
        RECT 72.540 250.160 72.710 257.040 ;
        RECT 80.830 250.160 81.000 257.040 ;
        RECT 89.120 250.160 89.290 257.040 ;
        RECT 92.380 253.190 95.810 256.180 ;
        RECT 98.540 250.160 98.710 257.040 ;
        RECT 106.830 250.160 107.000 257.040 ;
        RECT 115.120 250.160 115.290 257.040 ;
        RECT 118.380 253.190 121.810 256.180 ;
        RECT 124.540 250.160 124.710 257.040 ;
        RECT 132.830 250.160 133.000 257.040 ;
        RECT 141.120 250.160 141.290 257.040 ;
        RECT 144.380 253.190 147.810 256.180 ;
        RECT 150.540 250.160 150.710 257.040 ;
        RECT 158.830 250.160 159.000 257.040 ;
        RECT 167.120 250.160 167.290 257.040 ;
        RECT 170.380 253.190 173.810 256.180 ;
        RECT 176.540 250.160 176.710 257.040 ;
        RECT 184.830 250.160 185.000 257.040 ;
        RECT 193.120 250.160 193.290 257.040 ;
        RECT 196.380 253.190 199.810 256.180 ;
        RECT 202.540 250.160 202.710 257.040 ;
        RECT 210.830 250.160 211.000 257.040 ;
        RECT 219.120 250.160 219.290 257.040 ;
        RECT 222.380 253.190 225.810 256.180 ;
        RECT 228.540 250.160 228.710 257.040 ;
        RECT 236.830 250.160 237.000 257.040 ;
        RECT 245.120 250.160 245.290 257.040 ;
        RECT 248.380 253.190 251.810 256.180 ;
        RECT 254.540 250.160 254.710 257.040 ;
        RECT 262.830 250.160 263.000 257.040 ;
        RECT 271.120 250.160 271.290 257.040 ;
        RECT 274.380 253.190 277.810 256.180 ;
        RECT 280.540 250.160 280.710 257.040 ;
        RECT 288.830 250.160 289.000 257.040 ;
        RECT 297.120 250.160 297.290 257.040 ;
        RECT 300.380 253.190 303.810 256.180 ;
        RECT 688.570 249.600 715.340 249.770 ;
        RECT 40.380 241.190 43.810 244.180 ;
        RECT 46.540 241.980 46.710 248.860 ;
        RECT 54.830 241.980 55.000 248.860 ;
        RECT 63.120 241.980 63.290 248.860 ;
        RECT 66.380 241.190 69.810 244.180 ;
        RECT 72.540 241.980 72.710 248.860 ;
        RECT 80.830 241.980 81.000 248.860 ;
        RECT 89.120 241.980 89.290 248.860 ;
        RECT 40.380 231.190 43.810 234.180 ;
        RECT 46.540 233.800 46.710 240.680 ;
        RECT 54.830 233.800 55.000 240.680 ;
        RECT 63.120 233.800 63.290 240.680 ;
        RECT 92.380 241.190 95.810 244.180 ;
        RECT 98.540 241.980 98.710 248.860 ;
        RECT 106.830 241.980 107.000 248.860 ;
        RECT 115.120 241.980 115.290 248.860 ;
        RECT 46.540 225.620 46.710 232.500 ;
        RECT 54.830 225.620 55.000 232.500 ;
        RECT 63.120 225.620 63.290 232.500 ;
        RECT 66.380 231.190 69.810 234.180 ;
        RECT 72.540 233.800 72.710 240.680 ;
        RECT 80.830 233.800 81.000 240.680 ;
        RECT 89.120 233.800 89.290 240.680 ;
        RECT 118.380 241.190 121.810 244.180 ;
        RECT 124.540 241.980 124.710 248.860 ;
        RECT 132.830 241.980 133.000 248.860 ;
        RECT 141.120 241.980 141.290 248.860 ;
        RECT 72.540 225.620 72.710 232.500 ;
        RECT 80.830 225.620 81.000 232.500 ;
        RECT 89.120 225.620 89.290 232.500 ;
        RECT 92.380 231.190 95.810 234.180 ;
        RECT 98.540 233.800 98.710 240.680 ;
        RECT 106.830 233.800 107.000 240.680 ;
        RECT 115.120 233.800 115.290 240.680 ;
        RECT 144.380 241.190 147.810 244.180 ;
        RECT 150.540 241.980 150.710 248.860 ;
        RECT 158.830 241.980 159.000 248.860 ;
        RECT 167.120 241.980 167.290 248.860 ;
        RECT 98.540 225.620 98.710 232.500 ;
        RECT 106.830 225.620 107.000 232.500 ;
        RECT 115.120 225.620 115.290 232.500 ;
        RECT 118.380 231.190 121.810 234.180 ;
        RECT 124.540 233.800 124.710 240.680 ;
        RECT 132.830 233.800 133.000 240.680 ;
        RECT 141.120 233.800 141.290 240.680 ;
        RECT 170.380 241.190 173.810 244.180 ;
        RECT 176.540 241.980 176.710 248.860 ;
        RECT 184.830 241.980 185.000 248.860 ;
        RECT 193.120 241.980 193.290 248.860 ;
        RECT 124.540 225.620 124.710 232.500 ;
        RECT 132.830 225.620 133.000 232.500 ;
        RECT 141.120 225.620 141.290 232.500 ;
        RECT 144.380 231.190 147.810 234.180 ;
        RECT 150.540 233.800 150.710 240.680 ;
        RECT 158.830 233.800 159.000 240.680 ;
        RECT 167.120 233.800 167.290 240.680 ;
        RECT 196.380 241.190 199.810 244.180 ;
        RECT 202.540 241.980 202.710 248.860 ;
        RECT 210.830 241.980 211.000 248.860 ;
        RECT 219.120 241.980 219.290 248.860 ;
        RECT 150.540 225.620 150.710 232.500 ;
        RECT 158.830 225.620 159.000 232.500 ;
        RECT 167.120 225.620 167.290 232.500 ;
        RECT 170.380 231.190 173.810 234.180 ;
        RECT 176.540 233.800 176.710 240.680 ;
        RECT 184.830 233.800 185.000 240.680 ;
        RECT 193.120 233.800 193.290 240.680 ;
        RECT 222.380 241.190 225.810 244.180 ;
        RECT 228.540 241.980 228.710 248.860 ;
        RECT 236.830 241.980 237.000 248.860 ;
        RECT 245.120 241.980 245.290 248.860 ;
        RECT 176.540 225.620 176.710 232.500 ;
        RECT 184.830 225.620 185.000 232.500 ;
        RECT 193.120 225.620 193.290 232.500 ;
        RECT 196.380 231.190 199.810 234.180 ;
        RECT 202.540 233.800 202.710 240.680 ;
        RECT 210.830 233.800 211.000 240.680 ;
        RECT 219.120 233.800 219.290 240.680 ;
        RECT 248.380 241.190 251.810 244.180 ;
        RECT 254.540 241.980 254.710 248.860 ;
        RECT 262.830 241.980 263.000 248.860 ;
        RECT 271.120 241.980 271.290 248.860 ;
        RECT 202.540 225.620 202.710 232.500 ;
        RECT 210.830 225.620 211.000 232.500 ;
        RECT 219.120 225.620 219.290 232.500 ;
        RECT 222.380 231.190 225.810 234.180 ;
        RECT 228.540 233.800 228.710 240.680 ;
        RECT 236.830 233.800 237.000 240.680 ;
        RECT 245.120 233.800 245.290 240.680 ;
        RECT 274.380 241.190 277.810 244.180 ;
        RECT 280.540 241.980 280.710 248.860 ;
        RECT 288.830 241.980 289.000 248.860 ;
        RECT 297.120 241.980 297.290 248.860 ;
        RECT 228.540 225.620 228.710 232.500 ;
        RECT 236.830 225.620 237.000 232.500 ;
        RECT 245.120 225.620 245.290 232.500 ;
        RECT 248.380 231.190 251.810 234.180 ;
        RECT 254.540 233.800 254.710 240.680 ;
        RECT 262.830 233.800 263.000 240.680 ;
        RECT 271.120 233.800 271.290 240.680 ;
        RECT 300.380 241.190 303.810 244.180 ;
        RECT 688.400 244.075 688.570 248.985 ;
        RECT 690.260 244.270 690.430 249.150 ;
        RECT 692.840 244.270 693.010 249.150 ;
        RECT 695.420 244.270 695.590 249.150 ;
        RECT 698.000 244.270 698.170 249.150 ;
        RECT 700.580 244.270 700.750 249.150 ;
        RECT 703.160 244.270 703.330 249.150 ;
        RECT 705.740 244.270 705.910 249.150 ;
        RECT 708.320 244.270 708.490 249.150 ;
        RECT 710.900 244.270 711.070 249.150 ;
        RECT 713.480 244.270 713.650 249.150 ;
        RECT 715.340 244.075 715.510 248.985 ;
        RECT 689.490 243.805 689.910 243.975 ;
        RECT 690.780 243.805 691.200 243.975 ;
        RECT 692.070 243.805 692.490 243.975 ;
        RECT 693.360 243.805 693.780 243.975 ;
        RECT 694.650 243.805 695.070 243.975 ;
        RECT 695.940 243.805 696.360 243.975 ;
        RECT 697.230 243.805 697.650 243.975 ;
        RECT 698.520 243.805 698.940 243.975 ;
        RECT 699.810 243.805 700.230 243.975 ;
        RECT 701.100 243.805 701.520 243.975 ;
        RECT 702.390 243.805 702.810 243.975 ;
        RECT 703.680 243.805 704.100 243.975 ;
        RECT 704.970 243.805 705.390 243.975 ;
        RECT 706.260 243.805 706.680 243.975 ;
        RECT 707.550 243.805 707.970 243.975 ;
        RECT 708.840 243.805 709.260 243.975 ;
        RECT 710.130 243.805 710.550 243.975 ;
        RECT 711.420 243.805 711.840 243.975 ;
        RECT 712.710 243.805 713.130 243.975 ;
        RECT 714.000 243.805 714.420 243.975 ;
        RECT 254.540 225.620 254.710 232.500 ;
        RECT 262.830 225.620 263.000 232.500 ;
        RECT 271.120 225.620 271.290 232.500 ;
        RECT 274.380 231.190 277.810 234.180 ;
        RECT 280.540 233.800 280.710 240.680 ;
        RECT 288.830 233.800 289.000 240.680 ;
        RECT 297.120 233.800 297.290 240.680 ;
        RECT 280.540 225.620 280.710 232.500 ;
        RECT 288.830 225.620 289.000 232.500 ;
        RECT 297.120 225.620 297.290 232.500 ;
        RECT 300.380 231.190 303.810 234.180 ;
        RECT 40.380 221.190 43.810 224.180 ;
        RECT 46.540 217.440 46.710 224.320 ;
        RECT 54.830 217.440 55.000 224.320 ;
        RECT 63.120 217.440 63.290 224.320 ;
        RECT 66.380 221.190 69.810 224.180 ;
        RECT 72.540 217.440 72.710 224.320 ;
        RECT 80.830 217.440 81.000 224.320 ;
        RECT 89.120 217.440 89.290 224.320 ;
        RECT 92.380 221.190 95.810 224.180 ;
        RECT 98.540 217.440 98.710 224.320 ;
        RECT 106.830 217.440 107.000 224.320 ;
        RECT 115.120 217.440 115.290 224.320 ;
        RECT 118.380 221.190 121.810 224.180 ;
        RECT 124.540 217.440 124.710 224.320 ;
        RECT 132.830 217.440 133.000 224.320 ;
        RECT 141.120 217.440 141.290 224.320 ;
        RECT 144.380 221.190 147.810 224.180 ;
        RECT 150.540 217.440 150.710 224.320 ;
        RECT 158.830 217.440 159.000 224.320 ;
        RECT 167.120 217.440 167.290 224.320 ;
        RECT 170.380 221.190 173.810 224.180 ;
        RECT 176.540 217.440 176.710 224.320 ;
        RECT 184.830 217.440 185.000 224.320 ;
        RECT 193.120 217.440 193.290 224.320 ;
        RECT 196.380 221.190 199.810 224.180 ;
        RECT 202.540 217.440 202.710 224.320 ;
        RECT 210.830 217.440 211.000 224.320 ;
        RECT 219.120 217.440 219.290 224.320 ;
        RECT 222.380 221.190 225.810 224.180 ;
        RECT 228.540 217.440 228.710 224.320 ;
        RECT 236.830 217.440 237.000 224.320 ;
        RECT 245.120 217.440 245.290 224.320 ;
        RECT 248.380 221.190 251.810 224.180 ;
        RECT 254.540 217.440 254.710 224.320 ;
        RECT 262.830 217.440 263.000 224.320 ;
        RECT 271.120 217.440 271.290 224.320 ;
        RECT 274.380 221.190 277.810 224.180 ;
        RECT 280.540 217.440 280.710 224.320 ;
        RECT 288.830 217.440 289.000 224.320 ;
        RECT 297.120 217.440 297.290 224.320 ;
        RECT 300.380 221.190 303.810 224.180 ;
        RECT 40.380 211.190 43.810 214.180 ;
        RECT 46.540 209.260 46.710 216.140 ;
        RECT 54.830 209.260 55.000 216.140 ;
        RECT 63.120 209.260 63.290 216.140 ;
        RECT 66.380 211.190 69.810 214.180 ;
        RECT 72.540 209.260 72.710 216.140 ;
        RECT 80.830 209.260 81.000 216.140 ;
        RECT 89.120 209.260 89.290 216.140 ;
        RECT 92.380 211.190 95.810 214.180 ;
        RECT 98.540 209.260 98.710 216.140 ;
        RECT 106.830 209.260 107.000 216.140 ;
        RECT 115.120 209.260 115.290 216.140 ;
        RECT 118.380 211.190 121.810 214.180 ;
        RECT 124.540 209.260 124.710 216.140 ;
        RECT 132.830 209.260 133.000 216.140 ;
        RECT 141.120 209.260 141.290 216.140 ;
        RECT 144.380 211.190 147.810 214.180 ;
        RECT 150.540 209.260 150.710 216.140 ;
        RECT 158.830 209.260 159.000 216.140 ;
        RECT 167.120 209.260 167.290 216.140 ;
        RECT 170.380 211.190 173.810 214.180 ;
        RECT 176.540 209.260 176.710 216.140 ;
        RECT 184.830 209.260 185.000 216.140 ;
        RECT 193.120 209.260 193.290 216.140 ;
        RECT 196.380 211.190 199.810 214.180 ;
        RECT 202.540 209.260 202.710 216.140 ;
        RECT 210.830 209.260 211.000 216.140 ;
        RECT 219.120 209.260 219.290 216.140 ;
        RECT 222.380 211.190 225.810 214.180 ;
        RECT 228.540 209.260 228.710 216.140 ;
        RECT 236.830 209.260 237.000 216.140 ;
        RECT 245.120 209.260 245.290 216.140 ;
        RECT 248.380 211.190 251.810 214.180 ;
        RECT 254.540 209.260 254.710 216.140 ;
        RECT 262.830 209.260 263.000 216.140 ;
        RECT 271.120 209.260 271.290 216.140 ;
        RECT 274.380 211.190 277.810 214.180 ;
        RECT 280.540 209.260 280.710 216.140 ;
        RECT 288.830 209.260 289.000 216.140 ;
        RECT 297.120 209.260 297.290 216.140 ;
        RECT 300.380 211.190 303.810 214.180 ;
        RECT 40.380 201.190 43.810 204.180 ;
        RECT 46.540 201.080 46.710 207.960 ;
        RECT 54.830 201.080 55.000 207.960 ;
        RECT 63.120 201.080 63.290 207.960 ;
        RECT 66.380 201.190 69.810 204.180 ;
        RECT 72.540 201.080 72.710 207.960 ;
        RECT 80.830 201.080 81.000 207.960 ;
        RECT 89.120 201.080 89.290 207.960 ;
        RECT 92.380 201.190 95.810 204.180 ;
        RECT 98.540 201.080 98.710 207.960 ;
        RECT 106.830 201.080 107.000 207.960 ;
        RECT 115.120 201.080 115.290 207.960 ;
        RECT 118.380 201.190 121.810 204.180 ;
        RECT 124.540 201.080 124.710 207.960 ;
        RECT 132.830 201.080 133.000 207.960 ;
        RECT 141.120 201.080 141.290 207.960 ;
        RECT 144.380 201.190 147.810 204.180 ;
        RECT 150.540 201.080 150.710 207.960 ;
        RECT 158.830 201.080 159.000 207.960 ;
        RECT 167.120 201.080 167.290 207.960 ;
        RECT 170.380 201.190 173.810 204.180 ;
        RECT 176.540 201.080 176.710 207.960 ;
        RECT 184.830 201.080 185.000 207.960 ;
        RECT 193.120 201.080 193.290 207.960 ;
        RECT 196.380 201.190 199.810 204.180 ;
        RECT 202.540 201.080 202.710 207.960 ;
        RECT 210.830 201.080 211.000 207.960 ;
        RECT 219.120 201.080 219.290 207.960 ;
        RECT 222.380 201.190 225.810 204.180 ;
        RECT 228.540 201.080 228.710 207.960 ;
        RECT 236.830 201.080 237.000 207.960 ;
        RECT 245.120 201.080 245.290 207.960 ;
        RECT 248.380 201.190 251.810 204.180 ;
        RECT 254.540 201.080 254.710 207.960 ;
        RECT 262.830 201.080 263.000 207.960 ;
        RECT 271.120 201.080 271.290 207.960 ;
        RECT 274.380 201.190 277.810 204.180 ;
        RECT 280.540 201.080 280.710 207.960 ;
        RECT 288.830 201.080 289.000 207.960 ;
        RECT 297.120 201.080 297.290 207.960 ;
        RECT 300.380 201.190 303.810 204.180 ;
        RECT 40.380 191.190 43.810 194.180 ;
        RECT 46.540 192.900 46.710 199.780 ;
        RECT 54.830 192.900 55.000 199.780 ;
        RECT 63.120 192.900 63.290 199.780 ;
        RECT 46.540 184.720 46.710 191.600 ;
        RECT 54.830 184.720 55.000 191.600 ;
        RECT 63.120 184.720 63.290 191.600 ;
        RECT 66.380 191.190 69.810 194.180 ;
        RECT 72.540 192.900 72.710 199.780 ;
        RECT 80.830 192.900 81.000 199.780 ;
        RECT 89.120 192.900 89.290 199.780 ;
        RECT 40.380 181.190 43.810 184.180 ;
        RECT 72.540 184.720 72.710 191.600 ;
        RECT 80.830 184.720 81.000 191.600 ;
        RECT 89.120 184.720 89.290 191.600 ;
        RECT 92.380 191.190 95.810 194.180 ;
        RECT 98.540 192.900 98.710 199.780 ;
        RECT 106.830 192.900 107.000 199.780 ;
        RECT 115.120 192.900 115.290 199.780 ;
        RECT 46.540 176.540 46.710 183.420 ;
        RECT 54.830 176.540 55.000 183.420 ;
        RECT 63.120 176.540 63.290 183.420 ;
        RECT 66.380 181.190 69.810 184.180 ;
        RECT 98.540 184.720 98.710 191.600 ;
        RECT 106.830 184.720 107.000 191.600 ;
        RECT 115.120 184.720 115.290 191.600 ;
        RECT 118.380 191.190 121.810 194.180 ;
        RECT 124.540 192.900 124.710 199.780 ;
        RECT 132.830 192.900 133.000 199.780 ;
        RECT 141.120 192.900 141.290 199.780 ;
        RECT 72.540 176.540 72.710 183.420 ;
        RECT 80.830 176.540 81.000 183.420 ;
        RECT 89.120 176.540 89.290 183.420 ;
        RECT 92.380 181.190 95.810 184.180 ;
        RECT 124.540 184.720 124.710 191.600 ;
        RECT 132.830 184.720 133.000 191.600 ;
        RECT 141.120 184.720 141.290 191.600 ;
        RECT 144.380 191.190 147.810 194.180 ;
        RECT 150.540 192.900 150.710 199.780 ;
        RECT 158.830 192.900 159.000 199.780 ;
        RECT 167.120 192.900 167.290 199.780 ;
        RECT 98.540 176.540 98.710 183.420 ;
        RECT 106.830 176.540 107.000 183.420 ;
        RECT 115.120 176.540 115.290 183.420 ;
        RECT 118.380 181.190 121.810 184.180 ;
        RECT 150.540 184.720 150.710 191.600 ;
        RECT 158.830 184.720 159.000 191.600 ;
        RECT 167.120 184.720 167.290 191.600 ;
        RECT 170.380 191.190 173.810 194.180 ;
        RECT 176.540 192.900 176.710 199.780 ;
        RECT 184.830 192.900 185.000 199.780 ;
        RECT 193.120 192.900 193.290 199.780 ;
        RECT 124.540 176.540 124.710 183.420 ;
        RECT 132.830 176.540 133.000 183.420 ;
        RECT 141.120 176.540 141.290 183.420 ;
        RECT 144.380 181.190 147.810 184.180 ;
        RECT 176.540 184.720 176.710 191.600 ;
        RECT 184.830 184.720 185.000 191.600 ;
        RECT 193.120 184.720 193.290 191.600 ;
        RECT 196.380 191.190 199.810 194.180 ;
        RECT 202.540 192.900 202.710 199.780 ;
        RECT 210.830 192.900 211.000 199.780 ;
        RECT 219.120 192.900 219.290 199.780 ;
        RECT 150.540 176.540 150.710 183.420 ;
        RECT 158.830 176.540 159.000 183.420 ;
        RECT 167.120 176.540 167.290 183.420 ;
        RECT 170.380 181.190 173.810 184.180 ;
        RECT 202.540 184.720 202.710 191.600 ;
        RECT 210.830 184.720 211.000 191.600 ;
        RECT 219.120 184.720 219.290 191.600 ;
        RECT 222.380 191.190 225.810 194.180 ;
        RECT 228.540 192.900 228.710 199.780 ;
        RECT 236.830 192.900 237.000 199.780 ;
        RECT 245.120 192.900 245.290 199.780 ;
        RECT 176.540 176.540 176.710 183.420 ;
        RECT 184.830 176.540 185.000 183.420 ;
        RECT 193.120 176.540 193.290 183.420 ;
        RECT 196.380 181.190 199.810 184.180 ;
        RECT 228.540 184.720 228.710 191.600 ;
        RECT 236.830 184.720 237.000 191.600 ;
        RECT 245.120 184.720 245.290 191.600 ;
        RECT 248.380 191.190 251.810 194.180 ;
        RECT 254.540 192.900 254.710 199.780 ;
        RECT 262.830 192.900 263.000 199.780 ;
        RECT 271.120 192.900 271.290 199.780 ;
        RECT 202.540 176.540 202.710 183.420 ;
        RECT 210.830 176.540 211.000 183.420 ;
        RECT 219.120 176.540 219.290 183.420 ;
        RECT 222.380 181.190 225.810 184.180 ;
        RECT 254.540 184.720 254.710 191.600 ;
        RECT 262.830 184.720 263.000 191.600 ;
        RECT 271.120 184.720 271.290 191.600 ;
        RECT 274.380 191.190 277.810 194.180 ;
        RECT 280.540 192.900 280.710 199.780 ;
        RECT 288.830 192.900 289.000 199.780 ;
        RECT 297.120 192.900 297.290 199.780 ;
        RECT 228.540 176.540 228.710 183.420 ;
        RECT 236.830 176.540 237.000 183.420 ;
        RECT 245.120 176.540 245.290 183.420 ;
        RECT 248.380 181.190 251.810 184.180 ;
        RECT 280.540 184.720 280.710 191.600 ;
        RECT 288.830 184.720 289.000 191.600 ;
        RECT 297.120 184.720 297.290 191.600 ;
        RECT 300.380 191.190 303.810 194.180 ;
        RECT 254.540 176.540 254.710 183.420 ;
        RECT 262.830 176.540 263.000 183.420 ;
        RECT 271.120 176.540 271.290 183.420 ;
        RECT 274.380 181.190 277.810 184.180 ;
        RECT 280.540 176.540 280.710 183.420 ;
        RECT 288.830 176.540 289.000 183.420 ;
        RECT 297.120 176.540 297.290 183.420 ;
        RECT 300.380 181.190 303.810 184.180 ;
        RECT 40.380 171.190 43.810 174.180 ;
        RECT 46.540 168.360 46.710 175.240 ;
        RECT 54.830 168.360 55.000 175.240 ;
        RECT 63.120 168.360 63.290 175.240 ;
        RECT 66.380 171.190 69.810 174.180 ;
        RECT 72.540 168.360 72.710 175.240 ;
        RECT 80.830 168.360 81.000 175.240 ;
        RECT 89.120 168.360 89.290 175.240 ;
        RECT 92.380 171.190 95.810 174.180 ;
        RECT 98.540 168.360 98.710 175.240 ;
        RECT 106.830 168.360 107.000 175.240 ;
        RECT 115.120 168.360 115.290 175.240 ;
        RECT 118.380 171.190 121.810 174.180 ;
        RECT 124.540 168.360 124.710 175.240 ;
        RECT 132.830 168.360 133.000 175.240 ;
        RECT 141.120 168.360 141.290 175.240 ;
        RECT 144.380 171.190 147.810 174.180 ;
        RECT 150.540 168.360 150.710 175.240 ;
        RECT 158.830 168.360 159.000 175.240 ;
        RECT 167.120 168.360 167.290 175.240 ;
        RECT 170.380 171.190 173.810 174.180 ;
        RECT 176.540 168.360 176.710 175.240 ;
        RECT 184.830 168.360 185.000 175.240 ;
        RECT 193.120 168.360 193.290 175.240 ;
        RECT 196.380 171.190 199.810 174.180 ;
        RECT 202.540 168.360 202.710 175.240 ;
        RECT 210.830 168.360 211.000 175.240 ;
        RECT 219.120 168.360 219.290 175.240 ;
        RECT 222.380 171.190 225.810 174.180 ;
        RECT 228.540 168.360 228.710 175.240 ;
        RECT 236.830 168.360 237.000 175.240 ;
        RECT 245.120 168.360 245.290 175.240 ;
        RECT 248.380 171.190 251.810 174.180 ;
        RECT 254.540 168.360 254.710 175.240 ;
        RECT 262.830 168.360 263.000 175.240 ;
        RECT 271.120 168.360 271.290 175.240 ;
        RECT 274.380 171.190 277.810 174.180 ;
        RECT 280.540 168.360 280.710 175.240 ;
        RECT 288.830 168.360 289.000 175.240 ;
        RECT 297.120 168.360 297.290 175.240 ;
        RECT 300.380 171.190 303.810 174.180 ;
        RECT 129.120 135.820 129.290 136.600 ;
        RECT 151.020 135.380 151.190 136.160 ;
        RECT 171.810 135.150 171.980 135.930 ;
        RECT 309.345 133.455 309.515 133.625 ;
        RECT 309.825 133.455 309.995 133.625 ;
        RECT 310.305 133.455 310.475 133.625 ;
        RECT 310.785 133.455 310.955 133.625 ;
        RECT 311.265 133.455 311.435 133.625 ;
        RECT 311.745 133.455 311.915 133.625 ;
        RECT 312.225 133.455 312.395 133.625 ;
        RECT 312.705 133.455 312.875 133.625 ;
        RECT 313.185 133.455 313.355 133.625 ;
        RECT 313.665 133.455 313.835 133.625 ;
        RECT 314.145 133.455 314.315 133.625 ;
        RECT 314.625 133.455 314.795 133.625 ;
        RECT 315.105 133.455 315.275 133.625 ;
        RECT 315.585 133.455 315.755 133.625 ;
        RECT 316.065 133.455 316.235 133.625 ;
        RECT 316.545 133.455 316.715 133.625 ;
        RECT 317.025 133.455 317.195 133.625 ;
        RECT 317.505 133.455 317.675 133.625 ;
        RECT 317.985 133.455 318.155 133.625 ;
        RECT 318.465 133.455 318.635 133.625 ;
        RECT 318.945 133.455 319.115 133.625 ;
        RECT 319.425 133.455 319.595 133.625 ;
        RECT 319.905 133.455 320.075 133.625 ;
        RECT 320.385 133.455 320.555 133.625 ;
        RECT 320.865 133.455 321.035 133.625 ;
        RECT 323.035 133.490 323.205 133.660 ;
        RECT 323.515 133.490 323.685 133.660 ;
        RECT 323.995 133.490 324.165 133.660 ;
        RECT 324.475 133.490 324.645 133.660 ;
        RECT 324.955 133.490 325.125 133.660 ;
        RECT 325.435 133.490 325.605 133.660 ;
        RECT 325.915 133.490 326.085 133.660 ;
        RECT 326.395 133.490 326.565 133.660 ;
        RECT 326.875 133.490 327.045 133.660 ;
        RECT 327.355 133.490 327.525 133.660 ;
        RECT 327.835 133.490 328.005 133.660 ;
        RECT 328.315 133.490 328.485 133.660 ;
        RECT 328.795 133.490 328.965 133.660 ;
        RECT 329.275 133.490 329.445 133.660 ;
        RECT 329.755 133.490 329.925 133.660 ;
        RECT 330.235 133.490 330.405 133.660 ;
        RECT 330.715 133.490 330.885 133.660 ;
        RECT 331.195 133.490 331.365 133.660 ;
        RECT 331.675 133.490 331.845 133.660 ;
        RECT 332.155 133.490 332.325 133.660 ;
        RECT 332.635 133.490 332.805 133.660 ;
        RECT 333.115 133.490 333.285 133.660 ;
        RECT 333.595 133.490 333.765 133.660 ;
        RECT 334.075 133.490 334.245 133.660 ;
        RECT 334.555 133.490 334.725 133.660 ;
        RECT 321.145 127.390 321.315 127.560 ;
        RECT 321.625 127.390 321.795 127.560 ;
        RECT 322.105 127.390 322.275 127.560 ;
        RECT 322.585 127.390 322.755 127.560 ;
        RECT 323.065 127.390 323.235 127.560 ;
        RECT 323.545 127.390 323.715 127.560 ;
        RECT 324.025 127.390 324.195 127.560 ;
        RECT 324.505 127.390 324.675 127.560 ;
        RECT 324.985 127.390 325.155 127.560 ;
        RECT 325.465 127.390 325.635 127.560 ;
        RECT 325.945 127.390 326.115 127.560 ;
        RECT 326.425 127.390 326.595 127.560 ;
        RECT 326.905 127.390 327.075 127.560 ;
        RECT 327.385 127.390 327.555 127.560 ;
        RECT 327.865 127.390 328.035 127.560 ;
        RECT 328.345 127.390 328.515 127.560 ;
        RECT 328.825 127.390 328.995 127.560 ;
        RECT 329.305 127.390 329.475 127.560 ;
        RECT 329.785 127.390 329.955 127.560 ;
        RECT 330.265 127.390 330.435 127.560 ;
        RECT 330.745 127.390 330.915 127.560 ;
        RECT 331.225 127.390 331.395 127.560 ;
        RECT 331.705 127.390 331.875 127.560 ;
        RECT 332.185 127.390 332.355 127.560 ;
        RECT 332.665 127.390 332.835 127.560 ;
        RECT 123.755 116.590 125.740 116.780 ;
        RECT 120.935 114.870 122.920 115.060 ;
        RECT 122.940 110.380 124.420 110.800 ;
        RECT 148.640 110.090 149.390 110.910 ;
        RECT 234.370 104.370 236.355 104.560 ;
        RECT 234.370 102.780 236.355 102.970 ;
        RECT 234.370 101.190 236.355 101.380 ;
        RECT 260.350 99.610 262.335 99.800 ;
        RECT 281.755 98.020 283.740 98.210 ;
        RECT 234.370 94.830 236.355 95.020 ;
        RECT 214.310 86.000 215.940 87.200 ;
        RECT 221.060 86.935 221.480 87.105 ;
        RECT 233.870 86.995 234.290 87.165 ;
        RECT 238.750 86.390 240.380 87.590 ;
        RECT 220.540 82.980 220.710 85.420 ;
        RECT 221.830 82.980 222.000 85.420 ;
        RECT 233.350 83.040 233.520 85.480 ;
        RECT 234.640 83.040 234.810 85.480 ;
        RECT 265.310 85.330 266.940 86.530 ;
        RECT 277.110 84.995 277.530 85.165 ;
        RECT 285.050 85.055 285.470 85.225 ;
        RECT 292.490 85.040 294.120 86.240 ;
        RECT 276.590 81.040 276.760 83.480 ;
        RECT 277.880 81.040 278.050 83.480 ;
        RECT 284.530 81.100 284.700 83.540 ;
        RECT 285.820 81.100 285.990 83.540 ;
        RECT 49.610 72.640 51.570 74.640 ;
        RECT 28.070 70.650 28.600 71.370 ;
        RECT 45.790 70.730 47.350 70.900 ;
        RECT 27.710 69.500 29.270 69.670 ;
        RECT 27.740 66.970 29.300 67.140 ;
        RECT 27.730 64.380 29.290 64.550 ;
        RECT 27.730 61.830 29.290 62.000 ;
        RECT 27.730 59.280 29.290 59.450 ;
        RECT 27.730 56.730 29.290 56.900 ;
        RECT 27.730 54.180 29.290 54.350 ;
        RECT 27.730 51.630 29.290 51.800 ;
        RECT 27.730 49.080 29.290 49.250 ;
        RECT 45.980 69.710 47.540 69.880 ;
        RECT 45.830 67.670 47.390 67.840 ;
        RECT 46.020 66.650 47.580 66.820 ;
        RECT 45.810 64.780 47.370 64.950 ;
        RECT 46.000 63.760 47.560 63.930 ;
        RECT 45.850 61.910 47.410 62.080 ;
        RECT 46.040 60.890 47.600 61.060 ;
        RECT 45.850 59.020 47.410 59.190 ;
        RECT 46.040 58.000 47.600 58.170 ;
        RECT 45.850 56.130 47.410 56.300 ;
        RECT 46.040 55.110 47.600 55.280 ;
        RECT 45.870 53.220 47.430 53.390 ;
        RECT 46.060 52.200 47.620 52.370 ;
        RECT 45.850 50.340 47.410 50.510 ;
        RECT 46.040 49.320 47.600 49.490 ;
        RECT 45.830 47.490 47.390 47.660 ;
        RECT 85.460 73.530 86.340 74.420 ;
        RECT 81.230 70.590 81.400 71.370 ;
        RECT 193.150 58.970 194.030 59.860 ;
        RECT 197.420 54.440 197.590 55.220 ;
        RECT 147.585 49.490 148.595 49.920 ;
        RECT 147.580 48.770 148.595 49.490 ;
        RECT 147.585 48.345 148.595 48.770 ;
        RECT 46.020 46.470 47.580 46.640 ;
        RECT 85.170 46.780 86.050 47.670 ;
        RECT 111.200 45.870 111.915 47.190 ;
        RECT 81.620 44.840 81.790 45.620 ;
        RECT 250.650 40.240 252.635 40.430 ;
        RECT 250.940 35.300 252.925 35.490 ;
        RECT 284.320 26.690 284.490 28.290 ;
        RECT 242.950 22.900 244.460 24.580 ;
        RECT 249.580 23.900 249.750 24.780 ;
        RECT 270.430 23.890 270.620 25.430 ;
        RECT 275.360 23.880 275.530 25.420 ;
        RECT 283.850 24.640 284.020 25.060 ;
        RECT 119.420 18.640 120.280 19.270 ;
        RECT 123.610 14.190 123.780 14.970 ;
        RECT 140.520 14.100 140.690 14.880 ;
        RECT 158.990 14.190 159.160 14.970 ;
        RECT 693.860 6.880 720.630 7.050 ;
        RECT 693.690 1.355 693.860 6.265 ;
        RECT 695.550 1.550 695.720 6.430 ;
        RECT 698.130 1.550 698.300 6.430 ;
        RECT 700.710 1.550 700.880 6.430 ;
        RECT 703.290 1.550 703.460 6.430 ;
        RECT 705.870 1.550 706.040 6.430 ;
        RECT 708.450 1.550 708.620 6.430 ;
        RECT 711.030 1.550 711.200 6.430 ;
        RECT 713.610 1.550 713.780 6.430 ;
        RECT 716.190 1.550 716.360 6.430 ;
        RECT 718.770 1.550 718.940 6.430 ;
        RECT 720.630 1.355 720.800 6.265 ;
        RECT 694.780 1.085 695.200 1.255 ;
        RECT 696.070 1.085 696.490 1.255 ;
        RECT 697.360 1.085 697.780 1.255 ;
        RECT 698.650 1.085 699.070 1.255 ;
        RECT 699.940 1.085 700.360 1.255 ;
        RECT 701.230 1.085 701.650 1.255 ;
        RECT 702.520 1.085 702.940 1.255 ;
        RECT 703.810 1.085 704.230 1.255 ;
        RECT 705.100 1.085 705.520 1.255 ;
        RECT 706.390 1.085 706.810 1.255 ;
        RECT 707.680 1.085 708.100 1.255 ;
        RECT 708.970 1.085 709.390 1.255 ;
        RECT 710.260 1.085 710.680 1.255 ;
        RECT 711.550 1.085 711.970 1.255 ;
        RECT 712.840 1.085 713.260 1.255 ;
        RECT 714.130 1.085 714.550 1.255 ;
        RECT 715.420 1.085 715.840 1.255 ;
        RECT 716.710 1.085 717.130 1.255 ;
        RECT 718.000 1.085 718.420 1.255 ;
        RECT 719.290 1.085 719.710 1.255 ;
      LAYER met1 ;
        RECT 46.510 329.550 46.740 330.720 ;
        RECT 43.050 329.530 49.690 329.550 ;
        RECT 54.800 329.530 55.030 330.720 ;
        RECT 63.090 329.530 63.320 330.720 ;
        RECT 72.510 329.530 72.740 330.720 ;
        RECT 80.800 329.530 81.030 330.720 ;
        RECT 89.090 329.530 89.320 330.720 ;
        RECT 98.510 329.590 98.740 330.720 ;
        RECT 92.160 329.530 98.960 329.590 ;
        RECT 106.800 329.530 107.030 330.720 ;
        RECT 115.090 329.530 115.320 330.720 ;
        RECT 124.510 329.530 124.740 330.720 ;
        RECT 132.800 329.530 133.030 330.720 ;
        RECT 141.090 329.530 141.320 330.720 ;
        RECT 150.510 329.530 150.740 330.720 ;
        RECT 158.800 329.530 159.030 330.720 ;
        RECT 167.090 329.530 167.320 330.720 ;
        RECT 176.510 329.530 176.740 330.720 ;
        RECT 184.800 329.530 185.030 330.720 ;
        RECT 193.090 329.530 193.320 330.720 ;
        RECT 202.510 329.530 202.740 330.720 ;
        RECT 210.800 329.530 211.030 330.720 ;
        RECT 219.090 329.530 219.320 330.720 ;
        RECT 228.510 329.570 228.740 330.720 ;
        RECT 222.150 329.530 228.950 329.570 ;
        RECT 236.800 329.530 237.030 330.720 ;
        RECT 245.090 329.530 245.320 330.720 ;
        RECT 254.510 329.530 254.740 330.720 ;
        RECT 262.800 329.530 263.030 330.720 ;
        RECT 271.090 329.530 271.320 330.720 ;
        RECT 280.510 329.530 280.740 330.720 ;
        RECT 288.800 329.530 289.030 330.720 ;
        RECT 297.090 329.530 297.320 330.720 ;
        RECT 43.050 329.450 66.290 329.530 ;
        RECT 72.250 329.450 118.290 329.530 ;
        RECT 43.050 329.390 118.290 329.450 ;
        RECT 124.250 329.520 144.290 329.530 ;
        RECT 150.250 329.520 170.290 329.530 ;
        RECT 124.250 329.460 170.290 329.520 ;
        RECT 176.250 329.460 196.290 329.530 ;
        RECT 202.250 329.460 248.290 329.530 ;
        RECT 124.250 329.390 248.290 329.460 ;
        RECT 43.050 329.360 248.290 329.390 ;
        RECT 254.250 329.460 274.290 329.530 ;
        RECT 280.250 329.460 300.290 329.530 ;
        RECT 254.250 329.360 300.290 329.460 ;
        RECT 43.050 327.320 300.290 329.360 ;
        RECT 39.400 327.300 300.290 327.320 ;
        RECT 39.400 325.800 304.560 327.300 ;
        RECT 39.400 325.700 96.560 325.800 ;
        RECT 98.250 325.780 304.560 325.800 ;
        RECT 98.250 325.730 226.560 325.780 ;
        RECT 98.250 325.700 148.560 325.730 ;
        RECT 150.250 325.700 226.560 325.730 ;
        RECT 228.250 325.700 304.560 325.780 ;
        RECT 39.400 325.630 49.690 325.700 ;
        RECT 39.400 321.310 44.730 325.630 ;
        RECT 46.510 323.720 46.740 325.630 ;
        RECT 54.800 323.720 55.030 325.700 ;
        RECT 63.090 323.720 63.320 325.700 ;
        RECT 64.020 325.650 64.310 325.700 ;
        RECT 65.580 325.660 72.740 325.700 ;
        RECT 46.510 321.310 46.740 322.540 ;
        RECT 39.400 321.280 50.910 321.310 ;
        RECT 54.800 321.280 55.030 322.540 ;
        RECT 63.090 321.280 63.320 322.540 ;
        RECT 65.580 321.280 70.560 325.660 ;
        RECT 72.510 323.720 72.740 325.660 ;
        RECT 80.800 323.720 81.030 325.700 ;
        RECT 89.090 323.720 89.320 325.700 ;
        RECT 90.020 325.650 90.310 325.700 ;
        RECT 72.510 321.280 72.740 322.540 ;
        RECT 80.800 321.280 81.030 322.540 ;
        RECT 89.090 321.280 89.320 322.540 ;
        RECT 91.580 321.280 96.560 325.700 ;
        RECT 98.510 323.720 98.740 325.700 ;
        RECT 106.800 323.720 107.030 325.700 ;
        RECT 115.090 323.720 115.320 325.700 ;
        RECT 116.020 325.650 116.310 325.700 ;
        RECT 117.580 325.600 124.760 325.700 ;
        RECT 98.510 321.280 98.740 322.540 ;
        RECT 106.800 321.280 107.030 322.540 ;
        RECT 115.090 321.280 115.320 322.540 ;
        RECT 117.580 321.280 122.560 325.600 ;
        RECT 124.510 323.720 124.740 325.600 ;
        RECT 132.800 323.720 133.030 325.700 ;
        RECT 141.090 323.720 141.320 325.700 ;
        RECT 142.020 325.650 142.310 325.700 ;
        RECT 124.510 321.280 124.740 322.540 ;
        RECT 132.800 321.280 133.030 322.540 ;
        RECT 141.090 321.280 141.320 322.540 ;
        RECT 143.580 321.280 148.560 325.700 ;
        RECT 150.510 323.720 150.740 325.700 ;
        RECT 158.800 323.720 159.030 325.700 ;
        RECT 167.090 323.720 167.320 325.700 ;
        RECT 168.020 325.650 168.310 325.700 ;
        RECT 169.580 325.670 176.970 325.700 ;
        RECT 150.510 321.280 150.740 322.540 ;
        RECT 158.800 321.280 159.030 322.540 ;
        RECT 167.090 321.280 167.320 322.540 ;
        RECT 169.580 321.280 174.560 325.670 ;
        RECT 176.510 323.720 176.740 325.670 ;
        RECT 184.800 323.720 185.030 325.700 ;
        RECT 193.090 323.720 193.320 325.700 ;
        RECT 194.020 325.650 194.310 325.700 ;
        RECT 195.580 325.670 202.970 325.700 ;
        RECT 176.510 321.280 176.740 322.540 ;
        RECT 184.800 321.280 185.030 322.540 ;
        RECT 193.090 321.280 193.320 322.540 ;
        RECT 195.580 321.280 200.560 325.670 ;
        RECT 202.510 323.720 202.740 325.670 ;
        RECT 210.800 323.720 211.030 325.700 ;
        RECT 219.090 323.720 219.320 325.700 ;
        RECT 220.020 325.650 220.310 325.700 ;
        RECT 202.510 321.280 202.740 322.540 ;
        RECT 210.800 321.280 211.030 322.540 ;
        RECT 219.090 321.280 219.320 322.540 ;
        RECT 221.580 321.280 226.560 325.700 ;
        RECT 228.510 323.720 228.740 325.700 ;
        RECT 236.800 323.720 237.030 325.700 ;
        RECT 245.090 323.720 245.320 325.700 ;
        RECT 246.020 325.650 246.310 325.700 ;
        RECT 247.580 325.570 254.780 325.700 ;
        RECT 228.510 321.280 228.740 322.540 ;
        RECT 236.800 321.280 237.030 322.540 ;
        RECT 245.090 321.280 245.320 322.540 ;
        RECT 247.580 321.280 252.560 325.570 ;
        RECT 254.510 323.720 254.740 325.570 ;
        RECT 262.800 323.720 263.030 325.700 ;
        RECT 271.090 323.720 271.320 325.700 ;
        RECT 272.020 325.650 272.310 325.700 ;
        RECT 273.580 325.670 280.810 325.700 ;
        RECT 254.510 321.280 254.740 322.540 ;
        RECT 262.800 321.280 263.030 322.540 ;
        RECT 271.090 321.280 271.320 322.540 ;
        RECT 273.580 321.280 278.560 325.670 ;
        RECT 280.510 323.720 280.740 325.670 ;
        RECT 288.800 323.720 289.030 325.700 ;
        RECT 297.090 323.720 297.320 325.700 ;
        RECT 298.020 325.650 298.310 325.700 ;
        RECT 280.510 321.280 280.740 322.540 ;
        RECT 288.800 321.280 289.030 322.540 ;
        RECT 297.090 321.280 297.320 322.540 ;
        RECT 299.580 321.280 304.560 325.700 ;
        RECT 39.400 321.250 63.810 321.280 ;
        RECT 64.460 321.250 70.560 321.280 ;
        RECT 39.400 317.450 70.560 321.250 ;
        RECT 72.250 321.250 89.810 321.280 ;
        RECT 90.460 321.250 96.560 321.280 ;
        RECT 72.250 317.450 96.560 321.250 ;
        RECT 98.250 321.250 115.810 321.280 ;
        RECT 116.460 321.250 122.560 321.280 ;
        RECT 98.250 317.450 122.560 321.250 ;
        RECT 124.250 321.250 141.810 321.280 ;
        RECT 142.460 321.250 148.560 321.280 ;
        RECT 124.250 317.450 148.560 321.250 ;
        RECT 150.250 321.250 167.810 321.280 ;
        RECT 168.460 321.250 174.560 321.280 ;
        RECT 150.250 317.450 174.560 321.250 ;
        RECT 176.250 321.250 193.810 321.280 ;
        RECT 194.460 321.250 200.560 321.280 ;
        RECT 176.250 317.450 200.560 321.250 ;
        RECT 202.250 321.250 219.810 321.280 ;
        RECT 220.460 321.250 226.560 321.280 ;
        RECT 202.250 317.450 226.560 321.250 ;
        RECT 228.250 321.250 245.810 321.280 ;
        RECT 246.460 321.250 252.560 321.280 ;
        RECT 228.250 317.450 252.560 321.250 ;
        RECT 254.250 321.250 271.810 321.280 ;
        RECT 272.460 321.250 278.560 321.280 ;
        RECT 254.250 317.450 278.560 321.250 ;
        RECT 280.250 321.250 297.810 321.280 ;
        RECT 298.460 321.250 304.560 321.280 ;
        RECT 280.250 317.450 304.560 321.250 ;
        RECT 39.400 317.390 50.910 317.450 ;
        RECT 39.400 313.020 44.730 317.390 ;
        RECT 46.510 315.540 46.740 317.390 ;
        RECT 54.800 315.540 55.030 317.450 ;
        RECT 63.090 315.540 63.320 317.450 ;
        RECT 64.020 317.410 64.310 317.450 ;
        RECT 46.510 313.030 46.740 314.360 ;
        RECT 54.800 313.030 55.030 314.360 ;
        RECT 63.090 313.030 63.320 314.360 ;
        RECT 65.580 313.030 70.560 317.450 ;
        RECT 72.510 315.540 72.740 317.450 ;
        RECT 80.800 315.540 81.030 317.450 ;
        RECT 89.090 315.540 89.320 317.450 ;
        RECT 90.020 317.410 90.310 317.450 ;
        RECT 72.510 313.030 72.740 314.360 ;
        RECT 80.800 313.030 81.030 314.360 ;
        RECT 89.090 313.030 89.320 314.360 ;
        RECT 91.580 313.030 96.560 317.450 ;
        RECT 98.510 315.540 98.740 317.450 ;
        RECT 106.800 315.540 107.030 317.450 ;
        RECT 115.090 315.540 115.320 317.450 ;
        RECT 116.020 317.410 116.310 317.450 ;
        RECT 98.510 313.030 98.740 314.360 ;
        RECT 106.800 313.030 107.030 314.360 ;
        RECT 115.090 313.030 115.320 314.360 ;
        RECT 117.580 313.030 122.560 317.450 ;
        RECT 124.510 315.540 124.740 317.450 ;
        RECT 132.800 315.540 133.030 317.450 ;
        RECT 141.090 315.540 141.320 317.450 ;
        RECT 142.020 317.410 142.310 317.450 ;
        RECT 124.510 313.030 124.740 314.360 ;
        RECT 132.800 313.030 133.030 314.360 ;
        RECT 141.090 313.030 141.320 314.360 ;
        RECT 143.580 313.030 148.560 317.450 ;
        RECT 150.510 315.540 150.740 317.450 ;
        RECT 158.800 315.540 159.030 317.450 ;
        RECT 167.090 315.540 167.320 317.450 ;
        RECT 168.020 317.410 168.310 317.450 ;
        RECT 150.510 313.030 150.740 314.360 ;
        RECT 158.800 313.030 159.030 314.360 ;
        RECT 167.090 313.030 167.320 314.360 ;
        RECT 169.580 313.030 174.560 317.450 ;
        RECT 176.510 315.540 176.740 317.450 ;
        RECT 184.800 315.540 185.030 317.450 ;
        RECT 193.090 315.540 193.320 317.450 ;
        RECT 194.020 317.410 194.310 317.450 ;
        RECT 176.510 313.030 176.740 314.360 ;
        RECT 184.800 313.030 185.030 314.360 ;
        RECT 193.090 313.030 193.320 314.360 ;
        RECT 195.580 313.030 200.560 317.450 ;
        RECT 202.510 315.540 202.740 317.450 ;
        RECT 210.800 315.540 211.030 317.450 ;
        RECT 219.090 315.540 219.320 317.450 ;
        RECT 220.020 317.410 220.310 317.450 ;
        RECT 202.510 313.030 202.740 314.360 ;
        RECT 210.800 313.030 211.030 314.360 ;
        RECT 219.090 313.030 219.320 314.360 ;
        RECT 221.580 313.030 226.560 317.450 ;
        RECT 228.510 315.540 228.740 317.450 ;
        RECT 236.800 315.540 237.030 317.450 ;
        RECT 245.090 315.540 245.320 317.450 ;
        RECT 246.020 317.410 246.310 317.450 ;
        RECT 228.510 313.030 228.740 314.360 ;
        RECT 236.800 313.030 237.030 314.360 ;
        RECT 245.090 313.030 245.320 314.360 ;
        RECT 247.580 313.030 252.560 317.450 ;
        RECT 254.510 315.540 254.740 317.450 ;
        RECT 262.800 315.540 263.030 317.450 ;
        RECT 271.090 315.540 271.320 317.450 ;
        RECT 272.020 317.410 272.310 317.450 ;
        RECT 254.510 313.030 254.740 314.360 ;
        RECT 262.800 313.030 263.030 314.360 ;
        RECT 271.090 313.030 271.320 314.360 ;
        RECT 273.580 313.030 278.560 317.450 ;
        RECT 280.510 315.540 280.740 317.450 ;
        RECT 288.800 315.540 289.030 317.450 ;
        RECT 297.090 315.540 297.320 317.450 ;
        RECT 298.020 317.410 298.310 317.450 ;
        RECT 280.510 313.030 280.740 314.360 ;
        RECT 288.800 313.030 289.030 314.360 ;
        RECT 297.090 313.030 297.320 314.360 ;
        RECT 299.580 313.030 304.560 317.450 ;
        RECT 46.250 313.020 63.810 313.030 ;
        RECT 39.400 313.010 63.810 313.020 ;
        RECT 64.460 313.010 70.560 313.030 ;
        RECT 39.400 309.210 70.560 313.010 ;
        RECT 39.400 309.200 63.870 309.210 ;
        RECT 64.500 309.200 70.560 309.210 ;
        RECT 72.250 313.010 89.810 313.030 ;
        RECT 90.460 313.010 96.560 313.030 ;
        RECT 72.250 309.210 96.560 313.010 ;
        RECT 72.250 309.200 89.870 309.210 ;
        RECT 90.500 309.200 96.560 309.210 ;
        RECT 98.250 313.010 115.810 313.030 ;
        RECT 116.460 313.010 122.560 313.030 ;
        RECT 98.250 309.210 122.560 313.010 ;
        RECT 98.250 309.200 115.870 309.210 ;
        RECT 116.500 309.200 122.560 309.210 ;
        RECT 124.250 313.010 141.810 313.030 ;
        RECT 142.460 313.010 148.560 313.030 ;
        RECT 124.250 309.210 148.560 313.010 ;
        RECT 124.250 309.200 141.870 309.210 ;
        RECT 142.500 309.200 148.560 309.210 ;
        RECT 150.250 313.010 167.810 313.030 ;
        RECT 168.460 313.010 174.560 313.030 ;
        RECT 150.250 309.210 174.560 313.010 ;
        RECT 150.250 309.200 167.870 309.210 ;
        RECT 168.500 309.200 174.560 309.210 ;
        RECT 176.250 313.010 193.810 313.030 ;
        RECT 194.460 313.010 200.560 313.030 ;
        RECT 176.250 309.210 200.560 313.010 ;
        RECT 176.250 309.200 193.870 309.210 ;
        RECT 194.500 309.200 200.560 309.210 ;
        RECT 202.250 313.010 219.810 313.030 ;
        RECT 220.460 313.010 226.560 313.030 ;
        RECT 202.250 309.210 226.560 313.010 ;
        RECT 202.250 309.200 219.870 309.210 ;
        RECT 220.500 309.200 226.560 309.210 ;
        RECT 228.250 313.010 245.810 313.030 ;
        RECT 246.460 313.010 252.560 313.030 ;
        RECT 228.250 309.210 252.560 313.010 ;
        RECT 228.250 309.200 245.870 309.210 ;
        RECT 246.500 309.200 252.560 309.210 ;
        RECT 254.250 313.010 271.810 313.030 ;
        RECT 272.460 313.010 278.560 313.030 ;
        RECT 254.250 309.210 278.560 313.010 ;
        RECT 254.250 309.200 271.870 309.210 ;
        RECT 272.500 309.200 278.560 309.210 ;
        RECT 280.250 313.010 297.810 313.030 ;
        RECT 298.460 313.010 304.560 313.030 ;
        RECT 280.250 309.210 304.560 313.010 ;
        RECT 280.250 309.200 297.870 309.210 ;
        RECT 298.500 309.200 304.560 309.210 ;
        RECT 39.400 309.100 48.360 309.200 ;
        RECT 39.400 304.590 44.730 309.100 ;
        RECT 46.510 307.360 46.740 309.100 ;
        RECT 54.800 307.360 55.030 309.200 ;
        RECT 63.090 307.360 63.320 309.200 ;
        RECT 46.510 304.590 46.740 306.180 ;
        RECT 39.400 304.530 48.250 304.590 ;
        RECT 54.800 304.530 55.030 306.180 ;
        RECT 63.090 304.530 63.320 306.180 ;
        RECT 64.020 304.530 64.300 304.540 ;
        RECT 65.580 304.530 70.560 309.200 ;
        RECT 72.510 307.360 72.740 309.200 ;
        RECT 80.800 307.360 81.030 309.200 ;
        RECT 89.090 307.360 89.320 309.200 ;
        RECT 72.510 304.530 72.740 306.180 ;
        RECT 80.800 304.530 81.030 306.180 ;
        RECT 89.090 304.530 89.320 306.180 ;
        RECT 90.020 304.530 90.300 304.540 ;
        RECT 91.580 304.530 96.560 309.200 ;
        RECT 98.510 307.360 98.740 309.200 ;
        RECT 106.800 307.360 107.030 309.200 ;
        RECT 115.090 307.360 115.320 309.200 ;
        RECT 98.510 304.530 98.740 306.180 ;
        RECT 106.800 304.530 107.030 306.180 ;
        RECT 115.090 304.530 115.320 306.180 ;
        RECT 116.020 304.530 116.300 304.540 ;
        RECT 117.580 304.530 122.560 309.200 ;
        RECT 124.510 307.360 124.740 309.200 ;
        RECT 132.800 307.360 133.030 309.200 ;
        RECT 141.090 307.360 141.320 309.200 ;
        RECT 124.510 304.530 124.740 306.180 ;
        RECT 132.800 304.530 133.030 306.180 ;
        RECT 141.090 304.530 141.320 306.180 ;
        RECT 142.020 304.530 142.300 304.540 ;
        RECT 143.580 304.530 148.560 309.200 ;
        RECT 150.510 307.360 150.740 309.200 ;
        RECT 158.800 307.360 159.030 309.200 ;
        RECT 167.090 307.360 167.320 309.200 ;
        RECT 150.510 304.530 150.740 306.180 ;
        RECT 158.800 304.530 159.030 306.180 ;
        RECT 167.090 304.530 167.320 306.180 ;
        RECT 168.020 304.530 168.300 304.540 ;
        RECT 169.580 304.530 174.560 309.200 ;
        RECT 176.510 307.360 176.740 309.200 ;
        RECT 184.800 307.360 185.030 309.200 ;
        RECT 193.090 307.360 193.320 309.200 ;
        RECT 176.510 304.530 176.740 306.180 ;
        RECT 184.800 304.530 185.030 306.180 ;
        RECT 193.090 304.530 193.320 306.180 ;
        RECT 194.020 304.530 194.300 304.540 ;
        RECT 195.580 304.530 200.560 309.200 ;
        RECT 202.510 307.360 202.740 309.200 ;
        RECT 210.800 307.360 211.030 309.200 ;
        RECT 219.090 307.360 219.320 309.200 ;
        RECT 202.510 304.530 202.740 306.180 ;
        RECT 210.800 304.530 211.030 306.180 ;
        RECT 219.090 304.530 219.320 306.180 ;
        RECT 220.020 304.530 220.300 304.540 ;
        RECT 221.580 304.530 226.560 309.200 ;
        RECT 228.510 307.360 228.740 309.200 ;
        RECT 236.800 307.360 237.030 309.200 ;
        RECT 245.090 307.360 245.320 309.200 ;
        RECT 228.510 304.530 228.740 306.180 ;
        RECT 236.800 304.530 237.030 306.180 ;
        RECT 245.090 304.530 245.320 306.180 ;
        RECT 246.020 304.530 246.300 304.540 ;
        RECT 247.580 304.530 252.560 309.200 ;
        RECT 254.510 307.360 254.740 309.200 ;
        RECT 262.800 307.360 263.030 309.200 ;
        RECT 271.090 307.360 271.320 309.200 ;
        RECT 254.510 304.530 254.740 306.180 ;
        RECT 262.800 304.530 263.030 306.180 ;
        RECT 271.090 304.530 271.320 306.180 ;
        RECT 272.020 304.530 272.300 304.540 ;
        RECT 273.580 304.530 278.560 309.200 ;
        RECT 280.510 307.360 280.740 309.200 ;
        RECT 288.800 307.360 289.030 309.200 ;
        RECT 297.090 307.360 297.320 309.200 ;
        RECT 280.510 304.530 280.740 306.180 ;
        RECT 288.800 304.530 289.030 306.180 ;
        RECT 297.090 304.530 297.320 306.180 ;
        RECT 298.020 304.530 298.300 304.540 ;
        RECT 299.580 304.530 304.560 309.200 ;
        RECT 39.400 300.710 70.560 304.530 ;
        RECT 39.400 300.700 63.890 300.710 ;
        RECT 64.520 300.700 70.560 300.710 ;
        RECT 72.250 300.710 96.560 304.530 ;
        RECT 72.250 300.700 89.890 300.710 ;
        RECT 90.520 300.700 96.560 300.710 ;
        RECT 98.250 300.710 122.560 304.530 ;
        RECT 98.250 300.700 115.890 300.710 ;
        RECT 116.520 300.700 122.560 300.710 ;
        RECT 124.250 300.710 148.560 304.530 ;
        RECT 124.250 300.700 141.890 300.710 ;
        RECT 142.520 300.700 148.560 300.710 ;
        RECT 150.250 300.710 174.560 304.530 ;
        RECT 150.250 300.700 167.890 300.710 ;
        RECT 168.520 300.700 174.560 300.710 ;
        RECT 176.250 300.710 200.560 304.530 ;
        RECT 176.250 300.700 193.890 300.710 ;
        RECT 194.520 300.700 200.560 300.710 ;
        RECT 202.250 300.710 226.560 304.530 ;
        RECT 202.250 300.700 219.890 300.710 ;
        RECT 220.520 300.700 226.560 300.710 ;
        RECT 228.250 300.710 252.560 304.530 ;
        RECT 228.250 300.700 245.890 300.710 ;
        RECT 246.520 300.700 252.560 300.710 ;
        RECT 254.250 300.710 278.560 304.530 ;
        RECT 254.250 300.700 271.890 300.710 ;
        RECT 272.520 300.700 278.560 300.710 ;
        RECT 280.250 300.710 304.560 304.530 ;
        RECT 280.250 300.700 297.890 300.710 ;
        RECT 298.520 300.700 304.560 300.710 ;
        RECT 39.400 300.670 48.250 300.700 ;
        RECT 39.400 295.940 44.730 300.670 ;
        RECT 46.510 299.180 46.740 300.670 ;
        RECT 54.800 299.180 55.030 300.700 ;
        RECT 63.090 299.180 63.320 300.700 ;
        RECT 46.510 296.030 46.740 298.000 ;
        RECT 54.800 296.030 55.030 298.000 ;
        RECT 63.090 296.030 63.320 298.000 ;
        RECT 64.020 296.030 64.300 296.040 ;
        RECT 65.580 296.030 70.560 300.700 ;
        RECT 72.510 299.180 72.740 300.700 ;
        RECT 80.800 299.180 81.030 300.700 ;
        RECT 89.090 299.180 89.320 300.700 ;
        RECT 72.510 296.030 72.740 298.000 ;
        RECT 80.800 296.030 81.030 298.000 ;
        RECT 89.090 296.030 89.320 298.000 ;
        RECT 90.020 296.030 90.300 296.040 ;
        RECT 91.580 296.030 96.560 300.700 ;
        RECT 98.510 299.180 98.740 300.700 ;
        RECT 106.800 299.180 107.030 300.700 ;
        RECT 115.090 299.180 115.320 300.700 ;
        RECT 98.510 296.030 98.740 298.000 ;
        RECT 106.800 296.030 107.030 298.000 ;
        RECT 115.090 296.030 115.320 298.000 ;
        RECT 116.020 296.030 116.300 296.040 ;
        RECT 117.580 296.030 122.560 300.700 ;
        RECT 124.510 299.180 124.740 300.700 ;
        RECT 132.800 299.180 133.030 300.700 ;
        RECT 141.090 299.180 141.320 300.700 ;
        RECT 124.510 296.030 124.740 298.000 ;
        RECT 132.800 296.030 133.030 298.000 ;
        RECT 141.090 296.030 141.320 298.000 ;
        RECT 142.020 296.030 142.300 296.040 ;
        RECT 143.580 296.030 148.560 300.700 ;
        RECT 150.510 299.180 150.740 300.700 ;
        RECT 158.800 299.180 159.030 300.700 ;
        RECT 167.090 299.180 167.320 300.700 ;
        RECT 150.510 296.030 150.740 298.000 ;
        RECT 158.800 296.030 159.030 298.000 ;
        RECT 167.090 296.030 167.320 298.000 ;
        RECT 168.020 296.030 168.300 296.040 ;
        RECT 169.580 296.030 174.560 300.700 ;
        RECT 176.510 299.180 176.740 300.700 ;
        RECT 184.800 299.180 185.030 300.700 ;
        RECT 193.090 299.180 193.320 300.700 ;
        RECT 176.510 296.030 176.740 298.000 ;
        RECT 184.800 296.030 185.030 298.000 ;
        RECT 193.090 296.030 193.320 298.000 ;
        RECT 194.020 296.030 194.300 296.040 ;
        RECT 195.580 296.030 200.560 300.700 ;
        RECT 202.510 299.180 202.740 300.700 ;
        RECT 210.800 299.180 211.030 300.700 ;
        RECT 219.090 299.180 219.320 300.700 ;
        RECT 202.510 296.030 202.740 298.000 ;
        RECT 210.800 296.030 211.030 298.000 ;
        RECT 219.090 296.030 219.320 298.000 ;
        RECT 220.020 296.030 220.300 296.040 ;
        RECT 221.580 296.030 226.560 300.700 ;
        RECT 228.510 299.180 228.740 300.700 ;
        RECT 236.800 299.180 237.030 300.700 ;
        RECT 245.090 299.180 245.320 300.700 ;
        RECT 228.510 296.030 228.740 298.000 ;
        RECT 236.800 296.030 237.030 298.000 ;
        RECT 245.090 296.030 245.320 298.000 ;
        RECT 246.020 296.030 246.300 296.040 ;
        RECT 247.580 296.030 252.560 300.700 ;
        RECT 254.510 299.180 254.740 300.700 ;
        RECT 262.800 299.180 263.030 300.700 ;
        RECT 271.090 299.180 271.320 300.700 ;
        RECT 254.510 296.030 254.740 298.000 ;
        RECT 262.800 296.030 263.030 298.000 ;
        RECT 271.090 296.030 271.320 298.000 ;
        RECT 272.020 296.030 272.300 296.040 ;
        RECT 273.580 296.030 278.560 300.700 ;
        RECT 280.510 299.180 280.740 300.700 ;
        RECT 288.800 299.180 289.030 300.700 ;
        RECT 297.090 299.180 297.320 300.700 ;
        RECT 280.510 296.030 280.740 298.000 ;
        RECT 288.800 296.030 289.030 298.000 ;
        RECT 297.090 296.030 297.320 298.000 ;
        RECT 298.020 296.030 298.300 296.040 ;
        RECT 299.580 296.030 304.560 300.700 ;
        RECT 46.250 295.940 70.560 296.030 ;
        RECT 39.400 292.200 70.560 295.940 ;
        RECT 72.250 292.200 96.560 296.030 ;
        RECT 98.250 292.200 122.560 296.030 ;
        RECT 124.250 292.200 148.560 296.030 ;
        RECT 150.250 292.200 174.560 296.030 ;
        RECT 176.250 292.200 200.560 296.030 ;
        RECT 202.250 292.200 226.560 296.030 ;
        RECT 228.250 292.200 252.560 296.030 ;
        RECT 254.250 292.200 278.560 296.030 ;
        RECT 280.250 292.200 304.560 296.030 ;
        RECT 39.400 292.020 49.610 292.200 ;
        RECT 39.400 288.000 44.730 292.020 ;
        RECT 46.510 291.000 46.740 292.020 ;
        RECT 54.800 291.000 55.030 292.200 ;
        RECT 63.090 291.000 63.320 292.200 ;
        RECT 64.020 292.140 64.310 292.200 ;
        RECT 46.510 288.030 46.740 289.820 ;
        RECT 54.800 288.030 55.030 289.820 ;
        RECT 63.090 288.030 63.320 289.820 ;
        RECT 65.580 288.030 70.560 292.200 ;
        RECT 72.510 291.000 72.740 292.200 ;
        RECT 80.800 291.000 81.030 292.200 ;
        RECT 89.090 291.000 89.320 292.200 ;
        RECT 90.020 292.140 90.310 292.200 ;
        RECT 72.510 288.030 72.740 289.820 ;
        RECT 80.800 288.030 81.030 289.820 ;
        RECT 89.090 288.030 89.320 289.820 ;
        RECT 91.580 288.030 96.560 292.200 ;
        RECT 98.510 291.000 98.740 292.200 ;
        RECT 106.800 291.000 107.030 292.200 ;
        RECT 115.090 291.000 115.320 292.200 ;
        RECT 116.020 292.140 116.310 292.200 ;
        RECT 98.510 288.030 98.740 289.820 ;
        RECT 106.800 288.030 107.030 289.820 ;
        RECT 115.090 288.030 115.320 289.820 ;
        RECT 117.580 288.030 122.560 292.200 ;
        RECT 124.510 291.000 124.740 292.200 ;
        RECT 132.800 291.000 133.030 292.200 ;
        RECT 141.090 291.000 141.320 292.200 ;
        RECT 142.020 292.140 142.310 292.200 ;
        RECT 124.510 288.030 124.740 289.820 ;
        RECT 132.800 288.030 133.030 289.820 ;
        RECT 141.090 288.030 141.320 289.820 ;
        RECT 143.580 288.030 148.560 292.200 ;
        RECT 150.510 291.000 150.740 292.200 ;
        RECT 158.800 291.000 159.030 292.200 ;
        RECT 167.090 291.000 167.320 292.200 ;
        RECT 168.020 292.140 168.310 292.200 ;
        RECT 150.510 288.030 150.740 289.820 ;
        RECT 158.800 288.030 159.030 289.820 ;
        RECT 167.090 288.030 167.320 289.820 ;
        RECT 169.580 288.030 174.560 292.200 ;
        RECT 176.510 291.000 176.740 292.200 ;
        RECT 184.800 291.000 185.030 292.200 ;
        RECT 193.090 291.000 193.320 292.200 ;
        RECT 194.020 292.140 194.310 292.200 ;
        RECT 176.510 288.030 176.740 289.820 ;
        RECT 184.800 288.030 185.030 289.820 ;
        RECT 193.090 288.030 193.320 289.820 ;
        RECT 195.580 288.030 200.560 292.200 ;
        RECT 202.510 291.000 202.740 292.200 ;
        RECT 210.800 291.000 211.030 292.200 ;
        RECT 219.090 291.000 219.320 292.200 ;
        RECT 220.020 292.140 220.310 292.200 ;
        RECT 202.510 288.030 202.740 289.820 ;
        RECT 210.800 288.030 211.030 289.820 ;
        RECT 219.090 288.030 219.320 289.820 ;
        RECT 221.580 288.030 226.560 292.200 ;
        RECT 228.510 291.000 228.740 292.200 ;
        RECT 236.800 291.000 237.030 292.200 ;
        RECT 245.090 291.000 245.320 292.200 ;
        RECT 246.020 292.140 246.310 292.200 ;
        RECT 228.510 288.030 228.740 289.820 ;
        RECT 236.800 288.030 237.030 289.820 ;
        RECT 245.090 288.030 245.320 289.820 ;
        RECT 247.580 288.030 252.560 292.200 ;
        RECT 254.510 291.000 254.740 292.200 ;
        RECT 262.800 291.000 263.030 292.200 ;
        RECT 271.090 291.000 271.320 292.200 ;
        RECT 272.020 292.140 272.310 292.200 ;
        RECT 254.510 288.030 254.740 289.820 ;
        RECT 262.800 288.030 263.030 289.820 ;
        RECT 271.090 288.030 271.320 289.820 ;
        RECT 273.580 288.030 278.560 292.200 ;
        RECT 280.510 291.000 280.740 292.200 ;
        RECT 288.800 291.000 289.030 292.200 ;
        RECT 297.090 291.000 297.320 292.200 ;
        RECT 298.020 292.140 298.310 292.200 ;
        RECT 280.510 288.030 280.740 289.820 ;
        RECT 288.800 288.030 289.030 289.820 ;
        RECT 297.090 288.030 297.320 289.820 ;
        RECT 299.580 288.030 304.560 292.200 ;
        RECT 46.250 288.000 63.890 288.030 ;
        RECT 64.460 288.000 70.560 288.030 ;
        RECT 39.400 284.200 70.560 288.000 ;
        RECT 72.250 288.000 89.890 288.030 ;
        RECT 90.460 288.000 96.560 288.030 ;
        RECT 72.250 284.200 96.560 288.000 ;
        RECT 98.250 288.000 115.890 288.030 ;
        RECT 116.460 288.000 122.560 288.030 ;
        RECT 98.250 284.200 122.560 288.000 ;
        RECT 124.250 288.000 141.890 288.030 ;
        RECT 142.460 288.000 148.560 288.030 ;
        RECT 124.250 284.200 148.560 288.000 ;
        RECT 150.250 288.000 167.890 288.030 ;
        RECT 168.460 288.000 174.560 288.030 ;
        RECT 150.250 284.200 174.560 288.000 ;
        RECT 176.250 288.000 193.890 288.030 ;
        RECT 194.460 288.000 200.560 288.030 ;
        RECT 176.250 284.200 200.560 288.000 ;
        RECT 202.250 288.000 219.890 288.030 ;
        RECT 220.460 288.000 226.560 288.030 ;
        RECT 202.250 284.200 226.560 288.000 ;
        RECT 228.250 288.000 245.890 288.030 ;
        RECT 246.460 288.000 252.560 288.030 ;
        RECT 228.250 284.200 252.560 288.000 ;
        RECT 254.250 288.000 271.890 288.030 ;
        RECT 272.460 288.000 278.560 288.030 ;
        RECT 254.250 284.200 278.560 288.000 ;
        RECT 280.250 288.000 297.890 288.030 ;
        RECT 298.460 288.000 304.560 288.030 ;
        RECT 280.250 284.200 304.560 288.000 ;
        RECT 39.400 284.080 50.130 284.200 ;
        RECT 39.400 280.080 44.730 284.080 ;
        RECT 46.510 282.820 46.740 284.080 ;
        RECT 54.800 282.820 55.030 284.200 ;
        RECT 63.090 282.820 63.320 284.200 ;
        RECT 64.020 284.120 64.310 284.200 ;
        RECT 46.510 280.080 46.740 281.640 ;
        RECT 39.400 280.030 49.010 280.080 ;
        RECT 54.800 280.030 55.030 281.640 ;
        RECT 63.090 280.030 63.320 281.640 ;
        RECT 65.580 280.030 70.560 284.200 ;
        RECT 72.510 282.820 72.740 284.200 ;
        RECT 80.800 282.820 81.030 284.200 ;
        RECT 89.090 282.820 89.320 284.200 ;
        RECT 90.020 284.120 90.310 284.200 ;
        RECT 72.510 280.030 72.740 281.640 ;
        RECT 80.800 280.030 81.030 281.640 ;
        RECT 89.090 280.030 89.320 281.640 ;
        RECT 91.580 280.030 96.560 284.200 ;
        RECT 98.510 282.820 98.740 284.200 ;
        RECT 106.800 282.820 107.030 284.200 ;
        RECT 115.090 282.820 115.320 284.200 ;
        RECT 116.020 284.120 116.310 284.200 ;
        RECT 98.510 280.030 98.740 281.640 ;
        RECT 106.800 280.030 107.030 281.640 ;
        RECT 115.090 280.030 115.320 281.640 ;
        RECT 117.580 280.030 122.560 284.200 ;
        RECT 124.510 282.820 124.740 284.200 ;
        RECT 132.800 282.820 133.030 284.200 ;
        RECT 141.090 282.820 141.320 284.200 ;
        RECT 142.020 284.120 142.310 284.200 ;
        RECT 124.510 280.030 124.740 281.640 ;
        RECT 132.800 280.030 133.030 281.640 ;
        RECT 141.090 280.030 141.320 281.640 ;
        RECT 143.580 280.030 148.560 284.200 ;
        RECT 150.510 282.820 150.740 284.200 ;
        RECT 158.800 282.820 159.030 284.200 ;
        RECT 167.090 282.820 167.320 284.200 ;
        RECT 168.020 284.120 168.310 284.200 ;
        RECT 150.510 280.030 150.740 281.640 ;
        RECT 158.800 280.030 159.030 281.640 ;
        RECT 167.090 280.030 167.320 281.640 ;
        RECT 169.580 280.030 174.560 284.200 ;
        RECT 176.510 282.820 176.740 284.200 ;
        RECT 184.800 282.820 185.030 284.200 ;
        RECT 193.090 282.820 193.320 284.200 ;
        RECT 194.020 284.120 194.310 284.200 ;
        RECT 176.510 280.030 176.740 281.640 ;
        RECT 184.800 280.030 185.030 281.640 ;
        RECT 193.090 280.030 193.320 281.640 ;
        RECT 195.580 280.030 200.560 284.200 ;
        RECT 202.510 282.820 202.740 284.200 ;
        RECT 210.800 282.820 211.030 284.200 ;
        RECT 219.090 282.820 219.320 284.200 ;
        RECT 220.020 284.120 220.310 284.200 ;
        RECT 202.510 280.030 202.740 281.640 ;
        RECT 210.800 280.030 211.030 281.640 ;
        RECT 219.090 280.030 219.320 281.640 ;
        RECT 221.580 280.030 226.560 284.200 ;
        RECT 228.510 282.820 228.740 284.200 ;
        RECT 236.800 282.820 237.030 284.200 ;
        RECT 245.090 282.820 245.320 284.200 ;
        RECT 246.020 284.120 246.310 284.200 ;
        RECT 228.510 280.030 228.740 281.640 ;
        RECT 236.800 280.030 237.030 281.640 ;
        RECT 245.090 280.030 245.320 281.640 ;
        RECT 247.580 280.030 252.560 284.200 ;
        RECT 254.510 282.820 254.740 284.200 ;
        RECT 262.800 282.820 263.030 284.200 ;
        RECT 271.090 282.820 271.320 284.200 ;
        RECT 272.020 284.120 272.310 284.200 ;
        RECT 254.510 280.030 254.740 281.640 ;
        RECT 262.800 280.030 263.030 281.640 ;
        RECT 271.090 280.030 271.320 281.640 ;
        RECT 273.580 280.030 278.560 284.200 ;
        RECT 280.510 282.820 280.740 284.200 ;
        RECT 288.800 282.820 289.030 284.200 ;
        RECT 297.090 282.820 297.320 284.200 ;
        RECT 298.020 284.120 298.310 284.200 ;
        RECT 280.510 280.030 280.740 281.640 ;
        RECT 288.800 280.030 289.030 281.640 ;
        RECT 297.090 280.030 297.320 281.640 ;
        RECT 299.580 280.030 304.560 284.200 ;
        RECT 39.400 279.980 63.930 280.030 ;
        RECT 64.500 279.980 70.560 280.030 ;
        RECT 39.400 276.200 70.560 279.980 ;
        RECT 72.250 279.980 89.930 280.030 ;
        RECT 90.500 279.980 96.560 280.030 ;
        RECT 72.250 276.200 96.560 279.980 ;
        RECT 98.250 279.980 115.930 280.030 ;
        RECT 116.500 279.980 122.560 280.030 ;
        RECT 98.250 276.200 122.560 279.980 ;
        RECT 124.250 279.980 141.930 280.030 ;
        RECT 142.500 279.980 148.560 280.030 ;
        RECT 124.250 276.200 148.560 279.980 ;
        RECT 150.250 279.980 167.930 280.030 ;
        RECT 168.500 279.980 174.560 280.030 ;
        RECT 150.250 276.200 174.560 279.980 ;
        RECT 176.250 279.980 193.930 280.030 ;
        RECT 194.500 279.980 200.560 280.030 ;
        RECT 176.250 276.200 200.560 279.980 ;
        RECT 202.250 279.980 219.930 280.030 ;
        RECT 220.500 279.980 226.560 280.030 ;
        RECT 202.250 276.200 226.560 279.980 ;
        RECT 228.250 279.980 245.930 280.030 ;
        RECT 246.500 279.980 252.560 280.030 ;
        RECT 228.250 276.200 252.560 279.980 ;
        RECT 254.250 279.980 271.930 280.030 ;
        RECT 272.500 279.980 278.560 280.030 ;
        RECT 254.250 276.200 278.560 279.980 ;
        RECT 280.250 279.980 297.930 280.030 ;
        RECT 298.500 279.980 304.560 280.030 ;
        RECT 280.250 276.200 304.560 279.980 ;
        RECT 39.400 276.160 49.010 276.200 ;
        RECT 39.400 272.140 44.730 276.160 ;
        RECT 46.510 274.640 46.740 276.160 ;
        RECT 54.800 274.640 55.030 276.200 ;
        RECT 63.090 274.640 63.320 276.200 ;
        RECT 64.020 276.190 64.310 276.200 ;
        RECT 46.510 272.140 46.740 273.460 ;
        RECT 39.400 272.030 48.330 272.140 ;
        RECT 54.800 272.030 55.030 273.460 ;
        RECT 63.090 272.030 63.320 273.460 ;
        RECT 64.020 272.030 64.300 272.050 ;
        RECT 65.580 272.030 70.560 276.200 ;
        RECT 72.510 274.640 72.740 276.200 ;
        RECT 80.800 274.640 81.030 276.200 ;
        RECT 89.090 274.640 89.320 276.200 ;
        RECT 90.020 276.190 90.310 276.200 ;
        RECT 72.510 272.030 72.740 273.460 ;
        RECT 80.800 272.030 81.030 273.460 ;
        RECT 89.090 272.030 89.320 273.460 ;
        RECT 90.020 272.030 90.300 272.050 ;
        RECT 91.580 272.030 96.560 276.200 ;
        RECT 98.510 274.640 98.740 276.200 ;
        RECT 106.800 274.640 107.030 276.200 ;
        RECT 115.090 274.640 115.320 276.200 ;
        RECT 116.020 276.190 116.310 276.200 ;
        RECT 98.510 272.030 98.740 273.460 ;
        RECT 106.800 272.030 107.030 273.460 ;
        RECT 115.090 272.030 115.320 273.460 ;
        RECT 116.020 272.030 116.300 272.050 ;
        RECT 117.580 272.030 122.560 276.200 ;
        RECT 124.510 274.640 124.740 276.200 ;
        RECT 132.800 274.640 133.030 276.200 ;
        RECT 141.090 274.640 141.320 276.200 ;
        RECT 142.020 276.190 142.310 276.200 ;
        RECT 124.510 272.030 124.740 273.460 ;
        RECT 132.800 272.030 133.030 273.460 ;
        RECT 141.090 272.030 141.320 273.460 ;
        RECT 142.020 272.030 142.300 272.050 ;
        RECT 143.580 272.030 148.560 276.200 ;
        RECT 150.510 274.640 150.740 276.200 ;
        RECT 158.800 274.640 159.030 276.200 ;
        RECT 167.090 274.640 167.320 276.200 ;
        RECT 168.020 276.190 168.310 276.200 ;
        RECT 150.510 272.030 150.740 273.460 ;
        RECT 158.800 272.030 159.030 273.460 ;
        RECT 167.090 272.030 167.320 273.460 ;
        RECT 168.020 272.030 168.300 272.050 ;
        RECT 169.580 272.030 174.560 276.200 ;
        RECT 176.510 274.640 176.740 276.200 ;
        RECT 184.800 274.640 185.030 276.200 ;
        RECT 193.090 274.640 193.320 276.200 ;
        RECT 194.020 276.190 194.310 276.200 ;
        RECT 176.510 272.030 176.740 273.460 ;
        RECT 184.800 272.030 185.030 273.460 ;
        RECT 193.090 272.030 193.320 273.460 ;
        RECT 194.020 272.030 194.300 272.050 ;
        RECT 195.580 272.030 200.560 276.200 ;
        RECT 202.510 274.640 202.740 276.200 ;
        RECT 210.800 274.640 211.030 276.200 ;
        RECT 219.090 274.640 219.320 276.200 ;
        RECT 220.020 276.190 220.310 276.200 ;
        RECT 202.510 272.030 202.740 273.460 ;
        RECT 210.800 272.030 211.030 273.460 ;
        RECT 219.090 272.030 219.320 273.460 ;
        RECT 220.020 272.030 220.300 272.050 ;
        RECT 221.580 272.030 226.560 276.200 ;
        RECT 228.510 274.640 228.740 276.200 ;
        RECT 236.800 274.640 237.030 276.200 ;
        RECT 245.090 274.640 245.320 276.200 ;
        RECT 246.020 276.190 246.310 276.200 ;
        RECT 228.510 272.030 228.740 273.460 ;
        RECT 236.800 272.030 237.030 273.460 ;
        RECT 245.090 272.030 245.320 273.460 ;
        RECT 246.020 272.030 246.300 272.050 ;
        RECT 247.580 272.030 252.560 276.200 ;
        RECT 254.510 274.640 254.740 276.200 ;
        RECT 262.800 274.640 263.030 276.200 ;
        RECT 271.090 274.640 271.320 276.200 ;
        RECT 272.020 276.190 272.310 276.200 ;
        RECT 254.510 272.030 254.740 273.460 ;
        RECT 262.800 272.030 263.030 273.460 ;
        RECT 271.090 272.030 271.320 273.460 ;
        RECT 272.020 272.030 272.300 272.050 ;
        RECT 273.580 272.030 278.560 276.200 ;
        RECT 280.510 274.640 280.740 276.200 ;
        RECT 288.800 274.640 289.030 276.200 ;
        RECT 297.090 274.640 297.320 276.200 ;
        RECT 298.020 276.190 298.310 276.200 ;
        RECT 280.510 272.030 280.740 273.460 ;
        RECT 288.800 272.030 289.030 273.460 ;
        RECT 297.090 272.030 297.320 273.460 ;
        RECT 298.020 272.030 298.300 272.050 ;
        RECT 299.580 272.030 304.560 276.200 ;
        RECT 39.400 268.220 70.560 272.030 ;
        RECT 39.400 264.280 44.730 268.220 ;
        RECT 46.250 268.200 70.560 268.220 ;
        RECT 72.250 268.200 96.560 272.030 ;
        RECT 98.250 268.200 122.560 272.030 ;
        RECT 124.250 268.200 148.560 272.030 ;
        RECT 150.250 268.200 174.560 272.030 ;
        RECT 176.250 268.200 200.560 272.030 ;
        RECT 202.250 268.200 226.560 272.030 ;
        RECT 228.250 268.200 252.560 272.030 ;
        RECT 254.250 268.200 278.560 272.030 ;
        RECT 280.250 268.200 304.560 272.030 ;
        RECT 46.510 266.460 46.740 268.200 ;
        RECT 54.800 266.460 55.030 268.200 ;
        RECT 63.090 266.460 63.320 268.200 ;
        RECT 64.020 268.190 64.310 268.200 ;
        RECT 46.510 264.280 46.740 265.280 ;
        RECT 39.400 264.030 49.770 264.280 ;
        RECT 54.800 264.030 55.030 265.280 ;
        RECT 63.090 264.030 63.320 265.280 ;
        RECT 64.020 264.030 64.300 264.050 ;
        RECT 65.580 264.030 70.560 268.200 ;
        RECT 72.510 266.460 72.740 268.200 ;
        RECT 80.800 266.460 81.030 268.200 ;
        RECT 89.090 266.460 89.320 268.200 ;
        RECT 90.020 268.190 90.310 268.200 ;
        RECT 72.510 264.030 72.740 265.280 ;
        RECT 80.800 264.030 81.030 265.280 ;
        RECT 89.090 264.030 89.320 265.280 ;
        RECT 90.020 264.030 90.300 264.050 ;
        RECT 91.580 264.030 96.560 268.200 ;
        RECT 98.510 266.460 98.740 268.200 ;
        RECT 106.800 266.460 107.030 268.200 ;
        RECT 115.090 266.460 115.320 268.200 ;
        RECT 116.020 268.190 116.310 268.200 ;
        RECT 98.510 264.030 98.740 265.280 ;
        RECT 106.800 264.030 107.030 265.280 ;
        RECT 115.090 264.030 115.320 265.280 ;
        RECT 116.020 264.030 116.300 264.050 ;
        RECT 117.580 264.030 122.560 268.200 ;
        RECT 124.510 266.460 124.740 268.200 ;
        RECT 132.800 266.460 133.030 268.200 ;
        RECT 141.090 266.460 141.320 268.200 ;
        RECT 142.020 268.190 142.310 268.200 ;
        RECT 124.510 264.030 124.740 265.280 ;
        RECT 132.800 264.030 133.030 265.280 ;
        RECT 141.090 264.030 141.320 265.280 ;
        RECT 142.020 264.030 142.300 264.050 ;
        RECT 143.580 264.030 148.560 268.200 ;
        RECT 150.510 266.460 150.740 268.200 ;
        RECT 158.800 266.460 159.030 268.200 ;
        RECT 167.090 266.460 167.320 268.200 ;
        RECT 168.020 268.190 168.310 268.200 ;
        RECT 150.510 264.030 150.740 265.280 ;
        RECT 158.800 264.030 159.030 265.280 ;
        RECT 167.090 264.030 167.320 265.280 ;
        RECT 168.020 264.030 168.300 264.050 ;
        RECT 169.580 264.030 174.560 268.200 ;
        RECT 176.510 266.460 176.740 268.200 ;
        RECT 184.800 266.460 185.030 268.200 ;
        RECT 193.090 266.460 193.320 268.200 ;
        RECT 194.020 268.190 194.310 268.200 ;
        RECT 176.510 264.030 176.740 265.280 ;
        RECT 184.800 264.030 185.030 265.280 ;
        RECT 193.090 264.030 193.320 265.280 ;
        RECT 194.020 264.030 194.300 264.050 ;
        RECT 195.580 264.030 200.560 268.200 ;
        RECT 202.510 266.460 202.740 268.200 ;
        RECT 210.800 266.460 211.030 268.200 ;
        RECT 219.090 266.460 219.320 268.200 ;
        RECT 220.020 268.190 220.310 268.200 ;
        RECT 202.510 264.030 202.740 265.280 ;
        RECT 210.800 264.030 211.030 265.280 ;
        RECT 219.090 264.030 219.320 265.280 ;
        RECT 220.020 264.030 220.300 264.050 ;
        RECT 221.580 264.030 226.560 268.200 ;
        RECT 228.510 266.460 228.740 268.200 ;
        RECT 236.800 266.460 237.030 268.200 ;
        RECT 245.090 266.460 245.320 268.200 ;
        RECT 246.020 268.190 246.310 268.200 ;
        RECT 228.510 264.030 228.740 265.280 ;
        RECT 236.800 264.030 237.030 265.280 ;
        RECT 245.090 264.030 245.320 265.280 ;
        RECT 246.020 264.030 246.300 264.050 ;
        RECT 247.580 264.030 252.560 268.200 ;
        RECT 254.510 266.460 254.740 268.200 ;
        RECT 262.800 266.460 263.030 268.200 ;
        RECT 271.090 266.460 271.320 268.200 ;
        RECT 272.020 268.190 272.310 268.200 ;
        RECT 254.510 264.030 254.740 265.280 ;
        RECT 262.800 264.030 263.030 265.280 ;
        RECT 271.090 264.030 271.320 265.280 ;
        RECT 272.020 264.030 272.300 264.050 ;
        RECT 273.580 264.030 278.560 268.200 ;
        RECT 280.510 266.460 280.740 268.200 ;
        RECT 288.800 266.460 289.030 268.200 ;
        RECT 297.090 266.460 297.320 268.200 ;
        RECT 298.020 268.190 298.310 268.200 ;
        RECT 280.510 264.030 280.740 265.280 ;
        RECT 288.800 264.030 289.030 265.280 ;
        RECT 297.090 264.030 297.320 265.280 ;
        RECT 298.020 264.030 298.300 264.050 ;
        RECT 299.580 264.030 304.560 268.200 ;
        RECT 39.400 260.200 70.560 264.030 ;
        RECT 72.250 260.200 96.560 264.030 ;
        RECT 98.250 260.200 122.560 264.030 ;
        RECT 124.250 260.200 148.560 264.030 ;
        RECT 150.250 260.200 174.560 264.030 ;
        RECT 176.250 260.200 200.560 264.030 ;
        RECT 202.250 260.200 226.560 264.030 ;
        RECT 228.250 260.200 252.560 264.030 ;
        RECT 254.250 260.200 278.560 264.030 ;
        RECT 280.250 260.200 304.560 264.030 ;
        RECT 39.400 259.660 49.770 260.200 ;
        RECT 39.400 255.960 44.730 259.660 ;
        RECT 46.510 258.280 46.740 259.660 ;
        RECT 54.800 258.280 55.030 260.200 ;
        RECT 63.090 258.280 63.320 260.200 ;
        RECT 64.020 260.180 64.340 260.200 ;
        RECT 46.510 256.030 46.740 257.100 ;
        RECT 54.800 256.030 55.030 257.100 ;
        RECT 63.090 256.030 63.320 257.100 ;
        RECT 64.020 256.030 64.300 256.040 ;
        RECT 65.580 256.030 70.560 260.200 ;
        RECT 72.510 258.280 72.740 260.200 ;
        RECT 80.800 258.280 81.030 260.200 ;
        RECT 89.090 258.280 89.320 260.200 ;
        RECT 90.020 260.180 90.340 260.200 ;
        RECT 72.510 256.030 72.740 257.100 ;
        RECT 80.800 256.030 81.030 257.100 ;
        RECT 89.090 256.030 89.320 257.100 ;
        RECT 90.020 256.030 90.300 256.040 ;
        RECT 91.580 256.030 96.560 260.200 ;
        RECT 98.510 258.280 98.740 260.200 ;
        RECT 106.800 258.280 107.030 260.200 ;
        RECT 115.090 258.280 115.320 260.200 ;
        RECT 116.020 260.180 116.340 260.200 ;
        RECT 98.510 256.030 98.740 257.100 ;
        RECT 106.800 256.030 107.030 257.100 ;
        RECT 115.090 256.030 115.320 257.100 ;
        RECT 116.020 256.030 116.300 256.040 ;
        RECT 117.580 256.030 122.560 260.200 ;
        RECT 124.510 258.280 124.740 260.200 ;
        RECT 132.800 258.280 133.030 260.200 ;
        RECT 141.090 258.280 141.320 260.200 ;
        RECT 142.020 260.180 142.340 260.200 ;
        RECT 124.510 256.030 124.740 257.100 ;
        RECT 132.800 256.030 133.030 257.100 ;
        RECT 141.090 256.030 141.320 257.100 ;
        RECT 142.020 256.030 142.300 256.040 ;
        RECT 143.580 256.030 148.560 260.200 ;
        RECT 150.510 258.280 150.740 260.200 ;
        RECT 158.800 258.280 159.030 260.200 ;
        RECT 167.090 258.280 167.320 260.200 ;
        RECT 168.020 260.180 168.340 260.200 ;
        RECT 150.510 256.030 150.740 257.100 ;
        RECT 158.800 256.030 159.030 257.100 ;
        RECT 167.090 256.030 167.320 257.100 ;
        RECT 168.020 256.030 168.300 256.040 ;
        RECT 169.580 256.030 174.560 260.200 ;
        RECT 176.510 258.280 176.740 260.200 ;
        RECT 184.800 258.280 185.030 260.200 ;
        RECT 193.090 258.280 193.320 260.200 ;
        RECT 194.020 260.180 194.340 260.200 ;
        RECT 176.510 256.030 176.740 257.100 ;
        RECT 184.800 256.030 185.030 257.100 ;
        RECT 193.090 256.030 193.320 257.100 ;
        RECT 194.020 256.030 194.300 256.040 ;
        RECT 195.580 256.030 200.560 260.200 ;
        RECT 202.510 258.280 202.740 260.200 ;
        RECT 210.800 258.280 211.030 260.200 ;
        RECT 219.090 258.280 219.320 260.200 ;
        RECT 220.020 260.180 220.340 260.200 ;
        RECT 202.510 256.030 202.740 257.100 ;
        RECT 210.800 256.030 211.030 257.100 ;
        RECT 219.090 256.030 219.320 257.100 ;
        RECT 220.020 256.030 220.300 256.040 ;
        RECT 221.580 256.030 226.560 260.200 ;
        RECT 228.510 258.280 228.740 260.200 ;
        RECT 236.800 258.280 237.030 260.200 ;
        RECT 245.090 258.280 245.320 260.200 ;
        RECT 246.020 260.180 246.340 260.200 ;
        RECT 228.510 256.030 228.740 257.100 ;
        RECT 236.800 256.030 237.030 257.100 ;
        RECT 245.090 256.030 245.320 257.100 ;
        RECT 246.020 256.030 246.300 256.040 ;
        RECT 247.580 256.030 252.560 260.200 ;
        RECT 254.510 258.280 254.740 260.200 ;
        RECT 262.800 258.280 263.030 260.200 ;
        RECT 271.090 258.280 271.320 260.200 ;
        RECT 272.020 260.180 272.340 260.200 ;
        RECT 254.510 256.030 254.740 257.100 ;
        RECT 262.800 256.030 263.030 257.100 ;
        RECT 271.090 256.030 271.320 257.100 ;
        RECT 272.020 256.030 272.300 256.040 ;
        RECT 273.580 256.030 278.560 260.200 ;
        RECT 280.510 258.280 280.740 260.200 ;
        RECT 288.800 258.280 289.030 260.200 ;
        RECT 297.090 258.280 297.320 260.200 ;
        RECT 298.020 260.180 298.340 260.200 ;
        RECT 280.510 256.030 280.740 257.100 ;
        RECT 288.800 256.030 289.030 257.100 ;
        RECT 297.090 256.030 297.320 257.100 ;
        RECT 298.020 256.030 298.300 256.040 ;
        RECT 299.580 256.030 304.560 260.200 ;
        RECT 46.250 255.960 70.560 256.030 ;
        RECT 39.400 252.200 70.560 255.960 ;
        RECT 72.250 252.200 96.560 256.030 ;
        RECT 98.250 252.200 122.560 256.030 ;
        RECT 124.250 252.200 148.560 256.030 ;
        RECT 150.250 252.200 174.560 256.030 ;
        RECT 176.250 252.200 200.560 256.030 ;
        RECT 202.250 252.200 226.560 256.030 ;
        RECT 228.250 252.200 252.560 256.030 ;
        RECT 254.250 252.200 278.560 256.030 ;
        RECT 280.250 252.200 304.560 256.030 ;
        RECT 39.400 252.120 47.370 252.200 ;
        RECT 39.400 247.720 44.730 252.120 ;
        RECT 46.510 250.100 46.740 252.120 ;
        RECT 54.800 250.100 55.030 252.200 ;
        RECT 63.090 250.100 63.320 252.200 ;
        RECT 64.020 252.180 64.300 252.200 ;
        RECT 46.510 247.780 46.740 248.920 ;
        RECT 54.800 247.780 55.030 248.920 ;
        RECT 63.090 247.780 63.320 248.920 ;
        RECT 65.580 247.780 70.560 252.200 ;
        RECT 72.510 250.100 72.740 252.200 ;
        RECT 80.800 250.100 81.030 252.200 ;
        RECT 89.090 250.100 89.320 252.200 ;
        RECT 90.020 252.180 90.300 252.200 ;
        RECT 72.510 247.780 72.740 248.920 ;
        RECT 80.800 247.780 81.030 248.920 ;
        RECT 89.090 247.780 89.320 248.920 ;
        RECT 91.580 247.780 96.560 252.200 ;
        RECT 98.510 250.100 98.740 252.200 ;
        RECT 106.800 250.100 107.030 252.200 ;
        RECT 115.090 250.100 115.320 252.200 ;
        RECT 116.020 252.180 116.300 252.200 ;
        RECT 98.510 247.780 98.740 248.920 ;
        RECT 106.800 247.780 107.030 248.920 ;
        RECT 115.090 247.780 115.320 248.920 ;
        RECT 117.580 247.780 122.560 252.200 ;
        RECT 124.510 250.100 124.740 252.200 ;
        RECT 132.800 250.100 133.030 252.200 ;
        RECT 141.090 250.100 141.320 252.200 ;
        RECT 142.020 252.180 142.300 252.200 ;
        RECT 124.510 247.780 124.740 248.920 ;
        RECT 132.800 247.780 133.030 248.920 ;
        RECT 141.090 247.780 141.320 248.920 ;
        RECT 143.580 247.780 148.560 252.200 ;
        RECT 150.510 250.100 150.740 252.200 ;
        RECT 158.800 250.100 159.030 252.200 ;
        RECT 167.090 250.100 167.320 252.200 ;
        RECT 168.020 252.180 168.300 252.200 ;
        RECT 150.510 247.780 150.740 248.920 ;
        RECT 158.800 247.780 159.030 248.920 ;
        RECT 167.090 247.780 167.320 248.920 ;
        RECT 169.580 247.780 174.560 252.200 ;
        RECT 176.510 250.100 176.740 252.200 ;
        RECT 184.800 250.100 185.030 252.200 ;
        RECT 193.090 250.100 193.320 252.200 ;
        RECT 194.020 252.180 194.300 252.200 ;
        RECT 176.510 247.780 176.740 248.920 ;
        RECT 184.800 247.780 185.030 248.920 ;
        RECT 193.090 247.780 193.320 248.920 ;
        RECT 195.580 247.780 200.560 252.200 ;
        RECT 202.510 250.100 202.740 252.200 ;
        RECT 210.800 250.100 211.030 252.200 ;
        RECT 219.090 250.100 219.320 252.200 ;
        RECT 220.020 252.180 220.300 252.200 ;
        RECT 202.510 247.780 202.740 248.920 ;
        RECT 210.800 247.780 211.030 248.920 ;
        RECT 219.090 247.780 219.320 248.920 ;
        RECT 221.580 247.780 226.560 252.200 ;
        RECT 228.510 250.100 228.740 252.200 ;
        RECT 236.800 250.100 237.030 252.200 ;
        RECT 245.090 250.100 245.320 252.200 ;
        RECT 246.020 252.180 246.300 252.200 ;
        RECT 228.510 247.780 228.740 248.920 ;
        RECT 236.800 247.780 237.030 248.920 ;
        RECT 245.090 247.780 245.320 248.920 ;
        RECT 247.580 247.780 252.560 252.200 ;
        RECT 254.510 250.100 254.740 252.200 ;
        RECT 262.800 250.100 263.030 252.200 ;
        RECT 271.090 250.100 271.320 252.200 ;
        RECT 272.020 252.180 272.300 252.200 ;
        RECT 254.510 247.780 254.740 248.920 ;
        RECT 262.800 247.780 263.030 248.920 ;
        RECT 271.090 247.780 271.320 248.920 ;
        RECT 273.580 247.780 278.560 252.200 ;
        RECT 280.510 250.100 280.740 252.200 ;
        RECT 288.800 250.100 289.030 252.200 ;
        RECT 297.090 250.100 297.320 252.200 ;
        RECT 298.020 252.180 298.300 252.200 ;
        RECT 280.510 247.780 280.740 248.920 ;
        RECT 288.800 247.780 289.030 248.920 ;
        RECT 297.090 247.780 297.320 248.920 ;
        RECT 299.580 247.780 304.560 252.200 ;
        RECT 46.250 247.770 63.890 247.780 ;
        RECT 64.440 247.770 70.560 247.780 ;
        RECT 46.250 247.720 70.560 247.770 ;
        RECT 39.400 243.950 70.560 247.720 ;
        RECT 72.250 247.770 89.890 247.780 ;
        RECT 90.440 247.770 96.560 247.780 ;
        RECT 72.250 243.950 96.560 247.770 ;
        RECT 98.250 247.770 115.890 247.780 ;
        RECT 116.440 247.770 122.560 247.780 ;
        RECT 98.250 243.950 122.560 247.770 ;
        RECT 124.250 247.770 141.890 247.780 ;
        RECT 142.440 247.770 148.560 247.780 ;
        RECT 124.250 243.950 148.560 247.770 ;
        RECT 150.250 247.770 167.890 247.780 ;
        RECT 168.440 247.770 174.560 247.780 ;
        RECT 150.250 243.950 174.560 247.770 ;
        RECT 176.250 247.770 193.890 247.780 ;
        RECT 194.440 247.770 200.560 247.780 ;
        RECT 176.250 243.950 200.560 247.770 ;
        RECT 202.250 247.770 219.890 247.780 ;
        RECT 220.440 247.770 226.560 247.780 ;
        RECT 202.250 243.950 226.560 247.770 ;
        RECT 228.250 247.770 245.890 247.780 ;
        RECT 246.440 247.770 252.560 247.780 ;
        RECT 228.250 243.950 252.560 247.770 ;
        RECT 254.250 247.770 271.890 247.780 ;
        RECT 272.440 247.770 278.560 247.780 ;
        RECT 254.250 243.950 278.560 247.770 ;
        RECT 280.250 247.770 297.890 247.780 ;
        RECT 298.440 247.770 304.560 247.780 ;
        RECT 280.250 243.950 304.560 247.770 ;
        RECT 688.370 249.570 715.540 251.075 ;
        RECT 688.370 244.015 688.600 249.570 ;
        RECT 690.230 244.210 690.460 249.570 ;
        RECT 692.810 244.210 693.040 249.570 ;
        RECT 695.390 244.210 695.620 249.570 ;
        RECT 697.970 244.210 698.200 249.570 ;
        RECT 700.550 244.210 700.780 249.570 ;
        RECT 703.130 244.210 703.360 249.570 ;
        RECT 705.710 244.210 705.940 249.570 ;
        RECT 708.290 244.210 708.520 249.570 ;
        RECT 710.870 244.210 711.100 249.570 ;
        RECT 713.450 244.210 713.680 249.570 ;
        RECT 715.310 244.015 715.540 249.570 ;
        RECT 39.400 243.820 46.740 243.950 ;
        RECT 39.400 239.380 44.730 243.820 ;
        RECT 46.510 241.920 46.740 243.820 ;
        RECT 54.800 241.920 55.030 243.950 ;
        RECT 63.090 241.920 63.320 243.950 ;
        RECT 46.510 239.380 46.740 240.740 ;
        RECT 39.400 239.280 46.950 239.380 ;
        RECT 54.800 239.280 55.030 240.740 ;
        RECT 63.090 239.280 63.320 240.740 ;
        RECT 64.020 239.280 64.300 239.290 ;
        RECT 65.580 239.280 70.560 243.950 ;
        RECT 72.510 241.920 72.740 243.950 ;
        RECT 80.800 241.920 81.030 243.950 ;
        RECT 89.090 241.920 89.320 243.950 ;
        RECT 72.510 239.280 72.740 240.740 ;
        RECT 80.800 239.280 81.030 240.740 ;
        RECT 89.090 239.280 89.320 240.740 ;
        RECT 90.020 239.280 90.300 239.290 ;
        RECT 91.580 239.280 96.560 243.950 ;
        RECT 98.510 241.920 98.740 243.950 ;
        RECT 106.800 241.920 107.030 243.950 ;
        RECT 115.090 241.920 115.320 243.950 ;
        RECT 98.510 239.280 98.740 240.740 ;
        RECT 106.800 239.280 107.030 240.740 ;
        RECT 115.090 239.280 115.320 240.740 ;
        RECT 116.020 239.280 116.300 239.290 ;
        RECT 117.580 239.280 122.560 243.950 ;
        RECT 124.510 241.920 124.740 243.950 ;
        RECT 132.800 241.920 133.030 243.950 ;
        RECT 141.090 241.920 141.320 243.950 ;
        RECT 124.510 239.280 124.740 240.740 ;
        RECT 132.800 239.280 133.030 240.740 ;
        RECT 141.090 239.280 141.320 240.740 ;
        RECT 142.020 239.280 142.300 239.290 ;
        RECT 143.580 239.280 148.560 243.950 ;
        RECT 150.510 241.920 150.740 243.950 ;
        RECT 158.800 241.920 159.030 243.950 ;
        RECT 167.090 241.920 167.320 243.950 ;
        RECT 150.510 239.280 150.740 240.740 ;
        RECT 158.800 239.280 159.030 240.740 ;
        RECT 167.090 239.280 167.320 240.740 ;
        RECT 168.020 239.280 168.300 239.290 ;
        RECT 169.580 239.280 174.560 243.950 ;
        RECT 176.510 241.920 176.740 243.950 ;
        RECT 184.800 241.920 185.030 243.950 ;
        RECT 193.090 241.920 193.320 243.950 ;
        RECT 176.510 239.280 176.740 240.740 ;
        RECT 184.800 239.280 185.030 240.740 ;
        RECT 193.090 239.280 193.320 240.740 ;
        RECT 194.020 239.280 194.300 239.290 ;
        RECT 195.580 239.280 200.560 243.950 ;
        RECT 202.510 241.920 202.740 243.950 ;
        RECT 210.800 241.920 211.030 243.950 ;
        RECT 219.090 241.920 219.320 243.950 ;
        RECT 202.510 239.280 202.740 240.740 ;
        RECT 210.800 239.280 211.030 240.740 ;
        RECT 219.090 239.280 219.320 240.740 ;
        RECT 220.020 239.280 220.300 239.290 ;
        RECT 221.580 239.280 226.560 243.950 ;
        RECT 228.510 241.920 228.740 243.950 ;
        RECT 236.800 241.920 237.030 243.950 ;
        RECT 245.090 241.920 245.320 243.950 ;
        RECT 228.510 239.280 228.740 240.740 ;
        RECT 236.800 239.280 237.030 240.740 ;
        RECT 245.090 239.280 245.320 240.740 ;
        RECT 246.020 239.280 246.300 239.290 ;
        RECT 247.580 239.280 252.560 243.950 ;
        RECT 254.510 241.920 254.740 243.950 ;
        RECT 262.800 241.920 263.030 243.950 ;
        RECT 271.090 241.920 271.320 243.950 ;
        RECT 254.510 239.280 254.740 240.740 ;
        RECT 262.800 239.280 263.030 240.740 ;
        RECT 271.090 239.280 271.320 240.740 ;
        RECT 272.020 239.280 272.300 239.290 ;
        RECT 273.580 239.280 278.560 243.950 ;
        RECT 280.510 241.920 280.740 243.950 ;
        RECT 288.800 241.920 289.030 243.950 ;
        RECT 297.090 241.920 297.320 243.950 ;
        RECT 280.510 239.280 280.740 240.740 ;
        RECT 288.800 239.280 289.030 240.740 ;
        RECT 297.090 239.280 297.320 240.740 ;
        RECT 298.020 239.280 298.300 239.290 ;
        RECT 299.580 239.280 304.560 243.950 ;
        RECT 689.430 243.775 689.970 244.005 ;
        RECT 690.720 243.775 691.260 244.005 ;
        RECT 692.010 243.775 692.550 244.005 ;
        RECT 693.300 243.775 693.840 244.005 ;
        RECT 694.590 243.775 695.130 244.005 ;
        RECT 695.880 243.775 696.420 244.005 ;
        RECT 697.170 243.775 697.710 244.005 ;
        RECT 698.460 243.775 699.000 244.005 ;
        RECT 699.750 243.775 700.290 244.005 ;
        RECT 701.040 243.775 701.580 244.005 ;
        RECT 702.330 243.775 702.870 244.005 ;
        RECT 703.620 243.775 704.160 244.005 ;
        RECT 704.910 243.775 705.450 244.005 ;
        RECT 706.200 243.775 706.740 244.005 ;
        RECT 707.490 243.775 708.030 244.005 ;
        RECT 708.780 243.775 709.320 244.005 ;
        RECT 710.070 243.775 710.610 244.005 ;
        RECT 711.360 243.775 711.900 244.005 ;
        RECT 712.650 243.775 713.190 244.005 ;
        RECT 713.940 243.775 714.480 244.005 ;
        RECT 39.400 235.480 70.560 239.280 ;
        RECT 39.400 230.760 44.730 235.480 ;
        RECT 46.250 235.450 70.560 235.480 ;
        RECT 72.250 235.450 96.560 239.280 ;
        RECT 98.250 235.450 122.560 239.280 ;
        RECT 124.250 235.450 148.560 239.280 ;
        RECT 150.250 235.450 174.560 239.280 ;
        RECT 176.250 235.450 200.560 239.280 ;
        RECT 202.250 235.450 226.560 239.280 ;
        RECT 228.250 235.450 252.560 239.280 ;
        RECT 254.250 235.450 278.560 239.280 ;
        RECT 280.250 235.450 304.560 239.280 ;
        RECT 46.510 233.740 46.740 235.450 ;
        RECT 54.800 233.740 55.030 235.450 ;
        RECT 63.090 233.740 63.320 235.450 ;
        RECT 64.020 235.430 64.310 235.450 ;
        RECT 46.510 230.780 46.740 232.560 ;
        RECT 54.800 230.780 55.030 232.560 ;
        RECT 63.090 230.780 63.320 232.560 ;
        RECT 65.580 230.780 70.560 235.450 ;
        RECT 72.510 233.740 72.740 235.450 ;
        RECT 80.800 233.740 81.030 235.450 ;
        RECT 89.090 233.740 89.320 235.450 ;
        RECT 90.020 235.430 90.310 235.450 ;
        RECT 72.510 230.780 72.740 232.560 ;
        RECT 80.800 230.780 81.030 232.560 ;
        RECT 89.090 230.780 89.320 232.560 ;
        RECT 91.580 230.780 96.560 235.450 ;
        RECT 98.510 233.740 98.740 235.450 ;
        RECT 106.800 233.740 107.030 235.450 ;
        RECT 115.090 233.740 115.320 235.450 ;
        RECT 116.020 235.430 116.310 235.450 ;
        RECT 98.510 230.780 98.740 232.560 ;
        RECT 106.800 230.780 107.030 232.560 ;
        RECT 115.090 230.780 115.320 232.560 ;
        RECT 117.580 230.780 122.560 235.450 ;
        RECT 124.510 233.740 124.740 235.450 ;
        RECT 132.800 233.740 133.030 235.450 ;
        RECT 141.090 233.740 141.320 235.450 ;
        RECT 142.020 235.430 142.310 235.450 ;
        RECT 124.510 230.780 124.740 232.560 ;
        RECT 132.800 230.780 133.030 232.560 ;
        RECT 141.090 230.780 141.320 232.560 ;
        RECT 143.580 230.780 148.560 235.450 ;
        RECT 150.510 233.740 150.740 235.450 ;
        RECT 158.800 233.740 159.030 235.450 ;
        RECT 167.090 233.740 167.320 235.450 ;
        RECT 168.020 235.430 168.310 235.450 ;
        RECT 150.510 230.780 150.740 232.560 ;
        RECT 158.800 230.780 159.030 232.560 ;
        RECT 167.090 230.780 167.320 232.560 ;
        RECT 169.580 230.780 174.560 235.450 ;
        RECT 176.510 233.740 176.740 235.450 ;
        RECT 184.800 233.740 185.030 235.450 ;
        RECT 193.090 233.740 193.320 235.450 ;
        RECT 194.020 235.430 194.310 235.450 ;
        RECT 176.510 230.780 176.740 232.560 ;
        RECT 184.800 230.780 185.030 232.560 ;
        RECT 193.090 230.780 193.320 232.560 ;
        RECT 195.580 230.780 200.560 235.450 ;
        RECT 202.510 233.740 202.740 235.450 ;
        RECT 210.800 233.740 211.030 235.450 ;
        RECT 219.090 233.740 219.320 235.450 ;
        RECT 220.020 235.430 220.310 235.450 ;
        RECT 202.510 230.780 202.740 232.560 ;
        RECT 210.800 230.780 211.030 232.560 ;
        RECT 219.090 230.780 219.320 232.560 ;
        RECT 221.580 230.780 226.560 235.450 ;
        RECT 228.510 233.740 228.740 235.450 ;
        RECT 236.800 233.740 237.030 235.450 ;
        RECT 245.090 233.740 245.320 235.450 ;
        RECT 246.020 235.430 246.310 235.450 ;
        RECT 228.510 230.780 228.740 232.560 ;
        RECT 236.800 230.780 237.030 232.560 ;
        RECT 245.090 230.780 245.320 232.560 ;
        RECT 247.580 230.780 252.560 235.450 ;
        RECT 254.510 233.740 254.740 235.450 ;
        RECT 262.800 233.740 263.030 235.450 ;
        RECT 271.090 233.740 271.320 235.450 ;
        RECT 272.020 235.430 272.310 235.450 ;
        RECT 254.510 230.780 254.740 232.560 ;
        RECT 262.800 230.780 263.030 232.560 ;
        RECT 271.090 230.780 271.320 232.560 ;
        RECT 273.580 230.780 278.560 235.450 ;
        RECT 280.510 233.740 280.740 235.450 ;
        RECT 288.800 233.740 289.030 235.450 ;
        RECT 297.090 233.740 297.320 235.450 ;
        RECT 298.020 235.430 298.310 235.450 ;
        RECT 280.510 230.780 280.740 232.560 ;
        RECT 288.800 230.780 289.030 232.560 ;
        RECT 297.090 230.780 297.320 232.560 ;
        RECT 299.580 230.780 304.560 235.450 ;
        RECT 46.250 230.770 63.850 230.780 ;
        RECT 64.420 230.770 70.560 230.780 ;
        RECT 46.250 230.760 70.560 230.770 ;
        RECT 39.400 226.950 70.560 230.760 ;
        RECT 72.250 230.770 89.850 230.780 ;
        RECT 90.420 230.770 96.560 230.780 ;
        RECT 72.250 226.950 96.560 230.770 ;
        RECT 98.250 230.770 115.850 230.780 ;
        RECT 116.420 230.770 122.560 230.780 ;
        RECT 98.250 226.950 122.560 230.770 ;
        RECT 124.250 230.770 141.850 230.780 ;
        RECT 142.420 230.770 148.560 230.780 ;
        RECT 124.250 226.950 148.560 230.770 ;
        RECT 150.250 230.770 167.850 230.780 ;
        RECT 168.420 230.770 174.560 230.780 ;
        RECT 150.250 226.950 174.560 230.770 ;
        RECT 176.250 230.770 193.850 230.780 ;
        RECT 194.420 230.770 200.560 230.780 ;
        RECT 176.250 226.950 200.560 230.770 ;
        RECT 202.250 230.770 219.850 230.780 ;
        RECT 220.420 230.770 226.560 230.780 ;
        RECT 202.250 226.950 226.560 230.770 ;
        RECT 228.250 230.770 245.850 230.780 ;
        RECT 246.420 230.770 252.560 230.780 ;
        RECT 228.250 226.950 252.560 230.770 ;
        RECT 254.250 230.770 271.850 230.780 ;
        RECT 272.420 230.770 278.560 230.780 ;
        RECT 254.250 226.950 278.560 230.770 ;
        RECT 280.250 230.770 297.850 230.780 ;
        RECT 298.420 230.770 304.560 230.780 ;
        RECT 280.250 226.950 304.560 230.770 ;
        RECT 39.400 226.860 46.930 226.950 ;
        RECT 39.400 222.770 44.730 226.860 ;
        RECT 46.510 225.560 46.740 226.860 ;
        RECT 54.800 225.560 55.030 226.950 ;
        RECT 63.090 225.560 63.320 226.950 ;
        RECT 64.020 226.910 64.310 226.950 ;
        RECT 46.510 222.780 46.740 224.380 ;
        RECT 54.800 222.780 55.030 224.380 ;
        RECT 63.090 222.780 63.320 224.380 ;
        RECT 65.580 222.780 70.560 226.950 ;
        RECT 72.510 225.560 72.740 226.950 ;
        RECT 80.800 225.560 81.030 226.950 ;
        RECT 89.090 225.560 89.320 226.950 ;
        RECT 90.020 226.910 90.310 226.950 ;
        RECT 72.510 222.780 72.740 224.380 ;
        RECT 80.800 222.780 81.030 224.380 ;
        RECT 89.090 222.780 89.320 224.380 ;
        RECT 91.580 222.780 96.560 226.950 ;
        RECT 98.510 225.560 98.740 226.950 ;
        RECT 106.800 225.560 107.030 226.950 ;
        RECT 115.090 225.560 115.320 226.950 ;
        RECT 116.020 226.910 116.310 226.950 ;
        RECT 98.510 222.780 98.740 224.380 ;
        RECT 106.800 222.780 107.030 224.380 ;
        RECT 115.090 222.780 115.320 224.380 ;
        RECT 117.580 222.780 122.560 226.950 ;
        RECT 124.510 225.560 124.740 226.950 ;
        RECT 132.800 225.560 133.030 226.950 ;
        RECT 141.090 225.560 141.320 226.950 ;
        RECT 142.020 226.910 142.310 226.950 ;
        RECT 124.510 222.780 124.740 224.380 ;
        RECT 132.800 222.780 133.030 224.380 ;
        RECT 141.090 222.780 141.320 224.380 ;
        RECT 143.580 222.780 148.560 226.950 ;
        RECT 150.510 225.560 150.740 226.950 ;
        RECT 158.800 225.560 159.030 226.950 ;
        RECT 167.090 225.560 167.320 226.950 ;
        RECT 168.020 226.910 168.310 226.950 ;
        RECT 150.510 222.780 150.740 224.380 ;
        RECT 158.800 222.780 159.030 224.380 ;
        RECT 167.090 222.780 167.320 224.380 ;
        RECT 169.580 222.780 174.560 226.950 ;
        RECT 176.510 225.560 176.740 226.950 ;
        RECT 184.800 225.560 185.030 226.950 ;
        RECT 193.090 225.560 193.320 226.950 ;
        RECT 194.020 226.910 194.310 226.950 ;
        RECT 176.510 222.780 176.740 224.380 ;
        RECT 184.800 222.780 185.030 224.380 ;
        RECT 193.090 222.780 193.320 224.380 ;
        RECT 195.580 222.780 200.560 226.950 ;
        RECT 202.510 225.560 202.740 226.950 ;
        RECT 210.800 225.560 211.030 226.950 ;
        RECT 219.090 225.560 219.320 226.950 ;
        RECT 220.020 226.910 220.310 226.950 ;
        RECT 202.510 222.780 202.740 224.380 ;
        RECT 210.800 222.780 211.030 224.380 ;
        RECT 219.090 222.780 219.320 224.380 ;
        RECT 221.580 222.780 226.560 226.950 ;
        RECT 228.510 225.560 228.740 226.950 ;
        RECT 236.800 225.560 237.030 226.950 ;
        RECT 245.090 225.560 245.320 226.950 ;
        RECT 246.020 226.910 246.310 226.950 ;
        RECT 228.510 222.780 228.740 224.380 ;
        RECT 236.800 222.780 237.030 224.380 ;
        RECT 245.090 222.780 245.320 224.380 ;
        RECT 247.580 222.780 252.560 226.950 ;
        RECT 254.510 225.560 254.740 226.950 ;
        RECT 262.800 225.560 263.030 226.950 ;
        RECT 271.090 225.560 271.320 226.950 ;
        RECT 272.020 226.910 272.310 226.950 ;
        RECT 254.510 222.780 254.740 224.380 ;
        RECT 262.800 222.780 263.030 224.380 ;
        RECT 271.090 222.780 271.320 224.380 ;
        RECT 273.580 222.780 278.560 226.950 ;
        RECT 280.510 225.560 280.740 226.950 ;
        RECT 288.800 225.560 289.030 226.950 ;
        RECT 297.090 225.560 297.320 226.950 ;
        RECT 298.020 226.910 298.310 226.950 ;
        RECT 280.510 222.780 280.740 224.380 ;
        RECT 288.800 222.780 289.030 224.380 ;
        RECT 297.090 222.780 297.320 224.380 ;
        RECT 299.580 222.780 304.560 226.950 ;
        RECT 46.250 222.770 63.850 222.780 ;
        RECT 64.560 222.770 70.560 222.780 ;
        RECT 39.400 218.950 70.560 222.770 ;
        RECT 72.250 222.770 89.850 222.780 ;
        RECT 90.560 222.770 96.560 222.780 ;
        RECT 72.250 218.950 96.560 222.770 ;
        RECT 98.250 222.770 115.850 222.780 ;
        RECT 116.560 222.770 122.560 222.780 ;
        RECT 98.250 218.950 122.560 222.770 ;
        RECT 124.250 222.770 141.850 222.780 ;
        RECT 142.560 222.770 148.560 222.780 ;
        RECT 124.250 218.950 148.560 222.770 ;
        RECT 150.250 222.770 167.850 222.780 ;
        RECT 168.560 222.770 174.560 222.780 ;
        RECT 150.250 218.950 174.560 222.770 ;
        RECT 176.250 222.770 193.850 222.780 ;
        RECT 194.560 222.770 200.560 222.780 ;
        RECT 176.250 218.950 200.560 222.770 ;
        RECT 202.250 222.770 219.850 222.780 ;
        RECT 220.560 222.770 226.560 222.780 ;
        RECT 202.250 218.950 226.560 222.770 ;
        RECT 228.250 222.770 245.850 222.780 ;
        RECT 246.560 222.770 252.560 222.780 ;
        RECT 228.250 218.950 252.560 222.770 ;
        RECT 254.250 222.770 271.850 222.780 ;
        RECT 272.560 222.770 278.560 222.780 ;
        RECT 254.250 218.950 278.560 222.770 ;
        RECT 280.250 222.770 297.850 222.780 ;
        RECT 298.560 222.770 304.560 222.780 ;
        RECT 280.250 218.950 304.560 222.770 ;
        RECT 39.400 218.870 46.740 218.950 ;
        RECT 39.400 214.820 44.730 218.870 ;
        RECT 46.510 217.380 46.740 218.870 ;
        RECT 54.800 217.380 55.030 218.950 ;
        RECT 63.090 217.380 63.320 218.950 ;
        RECT 64.020 218.910 64.310 218.950 ;
        RECT 46.510 214.820 46.740 216.200 ;
        RECT 39.400 214.780 46.750 214.820 ;
        RECT 54.800 214.780 55.030 216.200 ;
        RECT 63.090 214.780 63.320 216.200 ;
        RECT 64.020 214.780 64.300 214.810 ;
        RECT 65.580 214.780 70.560 218.950 ;
        RECT 72.510 217.380 72.740 218.950 ;
        RECT 80.800 217.380 81.030 218.950 ;
        RECT 89.090 217.380 89.320 218.950 ;
        RECT 90.020 218.910 90.310 218.950 ;
        RECT 72.510 214.780 72.740 216.200 ;
        RECT 80.800 214.780 81.030 216.200 ;
        RECT 89.090 214.780 89.320 216.200 ;
        RECT 90.020 214.780 90.300 214.810 ;
        RECT 91.580 214.780 96.560 218.950 ;
        RECT 98.510 217.380 98.740 218.950 ;
        RECT 106.800 217.380 107.030 218.950 ;
        RECT 115.090 217.380 115.320 218.950 ;
        RECT 116.020 218.910 116.310 218.950 ;
        RECT 98.510 214.780 98.740 216.200 ;
        RECT 106.800 214.780 107.030 216.200 ;
        RECT 115.090 214.780 115.320 216.200 ;
        RECT 116.020 214.780 116.300 214.810 ;
        RECT 117.580 214.780 122.560 218.950 ;
        RECT 124.510 217.380 124.740 218.950 ;
        RECT 132.800 217.380 133.030 218.950 ;
        RECT 141.090 217.380 141.320 218.950 ;
        RECT 142.020 218.910 142.310 218.950 ;
        RECT 124.510 214.780 124.740 216.200 ;
        RECT 132.800 214.780 133.030 216.200 ;
        RECT 141.090 214.780 141.320 216.200 ;
        RECT 142.020 214.780 142.300 214.810 ;
        RECT 143.580 214.780 148.560 218.950 ;
        RECT 150.510 217.380 150.740 218.950 ;
        RECT 158.800 217.380 159.030 218.950 ;
        RECT 167.090 217.380 167.320 218.950 ;
        RECT 168.020 218.910 168.310 218.950 ;
        RECT 150.510 214.780 150.740 216.200 ;
        RECT 158.800 214.780 159.030 216.200 ;
        RECT 167.090 214.780 167.320 216.200 ;
        RECT 168.020 214.780 168.300 214.810 ;
        RECT 169.580 214.780 174.560 218.950 ;
        RECT 176.510 217.380 176.740 218.950 ;
        RECT 184.800 217.380 185.030 218.950 ;
        RECT 193.090 217.380 193.320 218.950 ;
        RECT 194.020 218.910 194.310 218.950 ;
        RECT 176.510 214.780 176.740 216.200 ;
        RECT 184.800 214.780 185.030 216.200 ;
        RECT 193.090 214.780 193.320 216.200 ;
        RECT 194.020 214.780 194.300 214.810 ;
        RECT 195.580 214.780 200.560 218.950 ;
        RECT 202.510 217.380 202.740 218.950 ;
        RECT 210.800 217.380 211.030 218.950 ;
        RECT 219.090 217.380 219.320 218.950 ;
        RECT 220.020 218.910 220.310 218.950 ;
        RECT 202.510 214.780 202.740 216.200 ;
        RECT 210.800 214.780 211.030 216.200 ;
        RECT 219.090 214.780 219.320 216.200 ;
        RECT 220.020 214.780 220.300 214.810 ;
        RECT 221.580 214.780 226.560 218.950 ;
        RECT 228.510 217.380 228.740 218.950 ;
        RECT 236.800 217.380 237.030 218.950 ;
        RECT 245.090 217.380 245.320 218.950 ;
        RECT 246.020 218.910 246.310 218.950 ;
        RECT 228.510 214.780 228.740 216.200 ;
        RECT 236.800 214.780 237.030 216.200 ;
        RECT 245.090 214.780 245.320 216.200 ;
        RECT 246.020 214.780 246.300 214.810 ;
        RECT 247.580 214.780 252.560 218.950 ;
        RECT 254.510 217.380 254.740 218.950 ;
        RECT 262.800 217.380 263.030 218.950 ;
        RECT 271.090 217.380 271.320 218.950 ;
        RECT 272.020 218.910 272.310 218.950 ;
        RECT 254.510 214.780 254.740 216.200 ;
        RECT 262.800 214.780 263.030 216.200 ;
        RECT 271.090 214.780 271.320 216.200 ;
        RECT 272.020 214.780 272.300 214.810 ;
        RECT 273.580 214.780 278.560 218.950 ;
        RECT 280.510 217.380 280.740 218.950 ;
        RECT 288.800 217.380 289.030 218.950 ;
        RECT 297.090 217.380 297.320 218.950 ;
        RECT 298.020 218.910 298.310 218.950 ;
        RECT 280.510 214.780 280.740 216.200 ;
        RECT 288.800 214.780 289.030 216.200 ;
        RECT 297.090 214.780 297.320 216.200 ;
        RECT 298.020 214.780 298.300 214.810 ;
        RECT 299.580 214.780 304.560 218.950 ;
        RECT 39.400 210.950 70.560 214.780 ;
        RECT 72.250 210.950 96.560 214.780 ;
        RECT 98.250 210.950 122.560 214.780 ;
        RECT 124.250 210.950 148.560 214.780 ;
        RECT 150.250 210.950 174.560 214.780 ;
        RECT 176.250 210.950 200.560 214.780 ;
        RECT 202.250 210.950 226.560 214.780 ;
        RECT 228.250 210.950 252.560 214.780 ;
        RECT 254.250 210.950 278.560 214.780 ;
        RECT 280.250 210.950 304.560 214.780 ;
        RECT 39.400 210.920 46.750 210.950 ;
        RECT 39.400 206.880 44.730 210.920 ;
        RECT 46.510 209.200 46.740 210.920 ;
        RECT 54.800 209.200 55.030 210.950 ;
        RECT 63.090 209.200 63.320 210.950 ;
        RECT 64.020 210.940 64.310 210.950 ;
        RECT 46.510 206.880 46.740 208.020 ;
        RECT 39.400 206.780 46.740 206.880 ;
        RECT 54.800 206.780 55.030 208.020 ;
        RECT 63.090 206.780 63.320 208.020 ;
        RECT 65.580 206.780 70.560 210.950 ;
        RECT 72.510 209.200 72.740 210.950 ;
        RECT 80.800 209.200 81.030 210.950 ;
        RECT 89.090 209.200 89.320 210.950 ;
        RECT 90.020 210.940 90.310 210.950 ;
        RECT 72.510 206.780 72.740 208.020 ;
        RECT 80.800 206.780 81.030 208.020 ;
        RECT 89.090 206.780 89.320 208.020 ;
        RECT 91.580 206.780 96.560 210.950 ;
        RECT 98.510 209.200 98.740 210.950 ;
        RECT 106.800 209.200 107.030 210.950 ;
        RECT 115.090 209.200 115.320 210.950 ;
        RECT 116.020 210.940 116.310 210.950 ;
        RECT 98.510 206.780 98.740 208.020 ;
        RECT 106.800 206.780 107.030 208.020 ;
        RECT 115.090 206.780 115.320 208.020 ;
        RECT 117.580 206.780 122.560 210.950 ;
        RECT 124.510 209.200 124.740 210.950 ;
        RECT 132.800 209.200 133.030 210.950 ;
        RECT 141.090 209.200 141.320 210.950 ;
        RECT 142.020 210.940 142.310 210.950 ;
        RECT 124.510 206.780 124.740 208.020 ;
        RECT 132.800 206.780 133.030 208.020 ;
        RECT 141.090 206.780 141.320 208.020 ;
        RECT 143.580 206.780 148.560 210.950 ;
        RECT 150.510 209.200 150.740 210.950 ;
        RECT 158.800 209.200 159.030 210.950 ;
        RECT 167.090 209.200 167.320 210.950 ;
        RECT 168.020 210.940 168.310 210.950 ;
        RECT 150.510 206.780 150.740 208.020 ;
        RECT 158.800 206.780 159.030 208.020 ;
        RECT 167.090 206.780 167.320 208.020 ;
        RECT 169.580 206.780 174.560 210.950 ;
        RECT 176.510 209.200 176.740 210.950 ;
        RECT 184.800 209.200 185.030 210.950 ;
        RECT 193.090 209.200 193.320 210.950 ;
        RECT 194.020 210.940 194.310 210.950 ;
        RECT 176.510 206.780 176.740 208.020 ;
        RECT 184.800 206.780 185.030 208.020 ;
        RECT 193.090 206.780 193.320 208.020 ;
        RECT 195.580 206.780 200.560 210.950 ;
        RECT 202.510 209.200 202.740 210.950 ;
        RECT 210.800 209.200 211.030 210.950 ;
        RECT 219.090 209.200 219.320 210.950 ;
        RECT 220.020 210.940 220.310 210.950 ;
        RECT 202.510 206.780 202.740 208.020 ;
        RECT 210.800 206.780 211.030 208.020 ;
        RECT 219.090 206.780 219.320 208.020 ;
        RECT 221.580 206.780 226.560 210.950 ;
        RECT 228.510 209.200 228.740 210.950 ;
        RECT 236.800 209.200 237.030 210.950 ;
        RECT 245.090 209.200 245.320 210.950 ;
        RECT 246.020 210.940 246.310 210.950 ;
        RECT 228.510 206.780 228.740 208.020 ;
        RECT 236.800 206.780 237.030 208.020 ;
        RECT 245.090 206.780 245.320 208.020 ;
        RECT 247.580 206.780 252.560 210.950 ;
        RECT 254.510 209.200 254.740 210.950 ;
        RECT 262.800 209.200 263.030 210.950 ;
        RECT 271.090 209.200 271.320 210.950 ;
        RECT 272.020 210.940 272.310 210.950 ;
        RECT 254.510 206.780 254.740 208.020 ;
        RECT 262.800 206.780 263.030 208.020 ;
        RECT 271.090 206.780 271.320 208.020 ;
        RECT 273.580 206.780 278.560 210.950 ;
        RECT 280.510 209.200 280.740 210.950 ;
        RECT 288.800 209.200 289.030 210.950 ;
        RECT 297.090 209.200 297.320 210.950 ;
        RECT 298.020 210.940 298.310 210.950 ;
        RECT 280.510 206.780 280.740 208.020 ;
        RECT 288.800 206.780 289.030 208.020 ;
        RECT 297.090 206.780 297.320 208.020 ;
        RECT 299.580 206.780 304.560 210.950 ;
        RECT 39.400 206.760 63.910 206.780 ;
        RECT 64.460 206.760 70.560 206.780 ;
        RECT 39.400 202.980 70.560 206.760 ;
        RECT 39.400 198.510 44.730 202.980 ;
        RECT 46.250 202.950 70.560 202.980 ;
        RECT 72.250 206.760 89.910 206.780 ;
        RECT 90.460 206.760 96.560 206.780 ;
        RECT 72.250 202.950 96.560 206.760 ;
        RECT 98.250 206.760 115.910 206.780 ;
        RECT 116.460 206.760 122.560 206.780 ;
        RECT 98.250 202.950 122.560 206.760 ;
        RECT 124.250 206.760 141.910 206.780 ;
        RECT 142.460 206.760 148.560 206.780 ;
        RECT 124.250 202.950 148.560 206.760 ;
        RECT 150.250 206.760 167.910 206.780 ;
        RECT 168.460 206.760 174.560 206.780 ;
        RECT 150.250 202.950 174.560 206.760 ;
        RECT 176.250 206.760 193.910 206.780 ;
        RECT 194.460 206.760 200.560 206.780 ;
        RECT 176.250 202.950 200.560 206.760 ;
        RECT 202.250 206.760 219.910 206.780 ;
        RECT 220.460 206.760 226.560 206.780 ;
        RECT 202.250 202.950 226.560 206.760 ;
        RECT 228.250 206.760 245.910 206.780 ;
        RECT 246.460 206.760 252.560 206.780 ;
        RECT 228.250 202.950 252.560 206.760 ;
        RECT 254.250 206.760 271.910 206.780 ;
        RECT 272.460 206.760 278.560 206.780 ;
        RECT 254.250 202.950 278.560 206.760 ;
        RECT 280.250 206.760 297.910 206.780 ;
        RECT 298.460 206.760 304.560 206.780 ;
        RECT 280.250 202.950 304.560 206.760 ;
        RECT 46.510 201.020 46.740 202.950 ;
        RECT 54.800 201.020 55.030 202.950 ;
        RECT 63.090 201.020 63.320 202.950 ;
        RECT 64.020 202.920 64.310 202.950 ;
        RECT 46.510 198.510 46.740 199.840 ;
        RECT 39.400 198.280 47.300 198.510 ;
        RECT 54.800 198.280 55.030 199.840 ;
        RECT 63.090 198.280 63.320 199.840 ;
        RECT 65.580 198.280 70.560 202.950 ;
        RECT 72.510 201.020 72.740 202.950 ;
        RECT 80.800 201.020 81.030 202.950 ;
        RECT 89.090 201.020 89.320 202.950 ;
        RECT 90.020 202.920 90.310 202.950 ;
        RECT 72.510 198.280 72.740 199.840 ;
        RECT 80.800 198.280 81.030 199.840 ;
        RECT 89.090 198.280 89.320 199.840 ;
        RECT 91.580 198.280 96.560 202.950 ;
        RECT 98.510 201.020 98.740 202.950 ;
        RECT 106.800 201.020 107.030 202.950 ;
        RECT 115.090 201.020 115.320 202.950 ;
        RECT 116.020 202.920 116.310 202.950 ;
        RECT 98.510 198.280 98.740 199.840 ;
        RECT 106.800 198.280 107.030 199.840 ;
        RECT 115.090 198.280 115.320 199.840 ;
        RECT 117.580 198.280 122.560 202.950 ;
        RECT 124.510 201.020 124.740 202.950 ;
        RECT 132.800 201.020 133.030 202.950 ;
        RECT 141.090 201.020 141.320 202.950 ;
        RECT 142.020 202.920 142.310 202.950 ;
        RECT 124.510 198.280 124.740 199.840 ;
        RECT 132.800 198.280 133.030 199.840 ;
        RECT 141.090 198.280 141.320 199.840 ;
        RECT 143.580 198.280 148.560 202.950 ;
        RECT 150.510 201.020 150.740 202.950 ;
        RECT 158.800 201.020 159.030 202.950 ;
        RECT 167.090 201.020 167.320 202.950 ;
        RECT 168.020 202.920 168.310 202.950 ;
        RECT 150.510 198.280 150.740 199.840 ;
        RECT 158.800 198.280 159.030 199.840 ;
        RECT 167.090 198.280 167.320 199.840 ;
        RECT 169.580 198.280 174.560 202.950 ;
        RECT 176.510 201.020 176.740 202.950 ;
        RECT 184.800 201.020 185.030 202.950 ;
        RECT 193.090 201.020 193.320 202.950 ;
        RECT 194.020 202.920 194.310 202.950 ;
        RECT 176.510 198.280 176.740 199.840 ;
        RECT 184.800 198.280 185.030 199.840 ;
        RECT 193.090 198.280 193.320 199.840 ;
        RECT 195.580 198.280 200.560 202.950 ;
        RECT 202.510 201.020 202.740 202.950 ;
        RECT 210.800 201.020 211.030 202.950 ;
        RECT 219.090 201.020 219.320 202.950 ;
        RECT 220.020 202.920 220.310 202.950 ;
        RECT 202.510 198.280 202.740 199.840 ;
        RECT 210.800 198.280 211.030 199.840 ;
        RECT 219.090 198.280 219.320 199.840 ;
        RECT 221.580 198.280 226.560 202.950 ;
        RECT 228.510 201.020 228.740 202.950 ;
        RECT 236.800 201.020 237.030 202.950 ;
        RECT 245.090 201.020 245.320 202.950 ;
        RECT 246.020 202.920 246.310 202.950 ;
        RECT 228.510 198.280 228.740 199.840 ;
        RECT 236.800 198.280 237.030 199.840 ;
        RECT 245.090 198.280 245.320 199.840 ;
        RECT 247.580 198.280 252.560 202.950 ;
        RECT 254.510 201.020 254.740 202.950 ;
        RECT 262.800 201.020 263.030 202.950 ;
        RECT 271.090 201.020 271.320 202.950 ;
        RECT 272.020 202.920 272.310 202.950 ;
        RECT 254.510 198.280 254.740 199.840 ;
        RECT 262.800 198.280 263.030 199.840 ;
        RECT 271.090 198.280 271.320 199.840 ;
        RECT 273.580 198.280 278.560 202.950 ;
        RECT 280.510 201.020 280.740 202.950 ;
        RECT 288.800 201.020 289.030 202.950 ;
        RECT 297.090 201.020 297.320 202.950 ;
        RECT 298.020 202.920 298.310 202.950 ;
        RECT 280.510 198.280 280.740 199.840 ;
        RECT 288.800 198.280 289.030 199.840 ;
        RECT 297.090 198.280 297.320 199.840 ;
        RECT 299.580 198.280 304.560 202.950 ;
        RECT 39.400 198.250 63.890 198.280 ;
        RECT 64.380 198.250 70.560 198.280 ;
        RECT 39.400 194.610 70.560 198.250 ;
        RECT 39.400 189.870 44.730 194.610 ;
        RECT 46.250 194.450 70.560 194.610 ;
        RECT 72.250 198.250 89.890 198.280 ;
        RECT 90.380 198.250 96.560 198.280 ;
        RECT 72.250 194.450 96.560 198.250 ;
        RECT 98.250 198.250 115.890 198.280 ;
        RECT 116.380 198.250 122.560 198.280 ;
        RECT 98.250 194.450 122.560 198.250 ;
        RECT 124.250 198.250 141.890 198.280 ;
        RECT 142.380 198.250 148.560 198.280 ;
        RECT 124.250 194.450 148.560 198.250 ;
        RECT 150.250 198.250 167.890 198.280 ;
        RECT 168.380 198.250 174.560 198.280 ;
        RECT 150.250 194.450 174.560 198.250 ;
        RECT 176.250 198.250 193.890 198.280 ;
        RECT 194.380 198.250 200.560 198.280 ;
        RECT 176.250 194.450 200.560 198.250 ;
        RECT 202.250 198.250 219.890 198.280 ;
        RECT 220.380 198.250 226.560 198.280 ;
        RECT 202.250 194.450 226.560 198.250 ;
        RECT 228.250 198.250 245.890 198.280 ;
        RECT 246.380 198.250 252.560 198.280 ;
        RECT 228.250 194.450 252.560 198.250 ;
        RECT 254.250 198.250 271.890 198.280 ;
        RECT 272.380 198.250 278.560 198.280 ;
        RECT 254.250 194.450 278.560 198.250 ;
        RECT 280.250 198.250 297.890 198.280 ;
        RECT 298.380 198.250 304.560 198.280 ;
        RECT 280.250 194.450 304.560 198.250 ;
        RECT 46.510 192.840 46.740 194.450 ;
        RECT 54.800 192.840 55.030 194.450 ;
        RECT 63.090 192.840 63.320 194.450 ;
        RECT 64.020 194.440 64.310 194.450 ;
        RECT 46.510 189.870 46.740 191.660 ;
        RECT 39.400 189.780 46.780 189.870 ;
        RECT 54.800 189.780 55.030 191.660 ;
        RECT 63.090 189.780 63.320 191.660 ;
        RECT 65.580 189.780 70.560 194.450 ;
        RECT 72.510 192.840 72.740 194.450 ;
        RECT 80.800 192.840 81.030 194.450 ;
        RECT 89.090 192.840 89.320 194.450 ;
        RECT 90.020 194.440 90.310 194.450 ;
        RECT 72.510 189.780 72.740 191.660 ;
        RECT 80.800 189.780 81.030 191.660 ;
        RECT 89.090 189.780 89.320 191.660 ;
        RECT 91.580 189.780 96.560 194.450 ;
        RECT 98.510 192.840 98.740 194.450 ;
        RECT 106.800 192.840 107.030 194.450 ;
        RECT 115.090 192.840 115.320 194.450 ;
        RECT 116.020 194.440 116.310 194.450 ;
        RECT 98.510 189.780 98.740 191.660 ;
        RECT 106.800 189.780 107.030 191.660 ;
        RECT 115.090 189.780 115.320 191.660 ;
        RECT 117.580 189.780 122.560 194.450 ;
        RECT 124.510 192.840 124.740 194.450 ;
        RECT 132.800 192.840 133.030 194.450 ;
        RECT 141.090 192.840 141.320 194.450 ;
        RECT 142.020 194.440 142.310 194.450 ;
        RECT 124.510 189.780 124.740 191.660 ;
        RECT 132.800 189.780 133.030 191.660 ;
        RECT 141.090 189.780 141.320 191.660 ;
        RECT 143.580 189.780 148.560 194.450 ;
        RECT 150.510 192.840 150.740 194.450 ;
        RECT 158.800 192.840 159.030 194.450 ;
        RECT 167.090 192.840 167.320 194.450 ;
        RECT 168.020 194.440 168.310 194.450 ;
        RECT 150.510 189.780 150.740 191.660 ;
        RECT 158.800 189.780 159.030 191.660 ;
        RECT 167.090 189.780 167.320 191.660 ;
        RECT 169.580 189.780 174.560 194.450 ;
        RECT 176.510 192.840 176.740 194.450 ;
        RECT 184.800 192.840 185.030 194.450 ;
        RECT 193.090 192.840 193.320 194.450 ;
        RECT 194.020 194.440 194.310 194.450 ;
        RECT 176.510 189.780 176.740 191.660 ;
        RECT 184.800 189.780 185.030 191.660 ;
        RECT 193.090 189.780 193.320 191.660 ;
        RECT 195.580 189.780 200.560 194.450 ;
        RECT 202.510 192.840 202.740 194.450 ;
        RECT 210.800 192.840 211.030 194.450 ;
        RECT 219.090 192.840 219.320 194.450 ;
        RECT 220.020 194.440 220.310 194.450 ;
        RECT 202.510 189.780 202.740 191.660 ;
        RECT 210.800 189.780 211.030 191.660 ;
        RECT 219.090 189.780 219.320 191.660 ;
        RECT 221.580 189.780 226.560 194.450 ;
        RECT 228.510 192.840 228.740 194.450 ;
        RECT 236.800 192.840 237.030 194.450 ;
        RECT 245.090 192.840 245.320 194.450 ;
        RECT 246.020 194.440 246.310 194.450 ;
        RECT 228.510 189.780 228.740 191.660 ;
        RECT 236.800 189.780 237.030 191.660 ;
        RECT 245.090 189.780 245.320 191.660 ;
        RECT 247.580 189.780 252.560 194.450 ;
        RECT 254.510 192.840 254.740 194.450 ;
        RECT 262.800 192.840 263.030 194.450 ;
        RECT 271.090 192.840 271.320 194.450 ;
        RECT 272.020 194.440 272.310 194.450 ;
        RECT 254.510 189.780 254.740 191.660 ;
        RECT 262.800 189.780 263.030 191.660 ;
        RECT 271.090 189.780 271.320 191.660 ;
        RECT 273.580 189.780 278.560 194.450 ;
        RECT 280.510 192.840 280.740 194.450 ;
        RECT 288.800 192.840 289.030 194.450 ;
        RECT 297.090 192.840 297.320 194.450 ;
        RECT 298.020 194.440 298.310 194.450 ;
        RECT 280.510 189.780 280.740 191.660 ;
        RECT 288.800 189.780 289.030 191.660 ;
        RECT 297.090 189.780 297.320 191.660 ;
        RECT 299.580 189.780 304.560 194.450 ;
        RECT 39.400 189.770 63.910 189.780 ;
        RECT 64.400 189.770 70.560 189.780 ;
        RECT 39.400 185.970 70.560 189.770 ;
        RECT 39.400 181.800 44.730 185.970 ;
        RECT 46.250 185.950 70.560 185.970 ;
        RECT 72.250 189.770 89.910 189.780 ;
        RECT 90.400 189.770 96.560 189.780 ;
        RECT 72.250 185.950 96.560 189.770 ;
        RECT 98.250 189.770 115.910 189.780 ;
        RECT 116.400 189.770 122.560 189.780 ;
        RECT 98.250 185.950 122.560 189.770 ;
        RECT 124.250 189.770 141.910 189.780 ;
        RECT 142.400 189.770 148.560 189.780 ;
        RECT 124.250 185.950 148.560 189.770 ;
        RECT 150.250 189.770 167.910 189.780 ;
        RECT 168.400 189.770 174.560 189.780 ;
        RECT 150.250 185.950 174.560 189.770 ;
        RECT 176.250 189.770 193.910 189.780 ;
        RECT 194.400 189.770 200.560 189.780 ;
        RECT 176.250 185.950 200.560 189.770 ;
        RECT 202.250 189.770 219.910 189.780 ;
        RECT 220.400 189.770 226.560 189.780 ;
        RECT 202.250 185.950 226.560 189.770 ;
        RECT 228.250 189.770 245.910 189.780 ;
        RECT 246.400 189.770 252.560 189.780 ;
        RECT 228.250 185.950 252.560 189.770 ;
        RECT 254.250 189.770 271.910 189.780 ;
        RECT 272.400 189.770 278.560 189.780 ;
        RECT 254.250 185.950 278.560 189.770 ;
        RECT 280.250 189.770 297.910 189.780 ;
        RECT 298.400 189.770 304.560 189.780 ;
        RECT 280.250 185.950 304.560 189.770 ;
        RECT 46.510 184.660 46.740 185.950 ;
        RECT 54.800 184.660 55.030 185.950 ;
        RECT 63.090 184.660 63.320 185.950 ;
        RECT 64.020 185.910 64.310 185.950 ;
        RECT 46.510 182.200 46.740 183.480 ;
        RECT 45.980 181.800 48.010 182.200 ;
        RECT 39.400 181.780 48.010 181.800 ;
        RECT 54.800 181.780 55.030 183.480 ;
        RECT 63.090 181.780 63.320 183.480 ;
        RECT 65.580 181.780 70.560 185.950 ;
        RECT 72.510 184.660 72.740 185.950 ;
        RECT 80.800 184.660 81.030 185.950 ;
        RECT 89.090 184.660 89.320 185.950 ;
        RECT 90.020 185.910 90.310 185.950 ;
        RECT 72.510 181.780 72.740 183.480 ;
        RECT 80.800 181.780 81.030 183.480 ;
        RECT 89.090 181.780 89.320 183.480 ;
        RECT 91.580 181.780 96.560 185.950 ;
        RECT 98.510 184.660 98.740 185.950 ;
        RECT 106.800 184.660 107.030 185.950 ;
        RECT 115.090 184.660 115.320 185.950 ;
        RECT 116.020 185.910 116.310 185.950 ;
        RECT 98.510 181.780 98.740 183.480 ;
        RECT 106.800 181.780 107.030 183.480 ;
        RECT 115.090 181.780 115.320 183.480 ;
        RECT 117.580 181.780 122.560 185.950 ;
        RECT 124.510 184.660 124.740 185.950 ;
        RECT 132.800 184.660 133.030 185.950 ;
        RECT 141.090 184.660 141.320 185.950 ;
        RECT 142.020 185.910 142.310 185.950 ;
        RECT 124.510 181.780 124.740 183.480 ;
        RECT 132.800 181.780 133.030 183.480 ;
        RECT 141.090 181.780 141.320 183.480 ;
        RECT 143.580 181.780 148.560 185.950 ;
        RECT 150.510 184.660 150.740 185.950 ;
        RECT 158.800 184.660 159.030 185.950 ;
        RECT 167.090 184.660 167.320 185.950 ;
        RECT 168.020 185.910 168.310 185.950 ;
        RECT 150.510 181.780 150.740 183.480 ;
        RECT 158.800 181.780 159.030 183.480 ;
        RECT 167.090 181.780 167.320 183.480 ;
        RECT 169.580 181.780 174.560 185.950 ;
        RECT 176.510 184.660 176.740 185.950 ;
        RECT 184.800 184.660 185.030 185.950 ;
        RECT 193.090 184.660 193.320 185.950 ;
        RECT 194.020 185.910 194.310 185.950 ;
        RECT 176.510 181.780 176.740 183.480 ;
        RECT 184.800 181.780 185.030 183.480 ;
        RECT 193.090 181.780 193.320 183.480 ;
        RECT 195.580 181.780 200.560 185.950 ;
        RECT 202.510 184.660 202.740 185.950 ;
        RECT 210.800 184.660 211.030 185.950 ;
        RECT 219.090 184.660 219.320 185.950 ;
        RECT 220.020 185.910 220.310 185.950 ;
        RECT 202.510 181.780 202.740 183.480 ;
        RECT 210.800 181.780 211.030 183.480 ;
        RECT 219.090 181.780 219.320 183.480 ;
        RECT 221.580 181.780 226.560 185.950 ;
        RECT 228.510 184.660 228.740 185.950 ;
        RECT 236.800 184.660 237.030 185.950 ;
        RECT 245.090 184.660 245.320 185.950 ;
        RECT 246.020 185.910 246.310 185.950 ;
        RECT 228.510 181.780 228.740 183.480 ;
        RECT 236.800 181.780 237.030 183.480 ;
        RECT 245.090 181.780 245.320 183.480 ;
        RECT 247.580 181.780 252.560 185.950 ;
        RECT 254.510 184.660 254.740 185.950 ;
        RECT 262.800 184.660 263.030 185.950 ;
        RECT 271.090 184.660 271.320 185.950 ;
        RECT 272.020 185.910 272.310 185.950 ;
        RECT 254.510 181.780 254.740 183.480 ;
        RECT 262.800 181.780 263.030 183.480 ;
        RECT 271.090 181.780 271.320 183.480 ;
        RECT 273.580 181.780 278.560 185.950 ;
        RECT 280.510 184.660 280.740 185.950 ;
        RECT 288.800 184.660 289.030 185.950 ;
        RECT 297.090 184.660 297.320 185.950 ;
        RECT 298.020 185.910 298.310 185.950 ;
        RECT 280.510 181.780 280.740 183.480 ;
        RECT 288.800 181.780 289.030 183.480 ;
        RECT 297.090 181.780 297.320 183.480 ;
        RECT 299.580 181.780 304.560 185.950 ;
        RECT 39.400 181.750 63.830 181.780 ;
        RECT 64.480 181.750 70.560 181.780 ;
        RECT 39.400 177.950 70.560 181.750 ;
        RECT 72.250 181.750 89.830 181.780 ;
        RECT 90.480 181.750 96.560 181.780 ;
        RECT 72.250 177.950 96.560 181.750 ;
        RECT 98.250 181.750 115.830 181.780 ;
        RECT 116.480 181.750 122.560 181.780 ;
        RECT 98.250 177.950 122.560 181.750 ;
        RECT 124.250 181.750 141.830 181.780 ;
        RECT 142.480 181.750 148.560 181.780 ;
        RECT 124.250 177.950 148.560 181.750 ;
        RECT 150.250 181.750 167.830 181.780 ;
        RECT 168.480 181.750 174.560 181.780 ;
        RECT 150.250 177.950 174.560 181.750 ;
        RECT 176.250 181.750 193.830 181.780 ;
        RECT 194.480 181.750 200.560 181.780 ;
        RECT 176.250 177.950 200.560 181.750 ;
        RECT 202.250 181.750 219.830 181.780 ;
        RECT 220.480 181.750 226.560 181.780 ;
        RECT 202.250 177.950 226.560 181.750 ;
        RECT 228.250 181.750 245.830 181.780 ;
        RECT 246.480 181.750 252.560 181.780 ;
        RECT 228.250 177.950 252.560 181.750 ;
        RECT 254.250 181.750 271.830 181.780 ;
        RECT 272.480 181.750 278.560 181.780 ;
        RECT 254.250 177.950 278.560 181.750 ;
        RECT 280.250 181.750 297.830 181.780 ;
        RECT 298.480 181.750 304.560 181.780 ;
        RECT 280.250 177.950 304.560 181.750 ;
        RECT 39.400 177.900 48.010 177.950 ;
        RECT 39.400 174.000 44.730 177.900 ;
        RECT 45.980 177.560 48.010 177.900 ;
        RECT 46.510 176.480 46.740 177.560 ;
        RECT 54.800 176.480 55.030 177.950 ;
        RECT 63.090 176.480 63.320 177.950 ;
        RECT 64.020 177.900 64.340 177.950 ;
        RECT 46.510 174.040 46.740 175.300 ;
        RECT 46.360 174.000 47.360 174.040 ;
        RECT 54.800 174.000 55.030 175.300 ;
        RECT 63.090 174.000 63.320 175.300 ;
        RECT 64.020 174.000 64.300 174.010 ;
        RECT 65.580 174.000 70.560 177.950 ;
        RECT 72.510 176.480 72.740 177.950 ;
        RECT 80.800 176.480 81.030 177.950 ;
        RECT 89.090 176.480 89.320 177.950 ;
        RECT 90.020 177.900 90.340 177.950 ;
        RECT 72.510 174.040 72.740 175.300 ;
        RECT 39.400 173.990 45.390 174.000 ;
        RECT 46.360 173.990 70.560 174.000 ;
        RECT 39.400 170.160 70.560 173.990 ;
        RECT 44.550 170.090 47.570 170.160 ;
        RECT 46.510 168.300 46.740 170.090 ;
        RECT 54.800 168.300 55.030 170.160 ;
        RECT 63.090 168.300 63.320 170.160 ;
        RECT 64.020 170.080 64.300 170.160 ;
        RECT 65.580 170.080 70.560 170.160 ;
        RECT 72.360 174.000 73.360 174.040 ;
        RECT 80.800 174.000 81.030 175.300 ;
        RECT 89.090 174.000 89.320 175.300 ;
        RECT 90.020 174.000 90.300 174.010 ;
        RECT 91.580 174.000 96.560 177.950 ;
        RECT 98.510 176.480 98.740 177.950 ;
        RECT 106.800 176.480 107.030 177.950 ;
        RECT 115.090 176.480 115.320 177.950 ;
        RECT 116.020 177.900 116.340 177.950 ;
        RECT 98.510 174.040 98.740 175.300 ;
        RECT 72.360 170.160 96.560 174.000 ;
        RECT 72.360 170.140 73.360 170.160 ;
        RECT 72.510 168.300 72.740 170.140 ;
        RECT 80.800 168.300 81.030 170.160 ;
        RECT 89.090 168.300 89.320 170.160 ;
        RECT 90.020 170.080 90.300 170.160 ;
        RECT 91.580 170.080 96.560 170.160 ;
        RECT 98.360 174.000 99.360 174.040 ;
        RECT 106.800 174.000 107.030 175.300 ;
        RECT 115.090 174.000 115.320 175.300 ;
        RECT 116.020 174.000 116.300 174.010 ;
        RECT 117.580 174.000 122.560 177.950 ;
        RECT 124.510 176.480 124.740 177.950 ;
        RECT 132.800 176.480 133.030 177.950 ;
        RECT 141.090 176.480 141.320 177.950 ;
        RECT 142.020 177.900 142.340 177.950 ;
        RECT 124.510 174.040 124.740 175.300 ;
        RECT 98.360 170.160 122.560 174.000 ;
        RECT 98.360 170.140 99.360 170.160 ;
        RECT 98.510 168.300 98.740 170.140 ;
        RECT 106.800 168.300 107.030 170.160 ;
        RECT 115.090 168.300 115.320 170.160 ;
        RECT 116.020 170.080 116.300 170.160 ;
        RECT 117.580 170.080 122.560 170.160 ;
        RECT 124.360 174.000 125.360 174.040 ;
        RECT 132.800 174.000 133.030 175.300 ;
        RECT 141.090 174.000 141.320 175.300 ;
        RECT 142.020 174.000 142.300 174.010 ;
        RECT 143.580 174.000 148.560 177.950 ;
        RECT 150.510 176.480 150.740 177.950 ;
        RECT 158.800 176.480 159.030 177.950 ;
        RECT 167.090 176.480 167.320 177.950 ;
        RECT 168.020 177.900 168.340 177.950 ;
        RECT 150.510 174.040 150.740 175.300 ;
        RECT 124.360 170.160 148.560 174.000 ;
        RECT 124.360 170.140 125.360 170.160 ;
        RECT 124.510 168.300 124.740 170.140 ;
        RECT 132.800 168.300 133.030 170.160 ;
        RECT 141.090 168.300 141.320 170.160 ;
        RECT 142.020 170.080 142.300 170.160 ;
        RECT 143.580 170.080 148.560 170.160 ;
        RECT 150.360 174.000 151.360 174.040 ;
        RECT 158.800 174.000 159.030 175.300 ;
        RECT 167.090 174.000 167.320 175.300 ;
        RECT 168.020 174.000 168.300 174.010 ;
        RECT 169.580 174.000 174.560 177.950 ;
        RECT 176.510 176.480 176.740 177.950 ;
        RECT 184.800 176.480 185.030 177.950 ;
        RECT 193.090 176.480 193.320 177.950 ;
        RECT 194.020 177.900 194.340 177.950 ;
        RECT 176.510 174.040 176.740 175.300 ;
        RECT 150.360 170.160 174.560 174.000 ;
        RECT 150.360 170.140 151.360 170.160 ;
        RECT 150.510 168.300 150.740 170.140 ;
        RECT 158.800 168.300 159.030 170.160 ;
        RECT 167.090 168.300 167.320 170.160 ;
        RECT 168.020 170.080 168.300 170.160 ;
        RECT 169.580 170.080 174.560 170.160 ;
        RECT 176.360 174.000 177.360 174.040 ;
        RECT 184.800 174.000 185.030 175.300 ;
        RECT 193.090 174.000 193.320 175.300 ;
        RECT 194.020 174.000 194.300 174.010 ;
        RECT 195.580 174.000 200.560 177.950 ;
        RECT 202.510 176.480 202.740 177.950 ;
        RECT 210.800 176.480 211.030 177.950 ;
        RECT 219.090 176.480 219.320 177.950 ;
        RECT 220.020 177.900 220.340 177.950 ;
        RECT 202.510 174.040 202.740 175.300 ;
        RECT 176.360 170.160 200.560 174.000 ;
        RECT 176.360 170.140 177.360 170.160 ;
        RECT 176.510 168.300 176.740 170.140 ;
        RECT 184.800 168.300 185.030 170.160 ;
        RECT 193.090 168.300 193.320 170.160 ;
        RECT 194.020 170.080 194.300 170.160 ;
        RECT 195.580 170.080 200.560 170.160 ;
        RECT 202.360 174.000 203.360 174.040 ;
        RECT 210.800 174.000 211.030 175.300 ;
        RECT 219.090 174.000 219.320 175.300 ;
        RECT 220.020 174.000 220.300 174.010 ;
        RECT 221.580 174.000 226.560 177.950 ;
        RECT 228.510 176.480 228.740 177.950 ;
        RECT 236.800 176.480 237.030 177.950 ;
        RECT 245.090 176.480 245.320 177.950 ;
        RECT 246.020 177.900 246.340 177.950 ;
        RECT 228.510 174.040 228.740 175.300 ;
        RECT 202.360 170.160 226.560 174.000 ;
        RECT 202.360 170.140 203.360 170.160 ;
        RECT 202.510 168.300 202.740 170.140 ;
        RECT 210.800 168.300 211.030 170.160 ;
        RECT 219.090 168.300 219.320 170.160 ;
        RECT 220.020 170.080 220.300 170.160 ;
        RECT 221.580 170.080 226.560 170.160 ;
        RECT 228.360 174.000 229.360 174.040 ;
        RECT 236.800 174.000 237.030 175.300 ;
        RECT 245.090 174.000 245.320 175.300 ;
        RECT 246.020 174.000 246.300 174.010 ;
        RECT 247.580 174.000 252.560 177.950 ;
        RECT 254.510 176.480 254.740 177.950 ;
        RECT 262.800 176.480 263.030 177.950 ;
        RECT 271.090 176.480 271.320 177.950 ;
        RECT 272.020 177.900 272.340 177.950 ;
        RECT 254.510 174.040 254.740 175.300 ;
        RECT 228.360 170.160 252.560 174.000 ;
        RECT 228.360 170.140 229.360 170.160 ;
        RECT 228.510 168.300 228.740 170.140 ;
        RECT 236.800 168.300 237.030 170.160 ;
        RECT 245.090 168.300 245.320 170.160 ;
        RECT 246.020 170.080 246.300 170.160 ;
        RECT 247.580 170.080 252.560 170.160 ;
        RECT 254.360 174.000 255.360 174.040 ;
        RECT 262.800 174.000 263.030 175.300 ;
        RECT 271.090 174.000 271.320 175.300 ;
        RECT 272.020 174.000 272.300 174.010 ;
        RECT 273.580 174.000 278.560 177.950 ;
        RECT 280.510 176.480 280.740 177.950 ;
        RECT 288.800 176.480 289.030 177.950 ;
        RECT 297.090 176.480 297.320 177.950 ;
        RECT 298.020 177.900 298.340 177.950 ;
        RECT 280.510 174.040 280.740 175.300 ;
        RECT 254.360 170.160 278.560 174.000 ;
        RECT 254.360 170.140 255.360 170.160 ;
        RECT 254.510 168.300 254.740 170.140 ;
        RECT 262.800 168.300 263.030 170.160 ;
        RECT 271.090 168.300 271.320 170.160 ;
        RECT 272.020 170.080 272.300 170.160 ;
        RECT 273.580 170.080 278.560 170.160 ;
        RECT 280.360 174.000 281.360 174.040 ;
        RECT 288.800 174.000 289.030 175.300 ;
        RECT 297.090 174.000 297.320 175.300 ;
        RECT 298.020 174.000 298.300 174.010 ;
        RECT 299.580 174.000 304.560 177.950 ;
        RECT 280.360 170.160 304.560 174.000 ;
        RECT 280.360 170.140 281.360 170.160 ;
        RECT 280.510 168.300 280.740 170.140 ;
        RECT 288.800 168.300 289.030 170.160 ;
        RECT 297.090 168.300 297.320 170.160 ;
        RECT 298.020 170.080 298.300 170.160 ;
        RECT 299.580 170.080 304.560 170.160 ;
        RECT 300.970 144.310 304.090 170.080 ;
        RECT 322.920 144.310 335.750 144.330 ;
        RECT 300.970 142.720 335.750 144.310 ;
        RECT 334.990 141.950 335.750 142.720 ;
        RECT 129.090 135.760 129.320 136.660 ;
        RECT 150.990 135.320 151.220 136.220 ;
        RECT 334.990 136.140 335.780 141.950 ;
        RECT 171.780 135.090 172.010 135.990 ;
        RECT 334.990 135.355 335.770 136.140 ;
        RECT 334.990 135.090 336.550 135.355 ;
        RECT 335.370 134.370 336.520 135.090 ;
        RECT 335.350 133.840 336.670 134.370 ;
        RECT 321.040 133.820 323.050 133.830 ;
        RECT 334.260 133.820 336.670 133.840 ;
        RECT 321.040 133.785 336.670 133.820 ;
        RECT 309.190 133.330 336.670 133.785 ;
        RECT 309.190 133.310 323.050 133.330 ;
        RECT 334.260 133.310 336.670 133.330 ;
        RECT 309.190 133.295 321.190 133.310 ;
        RECT 335.350 132.750 336.670 133.310 ;
        RECT 320.990 127.710 332.990 127.720 ;
        RECT 334.930 127.710 336.940 128.050 ;
        RECT 320.990 127.230 336.940 127.710 ;
        RECT 334.930 126.910 336.940 127.230 ;
        RECT 123.540 115.270 125.940 116.980 ;
        RECT 120.710 114.620 125.940 115.270 ;
        RECT 122.050 114.550 125.940 114.620 ;
        RECT 122.050 112.440 125.070 114.550 ;
        RECT 122.410 110.940 124.760 112.440 ;
        RECT 116.830 110.560 124.760 110.940 ;
        RECT 111.430 104.630 112.220 110.410 ;
        RECT 122.410 110.290 124.760 110.560 ;
        RECT 148.320 111.000 149.620 111.130 ;
        RECT 148.320 109.920 149.650 111.000 ;
        RECT 111.270 102.875 112.660 104.630 ;
        RECT 148.370 104.580 149.650 109.920 ;
        RECT 148.340 102.725 149.845 104.580 ;
        RECT 234.220 104.210 236.490 104.740 ;
        RECT 234.250 101.050 236.470 103.090 ;
        RECT 260.210 99.480 262.450 99.930 ;
        RECT 281.620 97.880 283.890 98.350 ;
        RECT 234.240 94.700 236.480 95.170 ;
        RECT 213.840 86.620 216.410 87.680 ;
        RECT 220.440 86.620 222.100 87.350 ;
        RECT 213.840 86.410 222.100 86.620 ;
        RECT 213.840 85.510 216.410 86.410 ;
        RECT 220.440 82.360 222.100 86.410 ;
        RECT 233.260 82.360 234.920 87.370 ;
        RECT 238.280 85.900 240.850 88.070 ;
        RECT 264.840 84.840 267.410 87.010 ;
        RECT 266.070 84.560 266.270 84.840 ;
        RECT 276.340 84.560 278.280 85.330 ;
        RECT 266.070 84.420 278.280 84.560 ;
        RECT 266.110 84.380 278.280 84.420 ;
        RECT 220.440 82.120 234.920 82.360 ;
        RECT 220.440 81.490 222.100 82.120 ;
        RECT 233.260 81.510 234.920 82.120 ;
        RECT 276.340 81.950 278.280 84.380 ;
        RECT 284.290 81.950 286.230 85.470 ;
        RECT 292.020 84.550 294.590 86.720 ;
        RECT 276.340 81.770 286.230 81.950 ;
        RECT 276.340 79.430 278.280 81.770 ;
        RECT 284.290 79.570 286.230 81.770 ;
        RECT 111.105 75.020 112.495 76.775 ;
        RECT 49.460 74.300 51.760 74.770 ;
        RECT 49.400 72.720 51.760 74.300 ;
        RECT 85.310 73.310 86.500 74.670 ;
        RECT 147.820 74.460 149.740 76.860 ;
        RECT 49.460 72.370 51.760 72.720 ;
        RECT 27.910 70.380 28.790 71.470 ;
        RECT 45.740 70.900 47.410 70.960 ;
        RECT 45.720 70.730 47.410 70.900 ;
        RECT 45.740 70.670 47.410 70.730 ;
        RECT 81.200 70.530 81.430 71.430 ;
        RECT 27.650 69.430 29.330 69.730 ;
        RECT 45.920 69.660 47.600 69.940 ;
        RECT 45.780 67.840 47.450 67.900 ;
        RECT 45.760 67.670 47.450 67.840 ;
        RECT 45.780 67.610 47.450 67.670 ;
        RECT 27.680 66.910 29.360 67.210 ;
        RECT 45.960 66.600 47.640 66.880 ;
        RECT 45.760 64.950 47.430 65.010 ;
        RECT 45.740 64.780 47.430 64.950 ;
        RECT 45.760 64.720 47.430 64.780 ;
        RECT 27.660 64.580 29.340 64.620 ;
        RECT 27.660 64.350 29.350 64.580 ;
        RECT 27.660 64.320 29.340 64.350 ;
        RECT 45.940 63.710 47.620 63.990 ;
        RECT 45.800 62.080 47.470 62.140 ;
        RECT 27.660 62.030 29.340 62.080 ;
        RECT 27.660 61.800 29.350 62.030 ;
        RECT 45.780 61.910 47.470 62.080 ;
        RECT 45.800 61.850 47.470 61.910 ;
        RECT 27.660 61.780 29.340 61.800 ;
        RECT 45.980 60.840 47.660 61.120 ;
        RECT 27.660 59.480 29.340 59.530 ;
        RECT 27.660 59.250 29.350 59.480 ;
        RECT 27.660 59.230 29.340 59.250 ;
        RECT 45.800 59.190 47.470 59.250 ;
        RECT 45.780 59.020 47.470 59.190 ;
        RECT 45.800 58.960 47.470 59.020 ;
        RECT 193.000 58.750 194.190 60.110 ;
        RECT 45.980 57.950 47.660 58.230 ;
        RECT 27.660 56.930 29.340 56.980 ;
        RECT 27.660 56.700 29.350 56.930 ;
        RECT 27.660 56.680 29.340 56.700 ;
        RECT 45.800 56.300 47.470 56.360 ;
        RECT 45.780 56.130 47.470 56.300 ;
        RECT 45.800 56.070 47.470 56.130 ;
        RECT 45.980 55.060 47.660 55.340 ;
        RECT 27.660 54.380 29.340 54.430 ;
        RECT 197.390 54.380 197.620 55.280 ;
        RECT 27.660 54.150 29.350 54.380 ;
        RECT 27.660 54.130 29.340 54.150 ;
        RECT 45.820 53.390 47.490 53.450 ;
        RECT 45.800 53.220 47.490 53.390 ;
        RECT 45.820 53.160 47.490 53.220 ;
        RECT 46.000 52.150 47.680 52.430 ;
        RECT 27.660 51.830 29.340 51.880 ;
        RECT 27.660 51.600 29.350 51.830 ;
        RECT 27.660 51.580 29.340 51.600 ;
        RECT 45.800 50.510 47.470 50.570 ;
        RECT 45.780 50.340 47.470 50.510 ;
        RECT 45.800 50.280 47.470 50.340 ;
        RECT 27.660 49.280 29.340 49.330 ;
        RECT 27.660 49.050 29.350 49.280 ;
        RECT 45.980 49.270 47.660 49.550 ;
        RECT 27.660 49.030 29.340 49.050 ;
        RECT 147.380 48.250 148.800 50.060 ;
        RECT 45.780 47.660 47.450 47.720 ;
        RECT 45.760 47.490 47.450 47.660 ;
        RECT 45.780 47.430 47.450 47.490 ;
        RECT 45.960 46.420 47.640 46.700 ;
        RECT 85.020 46.560 86.210 47.920 ;
        RECT 111.100 45.710 112.035 47.295 ;
        RECT 81.590 44.780 81.820 45.680 ;
        RECT 250.560 40.160 252.720 40.520 ;
        RECT 250.840 35.220 253.000 35.580 ;
        RECT 284.260 26.630 284.550 28.350 ;
        RECT 242.670 22.670 244.760 24.740 ;
        RECT 249.520 23.840 249.800 24.840 ;
        RECT 270.370 23.820 270.670 25.490 ;
        RECT 275.270 23.810 275.600 25.480 ;
        RECT 283.780 24.590 284.090 25.130 ;
        RECT 283.820 24.570 284.090 24.590 ;
        RECT 119.090 18.370 120.490 19.540 ;
        RECT 123.580 14.130 123.810 15.030 ;
        RECT 140.490 14.040 140.720 14.940 ;
        RECT 158.960 14.130 159.190 15.030 ;
        RECT 693.660 6.850 720.830 8.355 ;
        RECT 693.660 1.295 693.890 6.850 ;
        RECT 695.520 1.490 695.750 6.850 ;
        RECT 698.100 1.490 698.330 6.850 ;
        RECT 700.680 1.490 700.910 6.850 ;
        RECT 703.260 1.490 703.490 6.850 ;
        RECT 705.840 1.490 706.070 6.850 ;
        RECT 708.420 1.490 708.650 6.850 ;
        RECT 711.000 1.490 711.230 6.850 ;
        RECT 713.580 1.490 713.810 6.850 ;
        RECT 716.160 1.490 716.390 6.850 ;
        RECT 718.740 1.490 718.970 6.850 ;
        RECT 720.600 1.295 720.830 6.850 ;
        RECT 694.720 1.055 695.260 1.285 ;
        RECT 696.010 1.055 696.550 1.285 ;
        RECT 697.300 1.055 697.840 1.285 ;
        RECT 698.590 1.055 699.130 1.285 ;
        RECT 699.880 1.055 700.420 1.285 ;
        RECT 701.170 1.055 701.710 1.285 ;
        RECT 702.460 1.055 703.000 1.285 ;
        RECT 703.750 1.055 704.290 1.285 ;
        RECT 705.040 1.055 705.580 1.285 ;
        RECT 706.330 1.055 706.870 1.285 ;
        RECT 707.620 1.055 708.160 1.285 ;
        RECT 708.910 1.055 709.450 1.285 ;
        RECT 710.200 1.055 710.740 1.285 ;
        RECT 711.490 1.055 712.030 1.285 ;
        RECT 712.780 1.055 713.320 1.285 ;
        RECT 714.070 1.055 714.610 1.285 ;
        RECT 715.360 1.055 715.900 1.285 ;
        RECT 716.650 1.055 717.190 1.285 ;
        RECT 717.940 1.055 718.480 1.285 ;
        RECT 719.230 1.055 719.770 1.285 ;
      LAYER via ;
        RECT 40.380 323.190 43.810 326.180 ;
        RECT 66.380 323.190 69.810 326.180 ;
        RECT 92.380 323.190 95.810 326.180 ;
        RECT 118.380 323.190 121.810 326.180 ;
        RECT 144.380 323.190 147.810 326.180 ;
        RECT 170.380 323.190 173.810 326.180 ;
        RECT 196.380 323.190 199.810 326.180 ;
        RECT 222.380 323.190 225.810 326.180 ;
        RECT 248.380 323.190 251.810 326.180 ;
        RECT 274.380 323.190 277.810 326.180 ;
        RECT 300.380 323.190 303.810 326.180 ;
        RECT 40.380 313.190 43.810 316.180 ;
        RECT 66.380 313.190 69.810 316.180 ;
        RECT 92.380 313.190 95.810 316.180 ;
        RECT 118.380 313.190 121.810 316.180 ;
        RECT 144.380 313.190 147.810 316.180 ;
        RECT 170.380 313.190 173.810 316.180 ;
        RECT 196.380 313.190 199.810 316.180 ;
        RECT 222.380 313.190 225.810 316.180 ;
        RECT 248.380 313.190 251.810 316.180 ;
        RECT 274.380 313.190 277.810 316.180 ;
        RECT 300.380 313.190 303.810 316.180 ;
        RECT 40.380 303.190 43.810 306.180 ;
        RECT 66.380 303.190 69.810 306.180 ;
        RECT 92.380 303.190 95.810 306.180 ;
        RECT 118.380 303.190 121.810 306.180 ;
        RECT 144.380 303.190 147.810 306.180 ;
        RECT 170.380 303.190 173.810 306.180 ;
        RECT 196.380 303.190 199.810 306.180 ;
        RECT 222.380 303.190 225.810 306.180 ;
        RECT 248.380 303.190 251.810 306.180 ;
        RECT 274.380 303.190 277.810 306.180 ;
        RECT 300.380 303.190 303.810 306.180 ;
        RECT 40.380 293.190 43.810 296.180 ;
        RECT 66.380 293.190 69.810 296.180 ;
        RECT 92.380 293.190 95.810 296.180 ;
        RECT 118.380 293.190 121.810 296.180 ;
        RECT 144.380 293.190 147.810 296.180 ;
        RECT 170.380 293.190 173.810 296.180 ;
        RECT 196.380 293.190 199.810 296.180 ;
        RECT 222.380 293.190 225.810 296.180 ;
        RECT 248.380 293.190 251.810 296.180 ;
        RECT 274.380 293.190 277.810 296.180 ;
        RECT 300.380 293.190 303.810 296.180 ;
        RECT 40.380 283.190 43.810 286.180 ;
        RECT 66.380 283.190 69.810 286.180 ;
        RECT 92.380 283.190 95.810 286.180 ;
        RECT 118.380 283.190 121.810 286.180 ;
        RECT 144.380 283.190 147.810 286.180 ;
        RECT 170.380 283.190 173.810 286.180 ;
        RECT 196.380 283.190 199.810 286.180 ;
        RECT 222.380 283.190 225.810 286.180 ;
        RECT 248.380 283.190 251.810 286.180 ;
        RECT 274.380 283.190 277.810 286.180 ;
        RECT 300.380 283.190 303.810 286.180 ;
        RECT 40.380 273.190 43.810 276.180 ;
        RECT 66.380 273.190 69.810 276.180 ;
        RECT 92.380 273.190 95.810 276.180 ;
        RECT 118.380 273.190 121.810 276.180 ;
        RECT 144.380 273.190 147.810 276.180 ;
        RECT 170.380 273.190 173.810 276.180 ;
        RECT 196.380 273.190 199.810 276.180 ;
        RECT 222.380 273.190 225.810 276.180 ;
        RECT 248.380 273.190 251.810 276.180 ;
        RECT 274.380 273.190 277.810 276.180 ;
        RECT 300.380 273.190 303.810 276.180 ;
        RECT 40.380 263.190 43.810 266.180 ;
        RECT 66.380 263.190 69.810 266.180 ;
        RECT 92.380 263.190 95.810 266.180 ;
        RECT 118.380 263.190 121.810 266.180 ;
        RECT 144.380 263.190 147.810 266.180 ;
        RECT 170.380 263.190 173.810 266.180 ;
        RECT 196.380 263.190 199.810 266.180 ;
        RECT 222.380 263.190 225.810 266.180 ;
        RECT 248.380 263.190 251.810 266.180 ;
        RECT 274.380 263.190 277.810 266.180 ;
        RECT 300.380 263.190 303.810 266.180 ;
        RECT 40.380 253.190 43.810 256.180 ;
        RECT 66.380 253.190 69.810 256.180 ;
        RECT 92.380 253.190 95.810 256.180 ;
        RECT 118.380 253.190 121.810 256.180 ;
        RECT 144.380 253.190 147.810 256.180 ;
        RECT 170.380 253.190 173.810 256.180 ;
        RECT 196.380 253.190 199.810 256.180 ;
        RECT 222.380 253.190 225.810 256.180 ;
        RECT 248.380 253.190 251.810 256.180 ;
        RECT 274.380 253.190 277.810 256.180 ;
        RECT 300.380 253.190 303.810 256.180 ;
        RECT 40.380 241.190 43.810 244.180 ;
        RECT 66.380 241.190 69.810 244.180 ;
        RECT 92.380 241.190 95.810 244.180 ;
        RECT 118.380 241.190 121.810 244.180 ;
        RECT 144.380 241.190 147.810 244.180 ;
        RECT 170.380 241.190 173.810 244.180 ;
        RECT 196.380 241.190 199.810 244.180 ;
        RECT 222.380 241.190 225.810 244.180 ;
        RECT 248.380 241.190 251.810 244.180 ;
        RECT 274.380 241.190 277.810 244.180 ;
        RECT 300.380 241.190 303.810 244.180 ;
        RECT 690.020 250.510 690.420 250.910 ;
        RECT 690.820 250.510 691.220 250.910 ;
        RECT 691.620 250.510 692.020 250.910 ;
        RECT 692.420 250.510 692.820 250.910 ;
        RECT 693.220 250.510 693.620 250.910 ;
        RECT 694.020 250.510 694.420 250.910 ;
        RECT 694.820 250.510 695.220 250.910 ;
        RECT 695.620 250.510 696.020 250.910 ;
        RECT 696.420 250.510 696.820 250.910 ;
        RECT 697.220 250.510 697.620 250.910 ;
        RECT 698.020 250.510 698.420 250.910 ;
        RECT 698.820 250.510 699.220 250.910 ;
        RECT 699.620 250.510 700.020 250.910 ;
        RECT 700.420 250.510 700.820 250.910 ;
        RECT 701.220 250.510 701.620 250.910 ;
        RECT 702.020 250.510 702.420 250.910 ;
        RECT 702.820 250.510 703.220 250.910 ;
        RECT 703.620 250.510 704.020 250.910 ;
        RECT 704.420 250.510 704.820 250.910 ;
        RECT 705.220 250.510 705.620 250.910 ;
        RECT 706.020 250.510 706.420 250.910 ;
        RECT 706.820 250.510 707.220 250.910 ;
        RECT 707.620 250.510 708.020 250.910 ;
        RECT 708.420 250.510 708.820 250.910 ;
        RECT 709.220 250.510 709.620 250.910 ;
        RECT 710.020 250.510 710.420 250.910 ;
        RECT 710.820 250.510 711.220 250.910 ;
        RECT 711.620 250.510 712.020 250.910 ;
        RECT 712.420 250.510 712.820 250.910 ;
        RECT 713.220 250.510 713.620 250.910 ;
        RECT 714.020 250.510 714.420 250.910 ;
        RECT 690.020 249.710 690.420 250.110 ;
        RECT 690.820 249.710 691.220 250.110 ;
        RECT 691.620 249.710 692.020 250.110 ;
        RECT 692.420 249.710 692.820 250.110 ;
        RECT 693.220 249.710 693.620 250.110 ;
        RECT 694.020 249.710 694.420 250.110 ;
        RECT 694.820 249.710 695.220 250.110 ;
        RECT 695.620 249.710 696.020 250.110 ;
        RECT 696.420 249.710 696.820 250.110 ;
        RECT 697.220 249.710 697.620 250.110 ;
        RECT 698.020 249.710 698.420 250.110 ;
        RECT 698.820 249.710 699.220 250.110 ;
        RECT 699.620 249.710 700.020 250.110 ;
        RECT 700.420 249.710 700.820 250.110 ;
        RECT 701.220 249.710 701.620 250.110 ;
        RECT 702.020 249.710 702.420 250.110 ;
        RECT 702.820 249.710 703.220 250.110 ;
        RECT 703.620 249.710 704.020 250.110 ;
        RECT 704.420 249.710 704.820 250.110 ;
        RECT 705.220 249.710 705.620 250.110 ;
        RECT 706.020 249.710 706.420 250.110 ;
        RECT 706.820 249.710 707.220 250.110 ;
        RECT 707.620 249.710 708.020 250.110 ;
        RECT 708.420 249.710 708.820 250.110 ;
        RECT 709.220 249.710 709.620 250.110 ;
        RECT 710.020 249.710 710.420 250.110 ;
        RECT 710.820 249.710 711.220 250.110 ;
        RECT 711.620 249.710 712.020 250.110 ;
        RECT 712.420 249.710 712.820 250.110 ;
        RECT 713.220 249.710 713.620 250.110 ;
        RECT 714.020 249.710 714.420 250.110 ;
        RECT 40.380 231.190 43.810 234.180 ;
        RECT 66.380 231.190 69.810 234.180 ;
        RECT 92.380 231.190 95.810 234.180 ;
        RECT 118.380 231.190 121.810 234.180 ;
        RECT 144.380 231.190 147.810 234.180 ;
        RECT 170.380 231.190 173.810 234.180 ;
        RECT 196.380 231.190 199.810 234.180 ;
        RECT 222.380 231.190 225.810 234.180 ;
        RECT 248.380 231.190 251.810 234.180 ;
        RECT 274.380 231.190 277.810 234.180 ;
        RECT 300.380 231.190 303.810 234.180 ;
        RECT 40.380 221.190 43.810 224.180 ;
        RECT 66.380 221.190 69.810 224.180 ;
        RECT 92.380 221.190 95.810 224.180 ;
        RECT 118.380 221.190 121.810 224.180 ;
        RECT 144.380 221.190 147.810 224.180 ;
        RECT 170.380 221.190 173.810 224.180 ;
        RECT 196.380 221.190 199.810 224.180 ;
        RECT 222.380 221.190 225.810 224.180 ;
        RECT 248.380 221.190 251.810 224.180 ;
        RECT 274.380 221.190 277.810 224.180 ;
        RECT 300.380 221.190 303.810 224.180 ;
        RECT 40.380 211.190 43.810 214.180 ;
        RECT 66.380 211.190 69.810 214.180 ;
        RECT 92.380 211.190 95.810 214.180 ;
        RECT 118.380 211.190 121.810 214.180 ;
        RECT 144.380 211.190 147.810 214.180 ;
        RECT 170.380 211.190 173.810 214.180 ;
        RECT 196.380 211.190 199.810 214.180 ;
        RECT 222.380 211.190 225.810 214.180 ;
        RECT 248.380 211.190 251.810 214.180 ;
        RECT 274.380 211.190 277.810 214.180 ;
        RECT 300.380 211.190 303.810 214.180 ;
        RECT 40.380 201.190 43.810 204.180 ;
        RECT 66.380 201.190 69.810 204.180 ;
        RECT 92.380 201.190 95.810 204.180 ;
        RECT 118.380 201.190 121.810 204.180 ;
        RECT 144.380 201.190 147.810 204.180 ;
        RECT 170.380 201.190 173.810 204.180 ;
        RECT 196.380 201.190 199.810 204.180 ;
        RECT 222.380 201.190 225.810 204.180 ;
        RECT 248.380 201.190 251.810 204.180 ;
        RECT 274.380 201.190 277.810 204.180 ;
        RECT 300.380 201.190 303.810 204.180 ;
        RECT 40.380 191.190 43.810 194.180 ;
        RECT 66.380 191.190 69.810 194.180 ;
        RECT 92.380 191.190 95.810 194.180 ;
        RECT 118.380 191.190 121.810 194.180 ;
        RECT 144.380 191.190 147.810 194.180 ;
        RECT 170.380 191.190 173.810 194.180 ;
        RECT 196.380 191.190 199.810 194.180 ;
        RECT 222.380 191.190 225.810 194.180 ;
        RECT 248.380 191.190 251.810 194.180 ;
        RECT 274.380 191.190 277.810 194.180 ;
        RECT 300.380 191.190 303.810 194.180 ;
        RECT 40.380 181.190 43.810 184.180 ;
        RECT 66.380 181.190 69.810 184.180 ;
        RECT 92.380 181.190 95.810 184.180 ;
        RECT 118.380 181.190 121.810 184.180 ;
        RECT 144.380 181.190 147.810 184.180 ;
        RECT 170.380 181.190 173.810 184.180 ;
        RECT 196.380 181.190 199.810 184.180 ;
        RECT 222.380 181.190 225.810 184.180 ;
        RECT 248.380 181.190 251.810 184.180 ;
        RECT 274.380 181.190 277.810 184.180 ;
        RECT 300.380 181.190 303.810 184.180 ;
        RECT 40.380 171.190 43.810 174.180 ;
        RECT 66.380 171.190 69.810 174.180 ;
        RECT 92.380 171.190 95.810 174.180 ;
        RECT 118.380 171.190 121.810 174.180 ;
        RECT 144.380 171.190 147.810 174.180 ;
        RECT 170.380 171.190 173.810 174.180 ;
        RECT 196.380 171.190 199.810 174.180 ;
        RECT 222.380 171.190 225.810 174.180 ;
        RECT 248.380 171.190 251.810 174.180 ;
        RECT 274.380 171.190 277.810 174.180 ;
        RECT 300.380 171.190 303.810 174.180 ;
        RECT 335.740 133.170 336.410 133.950 ;
        RECT 335.750 127.210 336.320 127.730 ;
        RECT 111.360 102.970 112.555 104.535 ;
        RECT 148.515 102.855 149.625 104.460 ;
        RECT 234.280 104.290 236.440 104.640 ;
        RECT 234.280 102.680 236.450 103.050 ;
        RECT 234.270 101.100 236.440 101.470 ;
        RECT 260.260 99.530 262.420 99.880 ;
        RECT 281.670 97.940 283.830 98.290 ;
        RECT 234.280 94.750 236.440 95.110 ;
        RECT 214.310 86.000 215.940 87.200 ;
        RECT 238.750 86.390 240.380 87.590 ;
        RECT 265.310 85.330 266.940 86.530 ;
        RECT 292.490 85.040 294.120 86.240 ;
        RECT 111.305 75.180 112.220 76.705 ;
        RECT 148.340 75.070 149.310 76.610 ;
        RECT 49.610 72.640 51.570 74.640 ;
        RECT 85.460 73.530 86.340 74.420 ;
        RECT 28.070 70.650 28.600 71.370 ;
        RECT 45.770 70.690 47.360 70.950 ;
        RECT 27.700 69.450 29.280 69.710 ;
        RECT 45.980 69.660 47.540 69.920 ;
        RECT 45.810 67.630 47.400 67.890 ;
        RECT 27.740 66.920 29.320 67.180 ;
        RECT 46.020 66.600 47.580 66.860 ;
        RECT 45.790 64.740 47.380 65.000 ;
        RECT 27.730 64.330 29.310 64.590 ;
        RECT 46.000 63.710 47.560 63.970 ;
        RECT 27.730 61.790 29.310 62.050 ;
        RECT 45.830 61.870 47.420 62.130 ;
        RECT 46.040 60.840 47.600 61.100 ;
        RECT 27.730 59.240 29.310 59.500 ;
        RECT 45.830 58.980 47.420 59.240 ;
        RECT 193.150 58.970 194.030 59.860 ;
        RECT 46.040 57.950 47.600 58.210 ;
        RECT 27.730 56.690 29.310 56.950 ;
        RECT 45.830 56.090 47.420 56.350 ;
        RECT 46.040 55.060 47.600 55.320 ;
        RECT 27.730 54.140 29.310 54.400 ;
        RECT 45.850 53.180 47.440 53.440 ;
        RECT 46.060 52.150 47.620 52.410 ;
        RECT 27.730 51.590 29.310 51.850 ;
        RECT 45.830 50.300 47.420 50.560 ;
        RECT 27.730 49.040 29.310 49.300 ;
        RECT 46.040 49.270 47.600 49.530 ;
        RECT 147.560 48.330 148.640 49.915 ;
        RECT 45.810 47.450 47.400 47.710 ;
        RECT 85.170 46.780 86.050 47.670 ;
        RECT 46.020 46.420 47.580 46.680 ;
        RECT 111.165 45.850 111.945 47.210 ;
        RECT 250.650 40.190 252.660 40.480 ;
        RECT 250.940 35.250 252.930 35.550 ;
        RECT 284.270 26.690 284.550 28.300 ;
        RECT 242.950 22.900 244.460 24.580 ;
        RECT 249.530 23.900 249.800 24.780 ;
        RECT 270.400 23.890 270.660 25.440 ;
        RECT 275.310 23.880 275.590 25.430 ;
        RECT 283.810 24.640 284.080 25.060 ;
        RECT 119.420 18.640 120.280 19.270 ;
        RECT 695.310 7.790 695.710 8.190 ;
        RECT 696.110 7.790 696.510 8.190 ;
        RECT 696.910 7.790 697.310 8.190 ;
        RECT 697.710 7.790 698.110 8.190 ;
        RECT 698.510 7.790 698.910 8.190 ;
        RECT 699.310 7.790 699.710 8.190 ;
        RECT 700.110 7.790 700.510 8.190 ;
        RECT 700.910 7.790 701.310 8.190 ;
        RECT 701.710 7.790 702.110 8.190 ;
        RECT 702.510 7.790 702.910 8.190 ;
        RECT 703.310 7.790 703.710 8.190 ;
        RECT 704.110 7.790 704.510 8.190 ;
        RECT 704.910 7.790 705.310 8.190 ;
        RECT 705.710 7.790 706.110 8.190 ;
        RECT 706.510 7.790 706.910 8.190 ;
        RECT 707.310 7.790 707.710 8.190 ;
        RECT 708.110 7.790 708.510 8.190 ;
        RECT 708.910 7.790 709.310 8.190 ;
        RECT 709.710 7.790 710.110 8.190 ;
        RECT 710.510 7.790 710.910 8.190 ;
        RECT 711.310 7.790 711.710 8.190 ;
        RECT 712.110 7.790 712.510 8.190 ;
        RECT 712.910 7.790 713.310 8.190 ;
        RECT 713.710 7.790 714.110 8.190 ;
        RECT 714.510 7.790 714.910 8.190 ;
        RECT 715.310 7.790 715.710 8.190 ;
        RECT 716.110 7.790 716.510 8.190 ;
        RECT 716.910 7.790 717.310 8.190 ;
        RECT 717.710 7.790 718.110 8.190 ;
        RECT 718.510 7.790 718.910 8.190 ;
        RECT 719.310 7.790 719.710 8.190 ;
        RECT 695.310 6.990 695.710 7.390 ;
        RECT 696.110 6.990 696.510 7.390 ;
        RECT 696.910 6.990 697.310 7.390 ;
        RECT 697.710 6.990 698.110 7.390 ;
        RECT 698.510 6.990 698.910 7.390 ;
        RECT 699.310 6.990 699.710 7.390 ;
        RECT 700.110 6.990 700.510 7.390 ;
        RECT 700.910 6.990 701.310 7.390 ;
        RECT 701.710 6.990 702.110 7.390 ;
        RECT 702.510 6.990 702.910 7.390 ;
        RECT 703.310 6.990 703.710 7.390 ;
        RECT 704.110 6.990 704.510 7.390 ;
        RECT 704.910 6.990 705.310 7.390 ;
        RECT 705.710 6.990 706.110 7.390 ;
        RECT 706.510 6.990 706.910 7.390 ;
        RECT 707.310 6.990 707.710 7.390 ;
        RECT 708.110 6.990 708.510 7.390 ;
        RECT 708.910 6.990 709.310 7.390 ;
        RECT 709.710 6.990 710.110 7.390 ;
        RECT 710.510 6.990 710.910 7.390 ;
        RECT 711.310 6.990 711.710 7.390 ;
        RECT 712.110 6.990 712.510 7.390 ;
        RECT 712.910 6.990 713.310 7.390 ;
        RECT 713.710 6.990 714.110 7.390 ;
        RECT 714.510 6.990 714.910 7.390 ;
        RECT 715.310 6.990 715.710 7.390 ;
        RECT 716.110 6.990 716.510 7.390 ;
        RECT 716.910 6.990 717.310 7.390 ;
        RECT 717.710 6.990 718.110 7.390 ;
        RECT 718.510 6.990 718.910 7.390 ;
        RECT 719.310 6.990 719.710 7.390 ;
      LAYER met2 ;
        RECT 39.650 322.330 44.490 327.060 ;
        RECT 65.650 322.330 70.490 327.060 ;
        RECT 91.650 322.330 96.490 327.060 ;
        RECT 117.650 322.330 122.490 327.060 ;
        RECT 143.650 322.330 148.490 327.060 ;
        RECT 169.650 322.330 174.490 327.060 ;
        RECT 195.650 322.330 200.490 327.060 ;
        RECT 221.650 322.330 226.490 327.060 ;
        RECT 247.650 322.330 252.490 327.060 ;
        RECT 273.650 322.330 278.490 327.060 ;
        RECT 299.650 322.330 304.490 327.060 ;
        RECT 39.650 312.330 44.490 317.060 ;
        RECT 65.650 312.330 70.490 317.060 ;
        RECT 91.650 312.330 96.490 317.060 ;
        RECT 117.650 312.330 122.490 317.060 ;
        RECT 143.650 312.330 148.490 317.060 ;
        RECT 169.650 312.330 174.490 317.060 ;
        RECT 195.650 312.330 200.490 317.060 ;
        RECT 221.650 312.330 226.490 317.060 ;
        RECT 247.650 312.330 252.490 317.060 ;
        RECT 273.650 312.330 278.490 317.060 ;
        RECT 299.650 312.330 304.490 317.060 ;
        RECT 39.650 302.330 44.490 307.060 ;
        RECT 65.650 302.330 70.490 307.060 ;
        RECT 91.650 302.330 96.490 307.060 ;
        RECT 117.650 302.330 122.490 307.060 ;
        RECT 143.650 302.330 148.490 307.060 ;
        RECT 169.650 302.330 174.490 307.060 ;
        RECT 195.650 302.330 200.490 307.060 ;
        RECT 221.650 302.330 226.490 307.060 ;
        RECT 247.650 302.330 252.490 307.060 ;
        RECT 273.650 302.330 278.490 307.060 ;
        RECT 299.650 302.330 304.490 307.060 ;
        RECT 39.650 292.330 44.490 297.060 ;
        RECT 65.650 292.330 70.490 297.060 ;
        RECT 91.650 292.330 96.490 297.060 ;
        RECT 117.650 292.330 122.490 297.060 ;
        RECT 143.650 292.330 148.490 297.060 ;
        RECT 169.650 292.330 174.490 297.060 ;
        RECT 195.650 292.330 200.490 297.060 ;
        RECT 221.650 292.330 226.490 297.060 ;
        RECT 247.650 292.330 252.490 297.060 ;
        RECT 273.650 292.330 278.490 297.060 ;
        RECT 299.650 292.330 304.490 297.060 ;
        RECT 39.650 282.330 44.490 287.060 ;
        RECT 65.650 282.330 70.490 287.060 ;
        RECT 91.650 282.330 96.490 287.060 ;
        RECT 117.650 282.330 122.490 287.060 ;
        RECT 143.650 282.330 148.490 287.060 ;
        RECT 169.650 282.330 174.490 287.060 ;
        RECT 195.650 282.330 200.490 287.060 ;
        RECT 221.650 282.330 226.490 287.060 ;
        RECT 247.650 282.330 252.490 287.060 ;
        RECT 273.650 282.330 278.490 287.060 ;
        RECT 299.650 282.330 304.490 287.060 ;
        RECT 39.650 272.330 44.490 277.060 ;
        RECT 65.650 272.330 70.490 277.060 ;
        RECT 91.650 272.330 96.490 277.060 ;
        RECT 117.650 272.330 122.490 277.060 ;
        RECT 143.650 272.330 148.490 277.060 ;
        RECT 169.650 272.330 174.490 277.060 ;
        RECT 195.650 272.330 200.490 277.060 ;
        RECT 221.650 272.330 226.490 277.060 ;
        RECT 247.650 272.330 252.490 277.060 ;
        RECT 273.650 272.330 278.490 277.060 ;
        RECT 299.650 272.330 304.490 277.060 ;
        RECT 39.650 262.330 44.490 267.060 ;
        RECT 65.650 262.330 70.490 267.060 ;
        RECT 91.650 262.330 96.490 267.060 ;
        RECT 117.650 262.330 122.490 267.060 ;
        RECT 143.650 262.330 148.490 267.060 ;
        RECT 169.650 262.330 174.490 267.060 ;
        RECT 195.650 262.330 200.490 267.060 ;
        RECT 221.650 262.330 226.490 267.060 ;
        RECT 247.650 262.330 252.490 267.060 ;
        RECT 273.650 262.330 278.490 267.060 ;
        RECT 299.650 262.330 304.490 267.060 ;
        RECT 39.650 252.330 44.490 257.060 ;
        RECT 65.650 252.330 70.490 257.060 ;
        RECT 91.650 252.330 96.490 257.060 ;
        RECT 117.650 252.330 122.490 257.060 ;
        RECT 143.650 252.330 148.490 257.060 ;
        RECT 169.650 252.330 174.490 257.060 ;
        RECT 195.650 252.330 200.490 257.060 ;
        RECT 221.650 252.330 226.490 257.060 ;
        RECT 247.650 252.330 252.490 257.060 ;
        RECT 273.650 252.330 278.490 257.060 ;
        RECT 299.650 252.330 304.490 257.060 ;
        RECT 689.520 249.510 715.020 251.310 ;
        RECT 39.650 240.330 44.490 245.060 ;
        RECT 65.650 240.330 70.490 245.060 ;
        RECT 91.650 240.330 96.490 245.060 ;
        RECT 117.650 240.330 122.490 245.060 ;
        RECT 143.650 240.330 148.490 245.060 ;
        RECT 169.650 240.330 174.490 245.060 ;
        RECT 195.650 240.330 200.490 245.060 ;
        RECT 221.650 240.330 226.490 245.060 ;
        RECT 247.650 240.330 252.490 245.060 ;
        RECT 273.650 240.330 278.490 245.060 ;
        RECT 299.650 240.330 304.490 245.060 ;
        RECT 39.650 230.330 44.490 235.060 ;
        RECT 65.650 230.330 70.490 235.060 ;
        RECT 91.650 230.330 96.490 235.060 ;
        RECT 117.650 230.330 122.490 235.060 ;
        RECT 143.650 230.330 148.490 235.060 ;
        RECT 169.650 230.330 174.490 235.060 ;
        RECT 195.650 230.330 200.490 235.060 ;
        RECT 221.650 230.330 226.490 235.060 ;
        RECT 247.650 230.330 252.490 235.060 ;
        RECT 273.650 230.330 278.490 235.060 ;
        RECT 299.650 230.330 304.490 235.060 ;
        RECT 39.650 220.330 44.490 225.060 ;
        RECT 65.650 220.330 70.490 225.060 ;
        RECT 91.650 220.330 96.490 225.060 ;
        RECT 117.650 220.330 122.490 225.060 ;
        RECT 143.650 220.330 148.490 225.060 ;
        RECT 169.650 220.330 174.490 225.060 ;
        RECT 195.650 220.330 200.490 225.060 ;
        RECT 221.650 220.330 226.490 225.060 ;
        RECT 247.650 220.330 252.490 225.060 ;
        RECT 273.650 220.330 278.490 225.060 ;
        RECT 299.650 220.330 304.490 225.060 ;
        RECT 39.650 210.330 44.490 215.060 ;
        RECT 65.650 210.330 70.490 215.060 ;
        RECT 91.650 210.330 96.490 215.060 ;
        RECT 117.650 210.330 122.490 215.060 ;
        RECT 143.650 210.330 148.490 215.060 ;
        RECT 169.650 210.330 174.490 215.060 ;
        RECT 195.650 210.330 200.490 215.060 ;
        RECT 221.650 210.330 226.490 215.060 ;
        RECT 247.650 210.330 252.490 215.060 ;
        RECT 273.650 210.330 278.490 215.060 ;
        RECT 299.650 210.330 304.490 215.060 ;
        RECT 39.650 200.330 44.490 205.060 ;
        RECT 65.650 200.330 70.490 205.060 ;
        RECT 91.650 200.330 96.490 205.060 ;
        RECT 117.650 200.330 122.490 205.060 ;
        RECT 143.650 200.330 148.490 205.060 ;
        RECT 169.650 200.330 174.490 205.060 ;
        RECT 195.650 200.330 200.490 205.060 ;
        RECT 221.650 200.330 226.490 205.060 ;
        RECT 247.650 200.330 252.490 205.060 ;
        RECT 273.650 200.330 278.490 205.060 ;
        RECT 299.650 200.330 304.490 205.060 ;
        RECT 39.650 190.330 44.490 195.060 ;
        RECT 65.650 190.330 70.490 195.060 ;
        RECT 91.650 190.330 96.490 195.060 ;
        RECT 117.650 190.330 122.490 195.060 ;
        RECT 143.650 190.330 148.490 195.060 ;
        RECT 169.650 190.330 174.490 195.060 ;
        RECT 195.650 190.330 200.490 195.060 ;
        RECT 221.650 190.330 226.490 195.060 ;
        RECT 247.650 190.330 252.490 195.060 ;
        RECT 273.650 190.330 278.490 195.060 ;
        RECT 299.650 190.330 304.490 195.060 ;
        RECT 39.650 180.330 44.490 185.060 ;
        RECT 65.650 180.330 70.490 185.060 ;
        RECT 91.650 180.330 96.490 185.060 ;
        RECT 117.650 180.330 122.490 185.060 ;
        RECT 143.650 180.330 148.490 185.060 ;
        RECT 169.650 180.330 174.490 185.060 ;
        RECT 195.650 180.330 200.490 185.060 ;
        RECT 221.650 180.330 226.490 185.060 ;
        RECT 247.650 180.330 252.490 185.060 ;
        RECT 273.650 180.330 278.490 185.060 ;
        RECT 299.650 180.330 304.490 185.060 ;
        RECT 39.650 170.330 44.490 175.060 ;
        RECT 65.650 170.330 70.490 175.060 ;
        RECT 91.650 170.330 96.490 175.060 ;
        RECT 117.650 170.330 122.490 175.060 ;
        RECT 143.650 170.330 148.490 175.060 ;
        RECT 169.650 170.330 174.490 175.060 ;
        RECT 195.650 170.330 200.490 175.060 ;
        RECT 221.650 170.330 226.490 175.060 ;
        RECT 247.650 170.330 252.490 175.060 ;
        RECT 273.650 170.330 278.490 175.060 ;
        RECT 299.650 170.330 304.490 175.060 ;
        RECT 335.670 127.060 336.550 134.110 ;
        RECT 111.270 102.875 112.660 104.630 ;
        RECT 148.340 102.725 149.845 104.580 ;
        RECT 234.220 104.210 236.490 104.740 ;
        RECT 234.220 101.030 236.520 103.130 ;
        RECT 260.210 99.480 262.450 99.930 ;
        RECT 261.290 99.180 261.620 99.480 ;
        RECT 268.080 99.180 268.440 99.210 ;
        RECT 261.290 98.870 268.440 99.180 ;
        RECT 261.290 98.860 261.620 98.870 ;
        RECT 234.240 95.120 236.480 95.170 ;
        RECT 233.030 94.840 236.480 95.120 ;
        RECT 233.030 90.390 233.270 94.840 ;
        RECT 234.240 94.700 236.480 94.840 ;
        RECT 233.000 88.060 233.300 90.390 ;
        RECT 238.280 88.060 240.850 88.070 ;
        RECT 233.000 87.890 240.850 88.060 ;
        RECT 233.010 87.870 240.850 87.890 ;
        RECT 213.840 85.510 216.410 87.680 ;
        RECT 238.280 85.900 240.850 87.870 ;
        RECT 264.840 85.950 267.410 87.010 ;
        RECT 268.080 85.950 268.440 98.870 ;
        RECT 281.620 97.880 283.890 98.350 ;
        RECT 264.840 85.570 268.450 85.950 ;
        RECT 264.840 84.840 267.410 85.570 ;
        RECT 268.080 85.540 268.440 85.570 ;
        RECT 292.020 84.550 294.590 86.720 ;
        RECT 49.460 74.300 51.760 74.770 ;
        RECT 49.250 74.290 51.760 74.300 ;
        RECT 48.850 72.960 51.760 74.290 ;
        RECT 28.090 71.470 28.480 71.530 ;
        RECT 27.910 70.380 28.790 71.470 ;
        RECT 48.850 71.320 49.200 72.960 ;
        RECT 49.590 72.370 51.760 72.960 ;
        RECT 84.770 73.800 112.980 77.090 ;
        RECT 147.820 74.460 149.740 76.860 ;
        RECT 84.770 72.710 106.090 73.800 ;
        RECT 49.590 72.330 49.740 72.370 ;
        RECT 45.730 70.960 47.410 70.970 ;
        RECT 48.850 70.960 49.260 71.320 ;
        RECT 45.720 70.670 49.260 70.960 ;
        RECT 45.730 70.660 47.410 70.670 ;
        RECT 28.090 69.750 28.480 70.380 ;
        RECT 45.970 69.940 46.170 70.660 ;
        RECT 28.090 69.730 28.540 69.750 ;
        RECT 27.650 69.430 29.330 69.730 ;
        RECT 45.920 69.650 47.600 69.940 ;
        RECT 28.290 67.210 28.540 69.430 ;
        RECT 48.850 67.910 49.260 70.670 ;
        RECT 45.760 67.600 49.260 67.910 ;
        RECT 27.680 66.910 29.360 67.210 ;
        RECT 28.290 64.620 28.540 66.910 ;
        RECT 46.010 66.880 46.210 67.600 ;
        RECT 45.960 66.590 47.640 66.880 ;
        RECT 45.750 65.010 47.430 65.020 ;
        RECT 48.850 65.010 49.260 67.600 ;
        RECT 45.750 64.720 49.260 65.010 ;
        RECT 45.750 64.710 47.430 64.720 ;
        RECT 27.660 64.320 29.340 64.620 ;
        RECT 28.290 62.080 28.540 64.320 ;
        RECT 45.990 63.990 46.190 64.710 ;
        RECT 45.940 63.700 47.620 63.990 ;
        RECT 48.850 62.170 49.260 64.720 ;
        RECT 27.660 61.780 29.340 62.080 ;
        RECT 45.770 61.830 49.260 62.170 ;
        RECT 28.290 59.530 28.540 61.780 ;
        RECT 46.030 61.120 46.230 61.830 ;
        RECT 45.980 60.830 47.660 61.120 ;
        RECT 27.660 59.230 29.340 59.530 ;
        RECT 48.850 59.270 49.260 61.830 ;
        RECT 28.290 56.980 28.540 59.230 ;
        RECT 45.790 58.950 49.260 59.270 ;
        RECT 46.030 58.230 46.230 58.950 ;
        RECT 45.980 57.940 47.660 58.230 ;
        RECT 27.660 56.680 29.340 56.980 ;
        RECT 28.290 54.430 28.540 56.680 ;
        RECT 48.850 56.390 49.260 58.950 ;
        RECT 193.000 58.750 194.190 60.110 ;
        RECT 45.750 56.080 49.260 56.390 ;
        RECT 45.790 56.060 47.470 56.080 ;
        RECT 46.030 55.340 46.230 56.060 ;
        RECT 45.980 55.050 47.660 55.340 ;
        RECT 27.660 54.130 29.340 54.430 ;
        RECT 28.290 51.880 28.540 54.130 ;
        RECT 48.850 53.490 49.260 56.080 ;
        RECT 45.780 53.180 49.260 53.490 ;
        RECT 45.810 53.150 47.490 53.180 ;
        RECT 46.050 52.430 46.250 53.150 ;
        RECT 46.000 52.140 47.680 52.430 ;
        RECT 27.660 51.580 29.340 51.880 ;
        RECT 28.290 49.330 28.540 51.580 ;
        RECT 48.850 50.580 49.260 53.180 ;
        RECT 45.750 50.300 49.260 50.580 ;
        RECT 45.790 50.270 47.470 50.300 ;
        RECT 46.030 49.550 46.230 50.270 ;
        RECT 27.660 49.030 29.340 49.330 ;
        RECT 45.980 49.260 47.660 49.550 ;
        RECT 28.290 48.980 28.540 49.030 ;
        RECT 48.850 47.730 49.260 50.300 ;
        RECT 147.325 48.195 148.840 50.095 ;
        RECT 45.760 47.420 49.260 47.730 ;
        RECT 46.010 46.700 46.210 47.420 ;
        RECT 48.850 46.850 49.260 47.420 ;
        RECT 45.960 46.410 47.640 46.700 ;
        RECT 85.020 46.560 86.210 47.920 ;
        RECT 111.010 45.685 112.175 47.310 ;
        RECT 250.560 40.490 252.720 40.520 ;
        RECT 249.740 40.480 252.720 40.490 ;
        RECT 249.560 40.170 252.720 40.480 ;
        RECT 249.560 37.880 250.180 40.170 ;
        RECT 250.560 40.160 252.720 40.170 ;
        RECT 243.580 37.840 250.380 37.880 ;
        RECT 243.540 36.700 250.380 37.840 ;
        RECT 243.540 24.740 244.210 36.700 ;
        RECT 249.560 36.540 250.180 36.700 ;
        RECT 249.560 35.600 250.210 36.540 ;
        RECT 249.550 35.150 253.020 35.600 ;
        RECT 249.560 35.130 250.210 35.150 ;
        RECT 249.570 35.100 250.210 35.130 ;
        RECT 284.260 26.630 284.550 28.350 ;
        RECT 242.670 22.670 244.760 24.740 ;
        RECT 249.470 23.840 249.850 24.850 ;
        RECT 270.330 23.810 270.730 25.520 ;
        RECT 275.270 23.810 275.600 25.480 ;
        RECT 283.780 24.590 284.080 25.130 ;
        RECT 119.090 18.370 120.490 19.540 ;
        RECT 694.810 6.790 720.310 8.590 ;
      LAYER via2 ;
        RECT 40.380 323.190 43.810 326.180 ;
        RECT 66.380 323.190 69.810 326.180 ;
        RECT 92.380 323.190 95.810 326.180 ;
        RECT 118.380 323.190 121.810 326.180 ;
        RECT 144.380 323.190 147.810 326.180 ;
        RECT 170.380 323.190 173.810 326.180 ;
        RECT 196.380 323.190 199.810 326.180 ;
        RECT 222.380 323.190 225.810 326.180 ;
        RECT 248.380 323.190 251.810 326.180 ;
        RECT 274.380 323.190 277.810 326.180 ;
        RECT 300.380 323.190 303.810 326.180 ;
        RECT 40.380 313.190 43.810 316.180 ;
        RECT 66.380 313.190 69.810 316.180 ;
        RECT 92.380 313.190 95.810 316.180 ;
        RECT 118.380 313.190 121.810 316.180 ;
        RECT 144.380 313.190 147.810 316.180 ;
        RECT 170.380 313.190 173.810 316.180 ;
        RECT 196.380 313.190 199.810 316.180 ;
        RECT 222.380 313.190 225.810 316.180 ;
        RECT 248.380 313.190 251.810 316.180 ;
        RECT 274.380 313.190 277.810 316.180 ;
        RECT 300.380 313.190 303.810 316.180 ;
        RECT 40.380 303.190 43.810 306.180 ;
        RECT 66.380 303.190 69.810 306.180 ;
        RECT 92.380 303.190 95.810 306.180 ;
        RECT 118.380 303.190 121.810 306.180 ;
        RECT 144.380 303.190 147.810 306.180 ;
        RECT 170.380 303.190 173.810 306.180 ;
        RECT 196.380 303.190 199.810 306.180 ;
        RECT 222.380 303.190 225.810 306.180 ;
        RECT 248.380 303.190 251.810 306.180 ;
        RECT 274.380 303.190 277.810 306.180 ;
        RECT 300.380 303.190 303.810 306.180 ;
        RECT 40.380 293.190 43.810 296.180 ;
        RECT 66.380 293.190 69.810 296.180 ;
        RECT 92.380 293.190 95.810 296.180 ;
        RECT 118.380 293.190 121.810 296.180 ;
        RECT 144.380 293.190 147.810 296.180 ;
        RECT 170.380 293.190 173.810 296.180 ;
        RECT 196.380 293.190 199.810 296.180 ;
        RECT 222.380 293.190 225.810 296.180 ;
        RECT 248.380 293.190 251.810 296.180 ;
        RECT 274.380 293.190 277.810 296.180 ;
        RECT 300.380 293.190 303.810 296.180 ;
        RECT 40.380 283.190 43.810 286.180 ;
        RECT 66.380 283.190 69.810 286.180 ;
        RECT 92.380 283.190 95.810 286.180 ;
        RECT 118.380 283.190 121.810 286.180 ;
        RECT 144.380 283.190 147.810 286.180 ;
        RECT 170.380 283.190 173.810 286.180 ;
        RECT 196.380 283.190 199.810 286.180 ;
        RECT 222.380 283.190 225.810 286.180 ;
        RECT 248.380 283.190 251.810 286.180 ;
        RECT 274.380 283.190 277.810 286.180 ;
        RECT 300.380 283.190 303.810 286.180 ;
        RECT 40.380 273.190 43.810 276.180 ;
        RECT 66.380 273.190 69.810 276.180 ;
        RECT 92.380 273.190 95.810 276.180 ;
        RECT 118.380 273.190 121.810 276.180 ;
        RECT 144.380 273.190 147.810 276.180 ;
        RECT 170.380 273.190 173.810 276.180 ;
        RECT 196.380 273.190 199.810 276.180 ;
        RECT 222.380 273.190 225.810 276.180 ;
        RECT 248.380 273.190 251.810 276.180 ;
        RECT 274.380 273.190 277.810 276.180 ;
        RECT 300.380 273.190 303.810 276.180 ;
        RECT 40.380 263.190 43.810 266.180 ;
        RECT 66.380 263.190 69.810 266.180 ;
        RECT 92.380 263.190 95.810 266.180 ;
        RECT 118.380 263.190 121.810 266.180 ;
        RECT 144.380 263.190 147.810 266.180 ;
        RECT 170.380 263.190 173.810 266.180 ;
        RECT 196.380 263.190 199.810 266.180 ;
        RECT 222.380 263.190 225.810 266.180 ;
        RECT 248.380 263.190 251.810 266.180 ;
        RECT 274.380 263.190 277.810 266.180 ;
        RECT 300.380 263.190 303.810 266.180 ;
        RECT 40.380 253.190 43.810 256.180 ;
        RECT 66.380 253.190 69.810 256.180 ;
        RECT 92.380 253.190 95.810 256.180 ;
        RECT 118.380 253.190 121.810 256.180 ;
        RECT 144.380 253.190 147.810 256.180 ;
        RECT 170.380 253.190 173.810 256.180 ;
        RECT 196.380 253.190 199.810 256.180 ;
        RECT 222.380 253.190 225.810 256.180 ;
        RECT 248.380 253.190 251.810 256.180 ;
        RECT 274.380 253.190 277.810 256.180 ;
        RECT 300.380 253.190 303.810 256.180 ;
        RECT 690.020 250.510 690.420 250.910 ;
        RECT 690.820 250.510 691.220 250.910 ;
        RECT 691.620 250.510 692.020 250.910 ;
        RECT 692.420 250.510 692.820 250.910 ;
        RECT 693.220 250.510 693.620 250.910 ;
        RECT 694.020 250.510 694.420 250.910 ;
        RECT 694.820 250.510 695.220 250.910 ;
        RECT 695.620 250.510 696.020 250.910 ;
        RECT 696.420 250.510 696.820 250.910 ;
        RECT 697.220 250.510 697.620 250.910 ;
        RECT 698.020 250.510 698.420 250.910 ;
        RECT 698.820 250.510 699.220 250.910 ;
        RECT 699.620 250.510 700.020 250.910 ;
        RECT 700.420 250.510 700.820 250.910 ;
        RECT 701.220 250.510 701.620 250.910 ;
        RECT 702.020 250.510 702.420 250.910 ;
        RECT 702.820 250.510 703.220 250.910 ;
        RECT 703.620 250.510 704.020 250.910 ;
        RECT 704.420 250.510 704.820 250.910 ;
        RECT 705.220 250.510 705.620 250.910 ;
        RECT 706.020 250.510 706.420 250.910 ;
        RECT 706.820 250.510 707.220 250.910 ;
        RECT 707.620 250.510 708.020 250.910 ;
        RECT 708.420 250.510 708.820 250.910 ;
        RECT 709.220 250.510 709.620 250.910 ;
        RECT 710.020 250.510 710.420 250.910 ;
        RECT 710.820 250.510 711.220 250.910 ;
        RECT 711.620 250.510 712.020 250.910 ;
        RECT 712.420 250.510 712.820 250.910 ;
        RECT 713.220 250.510 713.620 250.910 ;
        RECT 714.020 250.510 714.420 250.910 ;
        RECT 690.020 249.710 690.420 250.110 ;
        RECT 690.820 249.710 691.220 250.110 ;
        RECT 691.620 249.710 692.020 250.110 ;
        RECT 692.420 249.710 692.820 250.110 ;
        RECT 693.220 249.710 693.620 250.110 ;
        RECT 694.020 249.710 694.420 250.110 ;
        RECT 694.820 249.710 695.220 250.110 ;
        RECT 695.620 249.710 696.020 250.110 ;
        RECT 696.420 249.710 696.820 250.110 ;
        RECT 697.220 249.710 697.620 250.110 ;
        RECT 698.020 249.710 698.420 250.110 ;
        RECT 698.820 249.710 699.220 250.110 ;
        RECT 699.620 249.710 700.020 250.110 ;
        RECT 700.420 249.710 700.820 250.110 ;
        RECT 701.220 249.710 701.620 250.110 ;
        RECT 702.020 249.710 702.420 250.110 ;
        RECT 702.820 249.710 703.220 250.110 ;
        RECT 703.620 249.710 704.020 250.110 ;
        RECT 704.420 249.710 704.820 250.110 ;
        RECT 705.220 249.710 705.620 250.110 ;
        RECT 706.020 249.710 706.420 250.110 ;
        RECT 706.820 249.710 707.220 250.110 ;
        RECT 707.620 249.710 708.020 250.110 ;
        RECT 708.420 249.710 708.820 250.110 ;
        RECT 709.220 249.710 709.620 250.110 ;
        RECT 710.020 249.710 710.420 250.110 ;
        RECT 710.820 249.710 711.220 250.110 ;
        RECT 711.620 249.710 712.020 250.110 ;
        RECT 712.420 249.710 712.820 250.110 ;
        RECT 713.220 249.710 713.620 250.110 ;
        RECT 714.020 249.710 714.420 250.110 ;
        RECT 40.380 241.190 43.810 244.180 ;
        RECT 66.380 241.190 69.810 244.180 ;
        RECT 92.380 241.190 95.810 244.180 ;
        RECT 118.380 241.190 121.810 244.180 ;
        RECT 144.380 241.190 147.810 244.180 ;
        RECT 170.380 241.190 173.810 244.180 ;
        RECT 196.380 241.190 199.810 244.180 ;
        RECT 222.380 241.190 225.810 244.180 ;
        RECT 248.380 241.190 251.810 244.180 ;
        RECT 274.380 241.190 277.810 244.180 ;
        RECT 300.380 241.190 303.810 244.180 ;
        RECT 40.380 231.190 43.810 234.180 ;
        RECT 66.380 231.190 69.810 234.180 ;
        RECT 92.380 231.190 95.810 234.180 ;
        RECT 118.380 231.190 121.810 234.180 ;
        RECT 144.380 231.190 147.810 234.180 ;
        RECT 170.380 231.190 173.810 234.180 ;
        RECT 196.380 231.190 199.810 234.180 ;
        RECT 222.380 231.190 225.810 234.180 ;
        RECT 248.380 231.190 251.810 234.180 ;
        RECT 274.380 231.190 277.810 234.180 ;
        RECT 300.380 231.190 303.810 234.180 ;
        RECT 40.380 221.190 43.810 224.180 ;
        RECT 66.380 221.190 69.810 224.180 ;
        RECT 92.380 221.190 95.810 224.180 ;
        RECT 118.380 221.190 121.810 224.180 ;
        RECT 144.380 221.190 147.810 224.180 ;
        RECT 170.380 221.190 173.810 224.180 ;
        RECT 196.380 221.190 199.810 224.180 ;
        RECT 222.380 221.190 225.810 224.180 ;
        RECT 248.380 221.190 251.810 224.180 ;
        RECT 274.380 221.190 277.810 224.180 ;
        RECT 300.380 221.190 303.810 224.180 ;
        RECT 40.380 211.190 43.810 214.180 ;
        RECT 66.380 211.190 69.810 214.180 ;
        RECT 92.380 211.190 95.810 214.180 ;
        RECT 118.380 211.190 121.810 214.180 ;
        RECT 144.380 211.190 147.810 214.180 ;
        RECT 170.380 211.190 173.810 214.180 ;
        RECT 196.380 211.190 199.810 214.180 ;
        RECT 222.380 211.190 225.810 214.180 ;
        RECT 248.380 211.190 251.810 214.180 ;
        RECT 274.380 211.190 277.810 214.180 ;
        RECT 300.380 211.190 303.810 214.180 ;
        RECT 40.380 201.190 43.810 204.180 ;
        RECT 66.380 201.190 69.810 204.180 ;
        RECT 92.380 201.190 95.810 204.180 ;
        RECT 118.380 201.190 121.810 204.180 ;
        RECT 144.380 201.190 147.810 204.180 ;
        RECT 170.380 201.190 173.810 204.180 ;
        RECT 196.380 201.190 199.810 204.180 ;
        RECT 222.380 201.190 225.810 204.180 ;
        RECT 248.380 201.190 251.810 204.180 ;
        RECT 274.380 201.190 277.810 204.180 ;
        RECT 300.380 201.190 303.810 204.180 ;
        RECT 40.380 191.190 43.810 194.180 ;
        RECT 66.380 191.190 69.810 194.180 ;
        RECT 92.380 191.190 95.810 194.180 ;
        RECT 118.380 191.190 121.810 194.180 ;
        RECT 144.380 191.190 147.810 194.180 ;
        RECT 170.380 191.190 173.810 194.180 ;
        RECT 196.380 191.190 199.810 194.180 ;
        RECT 222.380 191.190 225.810 194.180 ;
        RECT 248.380 191.190 251.810 194.180 ;
        RECT 274.380 191.190 277.810 194.180 ;
        RECT 300.380 191.190 303.810 194.180 ;
        RECT 40.380 181.190 43.810 184.180 ;
        RECT 66.380 181.190 69.810 184.180 ;
        RECT 92.380 181.190 95.810 184.180 ;
        RECT 118.380 181.190 121.810 184.180 ;
        RECT 144.380 181.190 147.810 184.180 ;
        RECT 170.380 181.190 173.810 184.180 ;
        RECT 196.380 181.190 199.810 184.180 ;
        RECT 222.380 181.190 225.810 184.180 ;
        RECT 248.380 181.190 251.810 184.180 ;
        RECT 274.380 181.190 277.810 184.180 ;
        RECT 300.380 181.190 303.810 184.180 ;
        RECT 40.380 171.190 43.810 174.180 ;
        RECT 66.380 171.190 69.810 174.180 ;
        RECT 92.380 171.190 95.810 174.180 ;
        RECT 118.380 171.190 121.810 174.180 ;
        RECT 144.380 171.190 147.810 174.180 ;
        RECT 170.380 171.190 173.810 174.180 ;
        RECT 196.380 171.190 199.810 174.180 ;
        RECT 222.380 171.190 225.810 174.180 ;
        RECT 248.380 171.190 251.810 174.180 ;
        RECT 274.380 171.190 277.810 174.180 ;
        RECT 300.380 171.190 303.810 174.180 ;
        RECT 111.360 102.970 112.555 104.535 ;
        RECT 148.410 102.775 149.775 104.525 ;
        RECT 234.280 104.290 236.440 104.660 ;
        RECT 234.280 102.690 236.440 103.060 ;
        RECT 234.280 101.090 236.450 101.470 ;
        RECT 214.310 86.000 215.940 87.200 ;
        RECT 238.750 86.390 240.380 87.590 ;
        RECT 265.310 85.330 266.940 86.530 ;
        RECT 281.670 97.940 283.830 98.290 ;
        RECT 292.490 85.040 294.120 86.240 ;
        RECT 111.305 75.180 112.220 76.705 ;
        RECT 49.610 72.640 51.570 74.640 ;
        RECT 148.340 75.070 149.310 76.610 ;
        RECT 85.460 73.530 86.340 74.420 ;
        RECT 193.150 58.970 194.030 59.860 ;
        RECT 147.500 48.250 148.730 49.995 ;
        RECT 85.170 46.780 86.050 47.670 ;
        RECT 111.110 45.880 112.015 47.160 ;
        RECT 284.270 26.690 284.550 28.300 ;
        RECT 242.950 22.900 244.460 24.580 ;
        RECT 249.530 23.900 249.810 24.780 ;
        RECT 270.400 23.890 270.680 25.440 ;
        RECT 275.310 23.880 275.590 25.430 ;
        RECT 283.790 24.640 284.080 25.060 ;
        RECT 119.420 18.640 120.280 19.270 ;
        RECT 695.310 7.790 695.710 8.190 ;
        RECT 696.110 7.790 696.510 8.190 ;
        RECT 696.910 7.790 697.310 8.190 ;
        RECT 697.710 7.790 698.110 8.190 ;
        RECT 698.510 7.790 698.910 8.190 ;
        RECT 699.310 7.790 699.710 8.190 ;
        RECT 700.110 7.790 700.510 8.190 ;
        RECT 700.910 7.790 701.310 8.190 ;
        RECT 701.710 7.790 702.110 8.190 ;
        RECT 702.510 7.790 702.910 8.190 ;
        RECT 703.310 7.790 703.710 8.190 ;
        RECT 704.110 7.790 704.510 8.190 ;
        RECT 704.910 7.790 705.310 8.190 ;
        RECT 705.710 7.790 706.110 8.190 ;
        RECT 706.510 7.790 706.910 8.190 ;
        RECT 707.310 7.790 707.710 8.190 ;
        RECT 708.110 7.790 708.510 8.190 ;
        RECT 708.910 7.790 709.310 8.190 ;
        RECT 709.710 7.790 710.110 8.190 ;
        RECT 710.510 7.790 710.910 8.190 ;
        RECT 711.310 7.790 711.710 8.190 ;
        RECT 712.110 7.790 712.510 8.190 ;
        RECT 712.910 7.790 713.310 8.190 ;
        RECT 713.710 7.790 714.110 8.190 ;
        RECT 714.510 7.790 714.910 8.190 ;
        RECT 715.310 7.790 715.710 8.190 ;
        RECT 716.110 7.790 716.510 8.190 ;
        RECT 716.910 7.790 717.310 8.190 ;
        RECT 717.710 7.790 718.110 8.190 ;
        RECT 718.510 7.790 718.910 8.190 ;
        RECT 719.310 7.790 719.710 8.190 ;
        RECT 695.310 6.990 695.710 7.390 ;
        RECT 696.110 6.990 696.510 7.390 ;
        RECT 696.910 6.990 697.310 7.390 ;
        RECT 697.710 6.990 698.110 7.390 ;
        RECT 698.510 6.990 698.910 7.390 ;
        RECT 699.310 6.990 699.710 7.390 ;
        RECT 700.110 6.990 700.510 7.390 ;
        RECT 700.910 6.990 701.310 7.390 ;
        RECT 701.710 6.990 702.110 7.390 ;
        RECT 702.510 6.990 702.910 7.390 ;
        RECT 703.310 6.990 703.710 7.390 ;
        RECT 704.110 6.990 704.510 7.390 ;
        RECT 704.910 6.990 705.310 7.390 ;
        RECT 705.710 6.990 706.110 7.390 ;
        RECT 706.510 6.990 706.910 7.390 ;
        RECT 707.310 6.990 707.710 7.390 ;
        RECT 708.110 6.990 708.510 7.390 ;
        RECT 708.910 6.990 709.310 7.390 ;
        RECT 709.710 6.990 710.110 7.390 ;
        RECT 710.510 6.990 710.910 7.390 ;
        RECT 711.310 6.990 711.710 7.390 ;
        RECT 712.110 6.990 712.510 7.390 ;
        RECT 712.910 6.990 713.310 7.390 ;
        RECT 713.710 6.990 714.110 7.390 ;
        RECT 714.510 6.990 714.910 7.390 ;
        RECT 715.310 6.990 715.710 7.390 ;
        RECT 716.110 6.990 716.510 7.390 ;
        RECT 716.910 6.990 717.310 7.390 ;
        RECT 717.710 6.990 718.110 7.390 ;
        RECT 718.510 6.990 718.910 7.390 ;
        RECT 719.310 6.990 719.710 7.390 ;
      LAYER met3 ;
        RECT 39.650 322.330 44.490 327.060 ;
        RECT 65.650 322.330 70.490 327.060 ;
        RECT 91.650 322.330 96.490 327.060 ;
        RECT 117.650 322.330 122.490 327.060 ;
        RECT 143.650 322.330 148.490 327.060 ;
        RECT 169.650 322.330 174.490 327.060 ;
        RECT 195.650 322.330 200.490 327.060 ;
        RECT 221.650 322.330 226.490 327.060 ;
        RECT 247.650 322.330 252.490 327.060 ;
        RECT 273.650 322.330 278.490 327.060 ;
        RECT 299.650 322.330 304.490 327.060 ;
        RECT 39.650 312.330 44.490 317.060 ;
        RECT 65.650 312.330 70.490 317.060 ;
        RECT 91.650 312.330 96.490 317.060 ;
        RECT 117.650 312.330 122.490 317.060 ;
        RECT 143.650 312.330 148.490 317.060 ;
        RECT 169.650 312.330 174.490 317.060 ;
        RECT 195.650 312.330 200.490 317.060 ;
        RECT 221.650 312.330 226.490 317.060 ;
        RECT 247.650 312.330 252.490 317.060 ;
        RECT 273.650 312.330 278.490 317.060 ;
        RECT 299.650 312.330 304.490 317.060 ;
        RECT 39.650 302.330 44.490 307.060 ;
        RECT 65.650 302.330 70.490 307.060 ;
        RECT 91.650 302.330 96.490 307.060 ;
        RECT 117.650 302.330 122.490 307.060 ;
        RECT 143.650 302.330 148.490 307.060 ;
        RECT 169.650 302.330 174.490 307.060 ;
        RECT 195.650 302.330 200.490 307.060 ;
        RECT 221.650 302.330 226.490 307.060 ;
        RECT 247.650 302.330 252.490 307.060 ;
        RECT 273.650 302.330 278.490 307.060 ;
        RECT 299.650 302.330 304.490 307.060 ;
        RECT 39.650 292.330 44.490 297.060 ;
        RECT 65.650 292.330 70.490 297.060 ;
        RECT 91.650 292.330 96.490 297.060 ;
        RECT 117.650 292.330 122.490 297.060 ;
        RECT 143.650 292.330 148.490 297.060 ;
        RECT 169.650 292.330 174.490 297.060 ;
        RECT 195.650 292.330 200.490 297.060 ;
        RECT 221.650 292.330 226.490 297.060 ;
        RECT 247.650 292.330 252.490 297.060 ;
        RECT 273.650 292.330 278.490 297.060 ;
        RECT 299.650 292.330 304.490 297.060 ;
        RECT 39.650 282.330 44.490 287.060 ;
        RECT 65.650 282.330 70.490 287.060 ;
        RECT 91.650 282.330 96.490 287.060 ;
        RECT 117.650 282.330 122.490 287.060 ;
        RECT 143.650 282.330 148.490 287.060 ;
        RECT 169.650 282.330 174.490 287.060 ;
        RECT 195.650 282.330 200.490 287.060 ;
        RECT 221.650 282.330 226.490 287.060 ;
        RECT 247.650 282.330 252.490 287.060 ;
        RECT 273.650 282.330 278.490 287.060 ;
        RECT 299.650 282.330 304.490 287.060 ;
        RECT 39.650 272.330 44.490 277.060 ;
        RECT 65.650 272.330 70.490 277.060 ;
        RECT 91.650 272.330 96.490 277.060 ;
        RECT 117.650 272.330 122.490 277.060 ;
        RECT 143.650 272.330 148.490 277.060 ;
        RECT 169.650 272.330 174.490 277.060 ;
        RECT 195.650 272.330 200.490 277.060 ;
        RECT 221.650 272.330 226.490 277.060 ;
        RECT 247.650 272.330 252.490 277.060 ;
        RECT 273.650 272.330 278.490 277.060 ;
        RECT 299.650 272.330 304.490 277.060 ;
        RECT 39.650 262.330 44.490 267.060 ;
        RECT 65.650 262.330 70.490 267.060 ;
        RECT 91.650 262.330 96.490 267.060 ;
        RECT 117.650 262.330 122.490 267.060 ;
        RECT 143.650 262.330 148.490 267.060 ;
        RECT 169.650 262.330 174.490 267.060 ;
        RECT 195.650 262.330 200.490 267.060 ;
        RECT 221.650 262.330 226.490 267.060 ;
        RECT 247.650 262.330 252.490 267.060 ;
        RECT 273.650 262.330 278.490 267.060 ;
        RECT 299.650 262.330 304.490 267.060 ;
        RECT 39.650 252.330 44.490 257.060 ;
        RECT 65.650 252.330 70.490 257.060 ;
        RECT 91.650 252.330 96.490 257.060 ;
        RECT 117.650 252.330 122.490 257.060 ;
        RECT 143.650 252.330 148.490 257.060 ;
        RECT 169.650 252.330 174.490 257.060 ;
        RECT 195.650 252.330 200.490 257.060 ;
        RECT 221.650 252.330 226.490 257.060 ;
        RECT 247.650 252.330 252.490 257.060 ;
        RECT 273.650 252.330 278.490 257.060 ;
        RECT 299.650 252.330 304.490 257.060 ;
        RECT 689.520 249.510 715.020 251.310 ;
        RECT 39.650 240.330 44.490 245.060 ;
        RECT 65.650 240.330 70.490 245.060 ;
        RECT 91.650 240.330 96.490 245.060 ;
        RECT 117.650 240.330 122.490 245.060 ;
        RECT 143.650 240.330 148.490 245.060 ;
        RECT 169.650 240.330 174.490 245.060 ;
        RECT 195.650 240.330 200.490 245.060 ;
        RECT 221.650 240.330 226.490 245.060 ;
        RECT 247.650 240.330 252.490 245.060 ;
        RECT 273.650 240.330 278.490 245.060 ;
        RECT 299.650 240.330 304.490 245.060 ;
        RECT 39.650 230.330 44.490 235.060 ;
        RECT 65.650 230.330 70.490 235.060 ;
        RECT 91.650 230.330 96.490 235.060 ;
        RECT 117.650 230.330 122.490 235.060 ;
        RECT 143.650 230.330 148.490 235.060 ;
        RECT 169.650 230.330 174.490 235.060 ;
        RECT 195.650 230.330 200.490 235.060 ;
        RECT 221.650 230.330 226.490 235.060 ;
        RECT 247.650 230.330 252.490 235.060 ;
        RECT 273.650 230.330 278.490 235.060 ;
        RECT 299.650 230.330 304.490 235.060 ;
        RECT 39.650 220.330 44.490 225.060 ;
        RECT 65.650 220.330 70.490 225.060 ;
        RECT 91.650 220.330 96.490 225.060 ;
        RECT 117.650 220.330 122.490 225.060 ;
        RECT 143.650 220.330 148.490 225.060 ;
        RECT 169.650 220.330 174.490 225.060 ;
        RECT 195.650 220.330 200.490 225.060 ;
        RECT 221.650 220.330 226.490 225.060 ;
        RECT 247.650 220.330 252.490 225.060 ;
        RECT 273.650 220.330 278.490 225.060 ;
        RECT 299.650 220.330 304.490 225.060 ;
        RECT 39.650 210.330 44.490 215.060 ;
        RECT 65.650 210.330 70.490 215.060 ;
        RECT 91.650 210.330 96.490 215.060 ;
        RECT 117.650 210.330 122.490 215.060 ;
        RECT 143.650 210.330 148.490 215.060 ;
        RECT 169.650 210.330 174.490 215.060 ;
        RECT 195.650 210.330 200.490 215.060 ;
        RECT 221.650 210.330 226.490 215.060 ;
        RECT 247.650 210.330 252.490 215.060 ;
        RECT 273.650 210.330 278.490 215.060 ;
        RECT 299.650 210.330 304.490 215.060 ;
        RECT 39.650 200.330 44.490 205.060 ;
        RECT 65.650 200.330 70.490 205.060 ;
        RECT 91.650 200.330 96.490 205.060 ;
        RECT 117.650 200.330 122.490 205.060 ;
        RECT 143.650 200.330 148.490 205.060 ;
        RECT 169.650 200.330 174.490 205.060 ;
        RECT 195.650 200.330 200.490 205.060 ;
        RECT 221.650 200.330 226.490 205.060 ;
        RECT 247.650 200.330 252.490 205.060 ;
        RECT 273.650 200.330 278.490 205.060 ;
        RECT 299.650 200.330 304.490 205.060 ;
        RECT 39.650 190.330 44.490 195.060 ;
        RECT 65.650 190.330 70.490 195.060 ;
        RECT 91.650 190.330 96.490 195.060 ;
        RECT 117.650 190.330 122.490 195.060 ;
        RECT 143.650 190.330 148.490 195.060 ;
        RECT 169.650 190.330 174.490 195.060 ;
        RECT 195.650 190.330 200.490 195.060 ;
        RECT 221.650 190.330 226.490 195.060 ;
        RECT 247.650 190.330 252.490 195.060 ;
        RECT 273.650 190.330 278.490 195.060 ;
        RECT 299.650 190.330 304.490 195.060 ;
        RECT 39.650 180.330 44.490 185.060 ;
        RECT 65.650 180.330 70.490 185.060 ;
        RECT 91.650 180.330 96.490 185.060 ;
        RECT 117.650 180.330 122.490 185.060 ;
        RECT 143.650 180.330 148.490 185.060 ;
        RECT 169.650 180.330 174.490 185.060 ;
        RECT 195.650 180.330 200.490 185.060 ;
        RECT 221.650 180.330 226.490 185.060 ;
        RECT 247.650 180.330 252.490 185.060 ;
        RECT 273.650 180.330 278.490 185.060 ;
        RECT 299.650 180.330 304.490 185.060 ;
        RECT 39.650 170.330 44.490 175.060 ;
        RECT 65.650 170.330 70.490 175.060 ;
        RECT 91.650 170.330 96.490 175.060 ;
        RECT 117.650 170.330 122.490 175.060 ;
        RECT 143.650 170.330 148.490 175.060 ;
        RECT 169.650 170.330 174.490 175.060 ;
        RECT 195.650 170.330 200.490 175.060 ;
        RECT 221.650 170.330 226.490 175.060 ;
        RECT 247.650 170.330 252.490 175.060 ;
        RECT 273.650 170.330 278.490 175.060 ;
        RECT 299.650 170.330 304.490 175.060 ;
        RECT 49.460 72.350 51.760 74.800 ;
        RECT 110.890 74.790 112.970 104.780 ;
        RECT 148.320 102.715 149.850 104.600 ;
        RECT 234.210 104.200 236.500 104.750 ;
        RECT 234.930 103.850 235.260 104.200 ;
        RECT 234.930 103.510 239.380 103.850 ;
        RECT 234.210 102.090 236.510 103.130 ;
        RECT 239.060 102.090 239.380 103.510 ;
        RECT 234.210 101.770 239.420 102.090 ;
        RECT 234.210 101.000 236.510 101.770 ;
        RECT 239.090 88.070 239.420 101.770 ;
        RECT 281.620 98.310 283.890 98.360 ;
        RECT 292.860 98.310 293.170 98.320 ;
        RECT 281.620 97.930 293.470 98.310 ;
        RECT 281.620 97.880 283.890 97.930 ;
        RECT 213.840 85.510 216.410 87.680 ;
        RECT 238.280 85.900 240.850 88.070 ;
        RECT 264.840 84.840 267.410 87.010 ;
        RECT 292.860 86.720 293.170 97.930 ;
        RECT 292.020 84.550 294.590 86.720 ;
        RECT 148.120 82.070 149.540 84.150 ;
        RECT 148.120 81.040 149.590 82.070 ;
        RECT 148.170 76.860 149.590 81.040 ;
        RECT 85.310 73.310 86.500 74.670 ;
        RECT 147.820 74.460 149.740 76.860 ;
        RECT 193.000 58.750 194.190 60.110 ;
        RECT 219.250 56.920 233.170 61.120 ;
        RECT 147.305 50.060 148.840 50.115 ;
        RECT 110.820 48.930 148.840 50.060 ;
        RECT 85.020 46.560 86.210 47.920 ;
        RECT 111.040 47.315 112.790 48.930 ;
        RECT 147.305 48.150 148.840 48.930 ;
        RECT 110.960 45.685 112.790 47.315 ;
        RECT 111.040 45.390 112.790 45.685 ;
        RECT 284.240 26.940 284.580 28.350 ;
        RECT 283.750 26.630 284.580 26.940 ;
        RECT 249.520 26.440 270.650 26.450 ;
        RECT 249.520 26.020 270.660 26.440 ;
        RECT 119.140 24.650 120.240 25.960 ;
        RECT 249.530 24.850 249.870 26.020 ;
        RECT 119.120 21.220 120.240 24.650 ;
        RECT 242.670 24.200 244.760 24.740 ;
        RECT 249.470 24.620 249.870 24.850 ;
        RECT 270.310 25.520 270.660 26.020 ;
        RECT 249.470 24.230 249.850 24.620 ;
        RECT 249.230 24.200 249.850 24.230 ;
        RECT 242.670 23.840 249.850 24.200 ;
        RECT 270.310 23.850 270.730 25.520 ;
        RECT 242.670 23.820 245.310 23.840 ;
        RECT 242.670 22.670 244.760 23.820 ;
        RECT 270.330 23.810 270.730 23.850 ;
        RECT 270.330 23.400 270.680 23.810 ;
        RECT 275.260 23.450 275.620 25.480 ;
        RECT 283.750 25.180 284.130 26.630 ;
        RECT 283.730 23.740 284.130 25.180 ;
        RECT 275.170 23.410 281.200 23.450 ;
        RECT 283.710 23.410 284.130 23.740 ;
        RECT 270.330 23.390 272.930 23.400 ;
        RECT 275.170 23.390 284.130 23.410 ;
        RECT 270.330 23.070 284.130 23.390 ;
        RECT 270.800 23.050 272.930 23.070 ;
        RECT 275.170 23.050 284.130 23.070 ;
        RECT 280.570 23.030 284.130 23.050 ;
        RECT 283.710 23.020 284.130 23.030 ;
        RECT 119.090 18.370 120.490 19.540 ;
        RECT 694.810 6.790 720.310 8.590 ;
      LAYER via3 ;
        RECT 40.380 323.190 43.810 326.180 ;
        RECT 66.380 323.190 69.810 326.180 ;
        RECT 92.380 323.190 95.810 326.180 ;
        RECT 118.380 323.190 121.810 326.180 ;
        RECT 144.380 323.190 147.810 326.180 ;
        RECT 170.380 323.190 173.810 326.180 ;
        RECT 196.380 323.190 199.810 326.180 ;
        RECT 222.380 323.190 225.810 326.180 ;
        RECT 248.380 323.190 251.810 326.180 ;
        RECT 274.380 323.190 277.810 326.180 ;
        RECT 300.380 323.190 303.810 326.180 ;
        RECT 40.380 313.190 43.810 316.180 ;
        RECT 66.380 313.190 69.810 316.180 ;
        RECT 92.380 313.190 95.810 316.180 ;
        RECT 118.380 313.190 121.810 316.180 ;
        RECT 144.380 313.190 147.810 316.180 ;
        RECT 170.380 313.190 173.810 316.180 ;
        RECT 196.380 313.190 199.810 316.180 ;
        RECT 222.380 313.190 225.810 316.180 ;
        RECT 248.380 313.190 251.810 316.180 ;
        RECT 274.380 313.190 277.810 316.180 ;
        RECT 300.380 313.190 303.810 316.180 ;
        RECT 40.380 303.190 43.810 306.180 ;
        RECT 66.380 303.190 69.810 306.180 ;
        RECT 92.380 303.190 95.810 306.180 ;
        RECT 118.380 303.190 121.810 306.180 ;
        RECT 144.380 303.190 147.810 306.180 ;
        RECT 170.380 303.190 173.810 306.180 ;
        RECT 196.380 303.190 199.810 306.180 ;
        RECT 222.380 303.190 225.810 306.180 ;
        RECT 248.380 303.190 251.810 306.180 ;
        RECT 274.380 303.190 277.810 306.180 ;
        RECT 300.380 303.190 303.810 306.180 ;
        RECT 40.380 293.190 43.810 296.180 ;
        RECT 66.380 293.190 69.810 296.180 ;
        RECT 92.380 293.190 95.810 296.180 ;
        RECT 118.380 293.190 121.810 296.180 ;
        RECT 144.380 293.190 147.810 296.180 ;
        RECT 170.380 293.190 173.810 296.180 ;
        RECT 196.380 293.190 199.810 296.180 ;
        RECT 222.380 293.190 225.810 296.180 ;
        RECT 248.380 293.190 251.810 296.180 ;
        RECT 274.380 293.190 277.810 296.180 ;
        RECT 300.380 293.190 303.810 296.180 ;
        RECT 40.380 283.190 43.810 286.180 ;
        RECT 66.380 283.190 69.810 286.180 ;
        RECT 92.380 283.190 95.810 286.180 ;
        RECT 118.380 283.190 121.810 286.180 ;
        RECT 144.380 283.190 147.810 286.180 ;
        RECT 170.380 283.190 173.810 286.180 ;
        RECT 196.380 283.190 199.810 286.180 ;
        RECT 222.380 283.190 225.810 286.180 ;
        RECT 248.380 283.190 251.810 286.180 ;
        RECT 274.380 283.190 277.810 286.180 ;
        RECT 300.380 283.190 303.810 286.180 ;
        RECT 40.380 273.190 43.810 276.180 ;
        RECT 66.380 273.190 69.810 276.180 ;
        RECT 92.380 273.190 95.810 276.180 ;
        RECT 118.380 273.190 121.810 276.180 ;
        RECT 144.380 273.190 147.810 276.180 ;
        RECT 170.380 273.190 173.810 276.180 ;
        RECT 196.380 273.190 199.810 276.180 ;
        RECT 222.380 273.190 225.810 276.180 ;
        RECT 248.380 273.190 251.810 276.180 ;
        RECT 274.380 273.190 277.810 276.180 ;
        RECT 300.380 273.190 303.810 276.180 ;
        RECT 40.380 263.190 43.810 266.180 ;
        RECT 66.380 263.190 69.810 266.180 ;
        RECT 92.380 263.190 95.810 266.180 ;
        RECT 118.380 263.190 121.810 266.180 ;
        RECT 144.380 263.190 147.810 266.180 ;
        RECT 170.380 263.190 173.810 266.180 ;
        RECT 196.380 263.190 199.810 266.180 ;
        RECT 222.380 263.190 225.810 266.180 ;
        RECT 248.380 263.190 251.810 266.180 ;
        RECT 274.380 263.190 277.810 266.180 ;
        RECT 300.380 263.190 303.810 266.180 ;
        RECT 40.380 253.190 43.810 256.180 ;
        RECT 66.380 253.190 69.810 256.180 ;
        RECT 92.380 253.190 95.810 256.180 ;
        RECT 118.380 253.190 121.810 256.180 ;
        RECT 144.380 253.190 147.810 256.180 ;
        RECT 170.380 253.190 173.810 256.180 ;
        RECT 196.380 253.190 199.810 256.180 ;
        RECT 222.380 253.190 225.810 256.180 ;
        RECT 248.380 253.190 251.810 256.180 ;
        RECT 274.380 253.190 277.810 256.180 ;
        RECT 300.380 253.190 303.810 256.180 ;
        RECT 690.020 250.510 690.420 250.910 ;
        RECT 690.820 250.510 691.220 250.910 ;
        RECT 691.620 250.510 692.020 250.910 ;
        RECT 692.420 250.510 692.820 250.910 ;
        RECT 693.220 250.510 693.620 250.910 ;
        RECT 694.020 250.510 694.420 250.910 ;
        RECT 694.820 250.510 695.220 250.910 ;
        RECT 695.620 250.510 696.020 250.910 ;
        RECT 696.420 250.510 696.820 250.910 ;
        RECT 697.220 250.510 697.620 250.910 ;
        RECT 698.020 250.510 698.420 250.910 ;
        RECT 698.820 250.510 699.220 250.910 ;
        RECT 699.620 250.510 700.020 250.910 ;
        RECT 700.420 250.510 700.820 250.910 ;
        RECT 701.220 250.510 701.620 250.910 ;
        RECT 702.020 250.510 702.420 250.910 ;
        RECT 702.820 250.510 703.220 250.910 ;
        RECT 703.620 250.510 704.020 250.910 ;
        RECT 704.420 250.510 704.820 250.910 ;
        RECT 705.220 250.510 705.620 250.910 ;
        RECT 706.020 250.510 706.420 250.910 ;
        RECT 706.820 250.510 707.220 250.910 ;
        RECT 707.620 250.510 708.020 250.910 ;
        RECT 708.420 250.510 708.820 250.910 ;
        RECT 709.220 250.510 709.620 250.910 ;
        RECT 710.020 250.510 710.420 250.910 ;
        RECT 710.820 250.510 711.220 250.910 ;
        RECT 711.620 250.510 712.020 250.910 ;
        RECT 712.420 250.510 712.820 250.910 ;
        RECT 713.220 250.510 713.620 250.910 ;
        RECT 714.020 250.510 714.420 250.910 ;
        RECT 690.020 249.710 690.420 250.110 ;
        RECT 690.820 249.710 691.220 250.110 ;
        RECT 691.620 249.710 692.020 250.110 ;
        RECT 692.420 249.710 692.820 250.110 ;
        RECT 693.220 249.710 693.620 250.110 ;
        RECT 694.020 249.710 694.420 250.110 ;
        RECT 694.820 249.710 695.220 250.110 ;
        RECT 695.620 249.710 696.020 250.110 ;
        RECT 696.420 249.710 696.820 250.110 ;
        RECT 697.220 249.710 697.620 250.110 ;
        RECT 698.020 249.710 698.420 250.110 ;
        RECT 698.820 249.710 699.220 250.110 ;
        RECT 699.620 249.710 700.020 250.110 ;
        RECT 700.420 249.710 700.820 250.110 ;
        RECT 701.220 249.710 701.620 250.110 ;
        RECT 702.020 249.710 702.420 250.110 ;
        RECT 702.820 249.710 703.220 250.110 ;
        RECT 703.620 249.710 704.020 250.110 ;
        RECT 704.420 249.710 704.820 250.110 ;
        RECT 705.220 249.710 705.620 250.110 ;
        RECT 706.020 249.710 706.420 250.110 ;
        RECT 706.820 249.710 707.220 250.110 ;
        RECT 707.620 249.710 708.020 250.110 ;
        RECT 708.420 249.710 708.820 250.110 ;
        RECT 709.220 249.710 709.620 250.110 ;
        RECT 710.020 249.710 710.420 250.110 ;
        RECT 710.820 249.710 711.220 250.110 ;
        RECT 711.620 249.710 712.020 250.110 ;
        RECT 712.420 249.710 712.820 250.110 ;
        RECT 713.220 249.710 713.620 250.110 ;
        RECT 714.020 249.710 714.420 250.110 ;
        RECT 40.380 241.190 43.810 244.180 ;
        RECT 66.380 241.190 69.810 244.180 ;
        RECT 92.380 241.190 95.810 244.180 ;
        RECT 118.380 241.190 121.810 244.180 ;
        RECT 144.380 241.190 147.810 244.180 ;
        RECT 170.380 241.190 173.810 244.180 ;
        RECT 196.380 241.190 199.810 244.180 ;
        RECT 222.380 241.190 225.810 244.180 ;
        RECT 248.380 241.190 251.810 244.180 ;
        RECT 274.380 241.190 277.810 244.180 ;
        RECT 300.380 241.190 303.810 244.180 ;
        RECT 40.380 231.190 43.810 234.180 ;
        RECT 66.380 231.190 69.810 234.180 ;
        RECT 92.380 231.190 95.810 234.180 ;
        RECT 118.380 231.190 121.810 234.180 ;
        RECT 144.380 231.190 147.810 234.180 ;
        RECT 170.380 231.190 173.810 234.180 ;
        RECT 196.380 231.190 199.810 234.180 ;
        RECT 222.380 231.190 225.810 234.180 ;
        RECT 248.380 231.190 251.810 234.180 ;
        RECT 274.380 231.190 277.810 234.180 ;
        RECT 300.380 231.190 303.810 234.180 ;
        RECT 40.380 221.190 43.810 224.180 ;
        RECT 66.380 221.190 69.810 224.180 ;
        RECT 92.380 221.190 95.810 224.180 ;
        RECT 118.380 221.190 121.810 224.180 ;
        RECT 144.380 221.190 147.810 224.180 ;
        RECT 170.380 221.190 173.810 224.180 ;
        RECT 196.380 221.190 199.810 224.180 ;
        RECT 222.380 221.190 225.810 224.180 ;
        RECT 248.380 221.190 251.810 224.180 ;
        RECT 274.380 221.190 277.810 224.180 ;
        RECT 300.380 221.190 303.810 224.180 ;
        RECT 40.380 211.190 43.810 214.180 ;
        RECT 66.380 211.190 69.810 214.180 ;
        RECT 92.380 211.190 95.810 214.180 ;
        RECT 118.380 211.190 121.810 214.180 ;
        RECT 144.380 211.190 147.810 214.180 ;
        RECT 170.380 211.190 173.810 214.180 ;
        RECT 196.380 211.190 199.810 214.180 ;
        RECT 222.380 211.190 225.810 214.180 ;
        RECT 248.380 211.190 251.810 214.180 ;
        RECT 274.380 211.190 277.810 214.180 ;
        RECT 300.380 211.190 303.810 214.180 ;
        RECT 40.380 201.190 43.810 204.180 ;
        RECT 66.380 201.190 69.810 204.180 ;
        RECT 92.380 201.190 95.810 204.180 ;
        RECT 118.380 201.190 121.810 204.180 ;
        RECT 144.380 201.190 147.810 204.180 ;
        RECT 170.380 201.190 173.810 204.180 ;
        RECT 196.380 201.190 199.810 204.180 ;
        RECT 222.380 201.190 225.810 204.180 ;
        RECT 248.380 201.190 251.810 204.180 ;
        RECT 274.380 201.190 277.810 204.180 ;
        RECT 300.380 201.190 303.810 204.180 ;
        RECT 40.380 191.190 43.810 194.180 ;
        RECT 66.380 191.190 69.810 194.180 ;
        RECT 92.380 191.190 95.810 194.180 ;
        RECT 118.380 191.190 121.810 194.180 ;
        RECT 144.380 191.190 147.810 194.180 ;
        RECT 170.380 191.190 173.810 194.180 ;
        RECT 196.380 191.190 199.810 194.180 ;
        RECT 222.380 191.190 225.810 194.180 ;
        RECT 248.380 191.190 251.810 194.180 ;
        RECT 274.380 191.190 277.810 194.180 ;
        RECT 300.380 191.190 303.810 194.180 ;
        RECT 40.380 181.190 43.810 184.180 ;
        RECT 66.380 181.190 69.810 184.180 ;
        RECT 92.380 181.190 95.810 184.180 ;
        RECT 118.380 181.190 121.810 184.180 ;
        RECT 144.380 181.190 147.810 184.180 ;
        RECT 170.380 181.190 173.810 184.180 ;
        RECT 196.380 181.190 199.810 184.180 ;
        RECT 222.380 181.190 225.810 184.180 ;
        RECT 248.380 181.190 251.810 184.180 ;
        RECT 274.380 181.190 277.810 184.180 ;
        RECT 300.380 181.190 303.810 184.180 ;
        RECT 40.380 171.190 43.810 174.180 ;
        RECT 66.380 171.190 69.810 174.180 ;
        RECT 92.380 171.190 95.810 174.180 ;
        RECT 118.380 171.190 121.810 174.180 ;
        RECT 144.380 171.190 147.810 174.180 ;
        RECT 170.380 171.190 173.810 174.180 ;
        RECT 196.380 171.190 199.810 174.180 ;
        RECT 222.380 171.190 225.810 174.180 ;
        RECT 248.380 171.190 251.810 174.180 ;
        RECT 274.380 171.190 277.810 174.180 ;
        RECT 300.380 171.190 303.810 174.180 ;
        RECT 111.360 102.970 112.555 104.535 ;
        RECT 148.410 102.775 149.775 104.525 ;
        RECT 214.310 86.000 215.940 87.200 ;
        RECT 238.750 86.390 240.380 87.590 ;
        RECT 265.310 85.330 266.940 86.530 ;
        RECT 292.490 85.040 294.120 86.240 ;
        RECT 148.350 83.330 149.400 83.960 ;
        RECT 111.305 75.180 112.220 76.705 ;
        RECT 148.340 75.070 149.310 76.610 ;
        RECT 49.610 72.640 51.570 74.640 ;
        RECT 193.150 58.970 194.030 59.860 ;
        RECT 220.320 58.080 223.210 60.090 ;
        RECT 230.400 58.170 232.900 60.140 ;
        RECT 119.820 49.380 120.550 49.980 ;
        RECT 85.170 46.780 86.050 47.670 ;
        RECT 147.500 48.250 148.730 49.995 ;
        RECT 111.110 45.880 112.015 47.160 ;
        RECT 119.480 24.890 119.920 25.460 ;
        RECT 242.950 22.900 244.460 24.580 ;
        RECT 119.300 21.460 120.040 22.100 ;
        RECT 119.420 18.640 120.280 19.270 ;
        RECT 695.310 7.790 695.710 8.190 ;
        RECT 696.110 7.790 696.510 8.190 ;
        RECT 696.910 7.790 697.310 8.190 ;
        RECT 697.710 7.790 698.110 8.190 ;
        RECT 698.510 7.790 698.910 8.190 ;
        RECT 699.310 7.790 699.710 8.190 ;
        RECT 700.110 7.790 700.510 8.190 ;
        RECT 700.910 7.790 701.310 8.190 ;
        RECT 701.710 7.790 702.110 8.190 ;
        RECT 702.510 7.790 702.910 8.190 ;
        RECT 703.310 7.790 703.710 8.190 ;
        RECT 704.110 7.790 704.510 8.190 ;
        RECT 704.910 7.790 705.310 8.190 ;
        RECT 705.710 7.790 706.110 8.190 ;
        RECT 706.510 7.790 706.910 8.190 ;
        RECT 707.310 7.790 707.710 8.190 ;
        RECT 708.110 7.790 708.510 8.190 ;
        RECT 708.910 7.790 709.310 8.190 ;
        RECT 709.710 7.790 710.110 8.190 ;
        RECT 710.510 7.790 710.910 8.190 ;
        RECT 711.310 7.790 711.710 8.190 ;
        RECT 712.110 7.790 712.510 8.190 ;
        RECT 712.910 7.790 713.310 8.190 ;
        RECT 713.710 7.790 714.110 8.190 ;
        RECT 714.510 7.790 714.910 8.190 ;
        RECT 715.310 7.790 715.710 8.190 ;
        RECT 716.110 7.790 716.510 8.190 ;
        RECT 716.910 7.790 717.310 8.190 ;
        RECT 717.710 7.790 718.110 8.190 ;
        RECT 718.510 7.790 718.910 8.190 ;
        RECT 719.310 7.790 719.710 8.190 ;
        RECT 695.310 6.990 695.710 7.390 ;
        RECT 696.110 6.990 696.510 7.390 ;
        RECT 696.910 6.990 697.310 7.390 ;
        RECT 697.710 6.990 698.110 7.390 ;
        RECT 698.510 6.990 698.910 7.390 ;
        RECT 699.310 6.990 699.710 7.390 ;
        RECT 700.110 6.990 700.510 7.390 ;
        RECT 700.910 6.990 701.310 7.390 ;
        RECT 701.710 6.990 702.110 7.390 ;
        RECT 702.510 6.990 702.910 7.390 ;
        RECT 703.310 6.990 703.710 7.390 ;
        RECT 704.110 6.990 704.510 7.390 ;
        RECT 704.910 6.990 705.310 7.390 ;
        RECT 705.710 6.990 706.110 7.390 ;
        RECT 706.510 6.990 706.910 7.390 ;
        RECT 707.310 6.990 707.710 7.390 ;
        RECT 708.110 6.990 708.510 7.390 ;
        RECT 708.910 6.990 709.310 7.390 ;
        RECT 709.710 6.990 710.110 7.390 ;
        RECT 710.510 6.990 710.910 7.390 ;
        RECT 711.310 6.990 711.710 7.390 ;
        RECT 712.110 6.990 712.510 7.390 ;
        RECT 712.910 6.990 713.310 7.390 ;
        RECT 713.710 6.990 714.110 7.390 ;
        RECT 714.510 6.990 714.910 7.390 ;
        RECT 715.310 6.990 715.710 7.390 ;
        RECT 716.110 6.990 716.510 7.390 ;
        RECT 716.910 6.990 717.310 7.390 ;
        RECT 717.710 6.990 718.110 7.390 ;
        RECT 718.510 6.990 718.910 7.390 ;
        RECT 719.310 6.990 719.710 7.390 ;
      LAYER met4 ;
        RECT 673.820 394.390 726.660 394.880 ;
        RECT -33.940 391.530 -17.650 391.620 ;
        RECT 667.260 391.550 726.660 394.390 ;
        RECT -12.400 391.530 726.660 391.550 ;
        RECT -33.940 375.370 726.660 391.530 ;
        RECT -33.940 372.040 726.220 375.370 ;
        RECT -33.940 372.010 -6.560 372.040 ;
        RECT -33.940 -3.880 -17.650 372.010 ;
        RECT 299.510 327.060 304.210 372.040 ;
        RECT 667.260 371.900 726.220 372.040 ;
        RECT 39.650 322.330 44.490 327.060 ;
        RECT 65.650 322.330 70.490 327.060 ;
        RECT 91.650 322.330 96.490 327.060 ;
        RECT 117.650 322.330 122.490 327.060 ;
        RECT 143.650 322.330 148.490 327.060 ;
        RECT 169.650 322.330 174.490 327.060 ;
        RECT 195.650 322.330 200.490 327.060 ;
        RECT 221.650 322.330 226.490 327.060 ;
        RECT 247.650 322.330 252.490 327.060 ;
        RECT 273.650 322.330 278.490 327.060 ;
        RECT 299.510 322.330 304.490 327.060 ;
        RECT 299.510 321.080 304.210 322.330 ;
        RECT 39.650 312.330 44.490 317.060 ;
        RECT 65.650 312.330 70.490 317.060 ;
        RECT 91.650 312.330 96.490 317.060 ;
        RECT 117.650 312.330 122.490 317.060 ;
        RECT 143.650 312.330 148.490 317.060 ;
        RECT 169.650 312.330 174.490 317.060 ;
        RECT 195.650 312.330 200.490 317.060 ;
        RECT 221.650 312.330 226.490 317.060 ;
        RECT 247.650 312.330 252.490 317.060 ;
        RECT 273.650 312.330 278.490 317.060 ;
        RECT 299.650 312.330 304.490 317.060 ;
        RECT 39.650 302.330 44.490 307.060 ;
        RECT 65.650 302.330 70.490 307.060 ;
        RECT 91.650 302.330 96.490 307.060 ;
        RECT 117.650 302.330 122.490 307.060 ;
        RECT 143.650 302.330 148.490 307.060 ;
        RECT 169.650 302.330 174.490 307.060 ;
        RECT 195.650 302.330 200.490 307.060 ;
        RECT 221.650 302.330 226.490 307.060 ;
        RECT 247.650 302.330 252.490 307.060 ;
        RECT 273.650 302.330 278.490 307.060 ;
        RECT 299.650 302.330 304.490 307.060 ;
        RECT 39.650 292.330 44.490 297.060 ;
        RECT 65.650 292.330 70.490 297.060 ;
        RECT 91.650 292.330 96.490 297.060 ;
        RECT 117.650 292.330 122.490 297.060 ;
        RECT 143.650 292.330 148.490 297.060 ;
        RECT 169.650 292.330 174.490 297.060 ;
        RECT 195.650 292.330 200.490 297.060 ;
        RECT 221.650 292.330 226.490 297.060 ;
        RECT 247.650 292.330 252.490 297.060 ;
        RECT 273.650 292.330 278.490 297.060 ;
        RECT 299.650 292.330 304.490 297.060 ;
        RECT 39.650 282.330 44.490 287.060 ;
        RECT 65.650 282.330 70.490 287.060 ;
        RECT 91.650 282.330 96.490 287.060 ;
        RECT 117.650 282.330 122.490 287.060 ;
        RECT 143.650 282.330 148.490 287.060 ;
        RECT 169.650 282.330 174.490 287.060 ;
        RECT 195.650 282.330 200.490 287.060 ;
        RECT 221.650 282.330 226.490 287.060 ;
        RECT 247.650 282.330 252.490 287.060 ;
        RECT 273.650 282.330 278.490 287.060 ;
        RECT 299.650 282.330 304.490 287.060 ;
        RECT 39.650 272.330 44.490 277.060 ;
        RECT 65.650 272.330 70.490 277.060 ;
        RECT 91.650 272.330 96.490 277.060 ;
        RECT 117.650 272.330 122.490 277.060 ;
        RECT 143.650 272.330 148.490 277.060 ;
        RECT 169.650 272.330 174.490 277.060 ;
        RECT 195.650 272.330 200.490 277.060 ;
        RECT 221.650 272.330 226.490 277.060 ;
        RECT 247.650 272.330 252.490 277.060 ;
        RECT 273.650 272.330 278.490 277.060 ;
        RECT 299.650 272.330 304.490 277.060 ;
        RECT 39.650 262.330 44.490 267.060 ;
        RECT 65.650 262.330 70.490 267.060 ;
        RECT 91.650 262.330 96.490 267.060 ;
        RECT 117.650 262.330 122.490 267.060 ;
        RECT 143.650 262.330 148.490 267.060 ;
        RECT 169.650 262.330 174.490 267.060 ;
        RECT 195.650 262.330 200.490 267.060 ;
        RECT 221.650 262.330 226.490 267.060 ;
        RECT 247.650 262.330 252.490 267.060 ;
        RECT 273.650 262.330 278.490 267.060 ;
        RECT 299.650 262.330 304.490 267.060 ;
        RECT 39.650 252.330 44.490 257.060 ;
        RECT 65.650 252.330 70.490 257.060 ;
        RECT 91.650 252.330 96.490 257.060 ;
        RECT 117.650 252.330 122.490 257.060 ;
        RECT 143.650 252.330 148.490 257.060 ;
        RECT 169.650 252.330 174.490 257.060 ;
        RECT 195.650 252.330 200.490 257.060 ;
        RECT 221.650 252.330 226.490 257.060 ;
        RECT 247.650 252.330 252.490 257.060 ;
        RECT 273.650 252.330 278.490 257.060 ;
        RECT 299.650 252.330 304.490 257.060 ;
        RECT 39.650 240.330 44.490 245.060 ;
        RECT 65.650 240.330 70.490 245.060 ;
        RECT 91.650 240.330 96.490 245.060 ;
        RECT 117.650 240.330 122.490 245.060 ;
        RECT 143.650 240.330 148.490 245.060 ;
        RECT 169.650 240.330 174.490 245.060 ;
        RECT 195.650 240.330 200.490 245.060 ;
        RECT 221.650 240.330 226.490 245.060 ;
        RECT 247.650 240.330 252.490 245.060 ;
        RECT 273.650 240.330 278.490 245.060 ;
        RECT 299.650 240.330 304.490 245.060 ;
        RECT 39.650 230.330 44.490 235.060 ;
        RECT 65.650 230.330 70.490 235.060 ;
        RECT 91.650 230.330 96.490 235.060 ;
        RECT 117.650 230.330 122.490 235.060 ;
        RECT 143.650 230.330 148.490 235.060 ;
        RECT 169.650 230.330 174.490 235.060 ;
        RECT 195.650 230.330 200.490 235.060 ;
        RECT 221.650 230.330 226.490 235.060 ;
        RECT 247.650 230.330 252.490 235.060 ;
        RECT 273.650 230.330 278.490 235.060 ;
        RECT 299.650 230.330 304.490 235.060 ;
        RECT 39.650 220.330 44.490 225.060 ;
        RECT 65.650 220.330 70.490 225.060 ;
        RECT 91.650 220.330 96.490 225.060 ;
        RECT 117.650 220.330 122.490 225.060 ;
        RECT 143.650 220.330 148.490 225.060 ;
        RECT 169.650 220.330 174.490 225.060 ;
        RECT 195.650 220.330 200.490 225.060 ;
        RECT 221.650 220.330 226.490 225.060 ;
        RECT 247.650 220.330 252.490 225.060 ;
        RECT 273.650 220.330 278.490 225.060 ;
        RECT 299.650 220.330 304.490 225.060 ;
        RECT 39.650 210.330 44.490 215.060 ;
        RECT 65.650 210.330 70.490 215.060 ;
        RECT 91.650 210.330 96.490 215.060 ;
        RECT 117.650 210.330 122.490 215.060 ;
        RECT 143.650 210.330 148.490 215.060 ;
        RECT 169.650 210.330 174.490 215.060 ;
        RECT 195.650 210.330 200.490 215.060 ;
        RECT 221.650 210.330 226.490 215.060 ;
        RECT 247.650 210.330 252.490 215.060 ;
        RECT 273.650 210.330 278.490 215.060 ;
        RECT 299.650 210.330 304.490 215.060 ;
        RECT 39.650 200.330 44.490 205.060 ;
        RECT 65.650 200.330 70.490 205.060 ;
        RECT 91.650 200.330 96.490 205.060 ;
        RECT 117.650 200.330 122.490 205.060 ;
        RECT 143.650 200.330 148.490 205.060 ;
        RECT 169.650 200.330 174.490 205.060 ;
        RECT 195.650 200.330 200.490 205.060 ;
        RECT 221.650 200.330 226.490 205.060 ;
        RECT 247.650 200.330 252.490 205.060 ;
        RECT 273.650 200.330 278.490 205.060 ;
        RECT 299.650 200.330 304.490 205.060 ;
        RECT 39.650 190.330 44.490 195.060 ;
        RECT 65.650 190.330 70.490 195.060 ;
        RECT 91.650 190.330 96.490 195.060 ;
        RECT 117.650 190.330 122.490 195.060 ;
        RECT 143.650 190.330 148.490 195.060 ;
        RECT 169.650 190.330 174.490 195.060 ;
        RECT 195.650 190.330 200.490 195.060 ;
        RECT 221.650 190.330 226.490 195.060 ;
        RECT 247.650 190.330 252.490 195.060 ;
        RECT 273.650 190.330 278.490 195.060 ;
        RECT 299.650 190.330 304.490 195.060 ;
        RECT 39.650 180.330 44.490 185.060 ;
        RECT 65.650 180.330 70.490 185.060 ;
        RECT 91.650 180.330 96.490 185.060 ;
        RECT 117.650 180.330 122.490 185.060 ;
        RECT 143.650 180.330 148.490 185.060 ;
        RECT 169.650 180.330 174.490 185.060 ;
        RECT 195.650 180.330 200.490 185.060 ;
        RECT 221.650 180.330 226.490 185.060 ;
        RECT 247.650 180.330 252.490 185.060 ;
        RECT 273.650 180.330 278.490 185.060 ;
        RECT 299.650 180.330 304.490 185.060 ;
        RECT 169.320 175.060 174.360 175.560 ;
        RECT 39.650 170.330 44.490 175.060 ;
        RECT 65.650 170.330 70.490 175.060 ;
        RECT 91.650 170.330 96.490 175.060 ;
        RECT 117.650 170.330 122.490 175.060 ;
        RECT 143.650 170.330 148.490 175.060 ;
        RECT 169.320 170.330 174.490 175.060 ;
        RECT 195.650 170.330 200.490 175.060 ;
        RECT 221.650 170.330 226.490 175.060 ;
        RECT 247.650 170.330 252.490 175.060 ;
        RECT 273.650 170.330 278.490 175.060 ;
        RECT 299.650 170.330 304.490 175.060 ;
        RECT 169.320 165.770 174.360 170.330 ;
        RECT 169.170 163.160 295.830 165.770 ;
        RECT 291.030 151.540 295.830 163.160 ;
        RECT 111.270 102.875 112.660 104.630 ;
        RECT 148.020 93.000 150.050 105.170 ;
        RECT 150.910 93.000 154.980 93.030 ;
        RECT 147.990 92.900 177.800 93.000 ;
        RECT 147.990 92.490 194.020 92.900 ;
        RECT 147.990 91.510 194.030 92.490 ;
        RECT 148.020 84.100 149.650 91.510 ;
        RECT 150.910 91.460 154.980 91.510 ;
        RECT 174.230 90.980 194.030 91.510 ;
        RECT 192.800 87.580 194.030 90.980 ;
        RECT 192.410 87.360 195.860 87.580 ;
        RECT 192.410 87.280 211.010 87.360 ;
        RECT 213.840 87.280 216.410 87.680 ;
        RECT 238.280 87.280 240.850 88.070 ;
        RECT 291.280 87.280 294.960 151.540 ;
        RECT 192.410 85.140 295.580 87.280 ;
        RECT 148.000 83.100 149.740 84.100 ;
        RECT 110.290 76.960 113.370 77.060 ;
        RECT 49.460 72.350 51.760 74.800 ;
        RECT 110.290 52.030 113.540 76.960 ;
        RECT 147.820 74.460 149.740 76.860 ;
        RECT 110.290 48.870 113.480 52.030 ;
        RECT 147.890 51.040 149.170 74.460 ;
        RECT 192.410 60.200 195.860 85.140 ;
        RECT 209.800 85.130 295.580 85.140 ;
        RECT 264.840 84.840 267.410 85.130 ;
        RECT 291.280 84.220 294.960 85.130 ;
        RECT 204.030 60.200 224.890 60.370 ;
        RECT 192.250 59.510 224.890 60.200 ;
        RECT 192.250 58.130 224.950 59.510 ;
        RECT 204.090 58.020 224.950 58.130 ;
        RECT 229.600 57.640 245.310 60.940 ;
        RECT 84.370 48.380 113.480 48.870 ;
        RECT 84.370 47.780 113.540 48.380 ;
        RECT 84.370 45.560 113.560 47.780 ;
        RECT 119.150 47.310 120.790 50.290 ;
        RECT 146.900 50.280 149.390 51.040 ;
        RECT 147.050 49.980 149.170 50.280 ;
        RECT 147.050 48.070 149.000 49.980 ;
        RECT 242.190 49.450 244.950 57.640 ;
        RECT 84.370 45.500 113.540 45.560 ;
        RECT 110.290 45.180 113.540 45.500 ;
        RECT 119.170 45.370 120.790 47.310 ;
        RECT 242.190 46.600 245.320 49.450 ;
        RECT 119.140 24.710 120.790 45.370 ;
        RECT 242.620 22.710 245.320 46.600 ;
        RECT 242.670 22.670 244.760 22.710 ;
        RECT 118.940 19.820 120.590 22.510 ;
        RECT 118.940 18.640 120.600 19.820 ;
        RECT 118.940 18.230 120.590 18.640 ;
        RECT 682.890 -5.210 726.220 371.900 ;
    END
  END vdda1
  OBS
      LAYER pwell ;
        RECT 148.890 44.310 150.960 44.400 ;
        RECT 148.890 44.290 153.110 44.310 ;
      LAYER li1 ;
        RECT 46.770 330.955 54.770 331.125 ;
        RECT 55.060 330.955 63.060 331.125 ;
        RECT 72.770 330.955 80.770 331.125 ;
        RECT 81.060 330.955 89.060 331.125 ;
        RECT 98.770 330.955 106.770 331.125 ;
        RECT 107.060 330.955 115.060 331.125 ;
        RECT 124.770 330.955 132.770 331.125 ;
        RECT 133.060 330.955 141.060 331.125 ;
        RECT 150.770 330.955 158.770 331.125 ;
        RECT 159.060 330.955 167.060 331.125 ;
        RECT 176.770 330.955 184.770 331.125 ;
        RECT 185.060 330.955 193.060 331.125 ;
        RECT 202.770 330.955 210.770 331.125 ;
        RECT 211.060 330.955 219.060 331.125 ;
        RECT 228.770 330.955 236.770 331.125 ;
        RECT 237.060 330.955 245.060 331.125 ;
        RECT 254.770 330.955 262.770 331.125 ;
        RECT 263.060 330.955 271.060 331.125 ;
        RECT 280.770 330.955 288.770 331.125 ;
        RECT 289.060 330.955 297.060 331.125 ;
        RECT 46.770 323.315 54.770 323.485 ;
        RECT 55.060 323.315 63.060 323.485 ;
        RECT 72.770 323.315 80.770 323.485 ;
        RECT 81.060 323.315 89.060 323.485 ;
        RECT 98.770 323.315 106.770 323.485 ;
        RECT 107.060 323.315 115.060 323.485 ;
        RECT 124.770 323.315 132.770 323.485 ;
        RECT 133.060 323.315 141.060 323.485 ;
        RECT 150.770 323.315 158.770 323.485 ;
        RECT 159.060 323.315 167.060 323.485 ;
        RECT 176.770 323.315 184.770 323.485 ;
        RECT 185.060 323.315 193.060 323.485 ;
        RECT 202.770 323.315 210.770 323.485 ;
        RECT 211.060 323.315 219.060 323.485 ;
        RECT 228.770 323.315 236.770 323.485 ;
        RECT 237.060 323.315 245.060 323.485 ;
        RECT 254.770 323.315 262.770 323.485 ;
        RECT 263.060 323.315 271.060 323.485 ;
        RECT 280.770 323.315 288.770 323.485 ;
        RECT 289.060 323.315 297.060 323.485 ;
        RECT 46.770 322.775 54.770 322.945 ;
        RECT 55.060 322.775 63.060 322.945 ;
        RECT 72.770 322.775 80.770 322.945 ;
        RECT 81.060 322.775 89.060 322.945 ;
        RECT 98.770 322.775 106.770 322.945 ;
        RECT 107.060 322.775 115.060 322.945 ;
        RECT 124.770 322.775 132.770 322.945 ;
        RECT 133.060 322.775 141.060 322.945 ;
        RECT 150.770 322.775 158.770 322.945 ;
        RECT 159.060 322.775 167.060 322.945 ;
        RECT 176.770 322.775 184.770 322.945 ;
        RECT 185.060 322.775 193.060 322.945 ;
        RECT 202.770 322.775 210.770 322.945 ;
        RECT 211.060 322.775 219.060 322.945 ;
        RECT 228.770 322.775 236.770 322.945 ;
        RECT 237.060 322.775 245.060 322.945 ;
        RECT 254.770 322.775 262.770 322.945 ;
        RECT 263.060 322.775 271.060 322.945 ;
        RECT 280.770 322.775 288.770 322.945 ;
        RECT 289.060 322.775 297.060 322.945 ;
        RECT 46.770 315.135 54.770 315.305 ;
        RECT 55.060 315.135 63.060 315.305 ;
        RECT 72.770 315.135 80.770 315.305 ;
        RECT 81.060 315.135 89.060 315.305 ;
        RECT 98.770 315.135 106.770 315.305 ;
        RECT 107.060 315.135 115.060 315.305 ;
        RECT 124.770 315.135 132.770 315.305 ;
        RECT 133.060 315.135 141.060 315.305 ;
        RECT 150.770 315.135 158.770 315.305 ;
        RECT 159.060 315.135 167.060 315.305 ;
        RECT 176.770 315.135 184.770 315.305 ;
        RECT 185.060 315.135 193.060 315.305 ;
        RECT 202.770 315.135 210.770 315.305 ;
        RECT 211.060 315.135 219.060 315.305 ;
        RECT 228.770 315.135 236.770 315.305 ;
        RECT 237.060 315.135 245.060 315.305 ;
        RECT 254.770 315.135 262.770 315.305 ;
        RECT 263.060 315.135 271.060 315.305 ;
        RECT 280.770 315.135 288.770 315.305 ;
        RECT 289.060 315.135 297.060 315.305 ;
        RECT 46.770 314.595 54.770 314.765 ;
        RECT 55.060 314.595 63.060 314.765 ;
        RECT 72.770 314.595 80.770 314.765 ;
        RECT 81.060 314.595 89.060 314.765 ;
        RECT 98.770 314.595 106.770 314.765 ;
        RECT 107.060 314.595 115.060 314.765 ;
        RECT 124.770 314.595 132.770 314.765 ;
        RECT 133.060 314.595 141.060 314.765 ;
        RECT 150.770 314.595 158.770 314.765 ;
        RECT 159.060 314.595 167.060 314.765 ;
        RECT 176.770 314.595 184.770 314.765 ;
        RECT 185.060 314.595 193.060 314.765 ;
        RECT 202.770 314.595 210.770 314.765 ;
        RECT 211.060 314.595 219.060 314.765 ;
        RECT 228.770 314.595 236.770 314.765 ;
        RECT 237.060 314.595 245.060 314.765 ;
        RECT 254.770 314.595 262.770 314.765 ;
        RECT 263.060 314.595 271.060 314.765 ;
        RECT 280.770 314.595 288.770 314.765 ;
        RECT 289.060 314.595 297.060 314.765 ;
        RECT 46.770 306.955 54.770 307.125 ;
        RECT 55.060 306.955 63.060 307.125 ;
        RECT 72.770 306.955 80.770 307.125 ;
        RECT 81.060 306.955 89.060 307.125 ;
        RECT 98.770 306.955 106.770 307.125 ;
        RECT 107.060 306.955 115.060 307.125 ;
        RECT 124.770 306.955 132.770 307.125 ;
        RECT 133.060 306.955 141.060 307.125 ;
        RECT 150.770 306.955 158.770 307.125 ;
        RECT 159.060 306.955 167.060 307.125 ;
        RECT 176.770 306.955 184.770 307.125 ;
        RECT 185.060 306.955 193.060 307.125 ;
        RECT 202.770 306.955 210.770 307.125 ;
        RECT 211.060 306.955 219.060 307.125 ;
        RECT 228.770 306.955 236.770 307.125 ;
        RECT 237.060 306.955 245.060 307.125 ;
        RECT 254.770 306.955 262.770 307.125 ;
        RECT 263.060 306.955 271.060 307.125 ;
        RECT 280.770 306.955 288.770 307.125 ;
        RECT 289.060 306.955 297.060 307.125 ;
        RECT 46.770 306.415 54.770 306.585 ;
        RECT 55.060 306.415 63.060 306.585 ;
        RECT 72.770 306.415 80.770 306.585 ;
        RECT 81.060 306.415 89.060 306.585 ;
        RECT 98.770 306.415 106.770 306.585 ;
        RECT 107.060 306.415 115.060 306.585 ;
        RECT 124.770 306.415 132.770 306.585 ;
        RECT 133.060 306.415 141.060 306.585 ;
        RECT 150.770 306.415 158.770 306.585 ;
        RECT 159.060 306.415 167.060 306.585 ;
        RECT 176.770 306.415 184.770 306.585 ;
        RECT 185.060 306.415 193.060 306.585 ;
        RECT 202.770 306.415 210.770 306.585 ;
        RECT 211.060 306.415 219.060 306.585 ;
        RECT 228.770 306.415 236.770 306.585 ;
        RECT 237.060 306.415 245.060 306.585 ;
        RECT 254.770 306.415 262.770 306.585 ;
        RECT 263.060 306.415 271.060 306.585 ;
        RECT 280.770 306.415 288.770 306.585 ;
        RECT 289.060 306.415 297.060 306.585 ;
        RECT 46.770 298.775 54.770 298.945 ;
        RECT 55.060 298.775 63.060 298.945 ;
        RECT 72.770 298.775 80.770 298.945 ;
        RECT 81.060 298.775 89.060 298.945 ;
        RECT 98.770 298.775 106.770 298.945 ;
        RECT 107.060 298.775 115.060 298.945 ;
        RECT 124.770 298.775 132.770 298.945 ;
        RECT 133.060 298.775 141.060 298.945 ;
        RECT 150.770 298.775 158.770 298.945 ;
        RECT 159.060 298.775 167.060 298.945 ;
        RECT 176.770 298.775 184.770 298.945 ;
        RECT 185.060 298.775 193.060 298.945 ;
        RECT 202.770 298.775 210.770 298.945 ;
        RECT 211.060 298.775 219.060 298.945 ;
        RECT 228.770 298.775 236.770 298.945 ;
        RECT 237.060 298.775 245.060 298.945 ;
        RECT 254.770 298.775 262.770 298.945 ;
        RECT 263.060 298.775 271.060 298.945 ;
        RECT 280.770 298.775 288.770 298.945 ;
        RECT 289.060 298.775 297.060 298.945 ;
        RECT 46.770 298.235 54.770 298.405 ;
        RECT 55.060 298.235 63.060 298.405 ;
        RECT 72.770 298.235 80.770 298.405 ;
        RECT 81.060 298.235 89.060 298.405 ;
        RECT 98.770 298.235 106.770 298.405 ;
        RECT 107.060 298.235 115.060 298.405 ;
        RECT 124.770 298.235 132.770 298.405 ;
        RECT 133.060 298.235 141.060 298.405 ;
        RECT 150.770 298.235 158.770 298.405 ;
        RECT 159.060 298.235 167.060 298.405 ;
        RECT 176.770 298.235 184.770 298.405 ;
        RECT 185.060 298.235 193.060 298.405 ;
        RECT 202.770 298.235 210.770 298.405 ;
        RECT 211.060 298.235 219.060 298.405 ;
        RECT 228.770 298.235 236.770 298.405 ;
        RECT 237.060 298.235 245.060 298.405 ;
        RECT 254.770 298.235 262.770 298.405 ;
        RECT 263.060 298.235 271.060 298.405 ;
        RECT 280.770 298.235 288.770 298.405 ;
        RECT 289.060 298.235 297.060 298.405 ;
        RECT 46.770 290.595 54.770 290.765 ;
        RECT 55.060 290.595 63.060 290.765 ;
        RECT 72.770 290.595 80.770 290.765 ;
        RECT 81.060 290.595 89.060 290.765 ;
        RECT 98.770 290.595 106.770 290.765 ;
        RECT 107.060 290.595 115.060 290.765 ;
        RECT 124.770 290.595 132.770 290.765 ;
        RECT 133.060 290.595 141.060 290.765 ;
        RECT 150.770 290.595 158.770 290.765 ;
        RECT 159.060 290.595 167.060 290.765 ;
        RECT 176.770 290.595 184.770 290.765 ;
        RECT 185.060 290.595 193.060 290.765 ;
        RECT 202.770 290.595 210.770 290.765 ;
        RECT 211.060 290.595 219.060 290.765 ;
        RECT 228.770 290.595 236.770 290.765 ;
        RECT 237.060 290.595 245.060 290.765 ;
        RECT 254.770 290.595 262.770 290.765 ;
        RECT 263.060 290.595 271.060 290.765 ;
        RECT 280.770 290.595 288.770 290.765 ;
        RECT 289.060 290.595 297.060 290.765 ;
        RECT 46.770 290.055 54.770 290.225 ;
        RECT 55.060 290.055 63.060 290.225 ;
        RECT 72.770 290.055 80.770 290.225 ;
        RECT 81.060 290.055 89.060 290.225 ;
        RECT 98.770 290.055 106.770 290.225 ;
        RECT 107.060 290.055 115.060 290.225 ;
        RECT 124.770 290.055 132.770 290.225 ;
        RECT 133.060 290.055 141.060 290.225 ;
        RECT 150.770 290.055 158.770 290.225 ;
        RECT 159.060 290.055 167.060 290.225 ;
        RECT 176.770 290.055 184.770 290.225 ;
        RECT 185.060 290.055 193.060 290.225 ;
        RECT 202.770 290.055 210.770 290.225 ;
        RECT 211.060 290.055 219.060 290.225 ;
        RECT 228.770 290.055 236.770 290.225 ;
        RECT 237.060 290.055 245.060 290.225 ;
        RECT 254.770 290.055 262.770 290.225 ;
        RECT 263.060 290.055 271.060 290.225 ;
        RECT 280.770 290.055 288.770 290.225 ;
        RECT 289.060 290.055 297.060 290.225 ;
        RECT 46.770 282.415 54.770 282.585 ;
        RECT 55.060 282.415 63.060 282.585 ;
        RECT 72.770 282.415 80.770 282.585 ;
        RECT 81.060 282.415 89.060 282.585 ;
        RECT 98.770 282.415 106.770 282.585 ;
        RECT 107.060 282.415 115.060 282.585 ;
        RECT 124.770 282.415 132.770 282.585 ;
        RECT 133.060 282.415 141.060 282.585 ;
        RECT 150.770 282.415 158.770 282.585 ;
        RECT 159.060 282.415 167.060 282.585 ;
        RECT 176.770 282.415 184.770 282.585 ;
        RECT 185.060 282.415 193.060 282.585 ;
        RECT 202.770 282.415 210.770 282.585 ;
        RECT 211.060 282.415 219.060 282.585 ;
        RECT 228.770 282.415 236.770 282.585 ;
        RECT 237.060 282.415 245.060 282.585 ;
        RECT 254.770 282.415 262.770 282.585 ;
        RECT 263.060 282.415 271.060 282.585 ;
        RECT 280.770 282.415 288.770 282.585 ;
        RECT 289.060 282.415 297.060 282.585 ;
        RECT 46.770 281.875 54.770 282.045 ;
        RECT 55.060 281.875 63.060 282.045 ;
        RECT 72.770 281.875 80.770 282.045 ;
        RECT 81.060 281.875 89.060 282.045 ;
        RECT 98.770 281.875 106.770 282.045 ;
        RECT 107.060 281.875 115.060 282.045 ;
        RECT 124.770 281.875 132.770 282.045 ;
        RECT 133.060 281.875 141.060 282.045 ;
        RECT 150.770 281.875 158.770 282.045 ;
        RECT 159.060 281.875 167.060 282.045 ;
        RECT 176.770 281.875 184.770 282.045 ;
        RECT 185.060 281.875 193.060 282.045 ;
        RECT 202.770 281.875 210.770 282.045 ;
        RECT 211.060 281.875 219.060 282.045 ;
        RECT 228.770 281.875 236.770 282.045 ;
        RECT 237.060 281.875 245.060 282.045 ;
        RECT 254.770 281.875 262.770 282.045 ;
        RECT 263.060 281.875 271.060 282.045 ;
        RECT 280.770 281.875 288.770 282.045 ;
        RECT 289.060 281.875 297.060 282.045 ;
        RECT 46.770 274.235 54.770 274.405 ;
        RECT 55.060 274.235 63.060 274.405 ;
        RECT 72.770 274.235 80.770 274.405 ;
        RECT 81.060 274.235 89.060 274.405 ;
        RECT 98.770 274.235 106.770 274.405 ;
        RECT 107.060 274.235 115.060 274.405 ;
        RECT 124.770 274.235 132.770 274.405 ;
        RECT 133.060 274.235 141.060 274.405 ;
        RECT 150.770 274.235 158.770 274.405 ;
        RECT 159.060 274.235 167.060 274.405 ;
        RECT 176.770 274.235 184.770 274.405 ;
        RECT 185.060 274.235 193.060 274.405 ;
        RECT 202.770 274.235 210.770 274.405 ;
        RECT 211.060 274.235 219.060 274.405 ;
        RECT 228.770 274.235 236.770 274.405 ;
        RECT 237.060 274.235 245.060 274.405 ;
        RECT 254.770 274.235 262.770 274.405 ;
        RECT 263.060 274.235 271.060 274.405 ;
        RECT 280.770 274.235 288.770 274.405 ;
        RECT 289.060 274.235 297.060 274.405 ;
        RECT 46.770 273.695 54.770 273.865 ;
        RECT 55.060 273.695 63.060 273.865 ;
        RECT 72.770 273.695 80.770 273.865 ;
        RECT 81.060 273.695 89.060 273.865 ;
        RECT 98.770 273.695 106.770 273.865 ;
        RECT 107.060 273.695 115.060 273.865 ;
        RECT 124.770 273.695 132.770 273.865 ;
        RECT 133.060 273.695 141.060 273.865 ;
        RECT 150.770 273.695 158.770 273.865 ;
        RECT 159.060 273.695 167.060 273.865 ;
        RECT 176.770 273.695 184.770 273.865 ;
        RECT 185.060 273.695 193.060 273.865 ;
        RECT 202.770 273.695 210.770 273.865 ;
        RECT 211.060 273.695 219.060 273.865 ;
        RECT 228.770 273.695 236.770 273.865 ;
        RECT 237.060 273.695 245.060 273.865 ;
        RECT 254.770 273.695 262.770 273.865 ;
        RECT 263.060 273.695 271.060 273.865 ;
        RECT 280.770 273.695 288.770 273.865 ;
        RECT 289.060 273.695 297.060 273.865 ;
        RECT 46.770 266.055 54.770 266.225 ;
        RECT 55.060 266.055 63.060 266.225 ;
        RECT 72.770 266.055 80.770 266.225 ;
        RECT 81.060 266.055 89.060 266.225 ;
        RECT 98.770 266.055 106.770 266.225 ;
        RECT 107.060 266.055 115.060 266.225 ;
        RECT 124.770 266.055 132.770 266.225 ;
        RECT 133.060 266.055 141.060 266.225 ;
        RECT 150.770 266.055 158.770 266.225 ;
        RECT 159.060 266.055 167.060 266.225 ;
        RECT 176.770 266.055 184.770 266.225 ;
        RECT 185.060 266.055 193.060 266.225 ;
        RECT 202.770 266.055 210.770 266.225 ;
        RECT 211.060 266.055 219.060 266.225 ;
        RECT 228.770 266.055 236.770 266.225 ;
        RECT 237.060 266.055 245.060 266.225 ;
        RECT 254.770 266.055 262.770 266.225 ;
        RECT 263.060 266.055 271.060 266.225 ;
        RECT 280.770 266.055 288.770 266.225 ;
        RECT 289.060 266.055 297.060 266.225 ;
        RECT 46.770 265.515 54.770 265.685 ;
        RECT 55.060 265.515 63.060 265.685 ;
        RECT 72.770 265.515 80.770 265.685 ;
        RECT 81.060 265.515 89.060 265.685 ;
        RECT 98.770 265.515 106.770 265.685 ;
        RECT 107.060 265.515 115.060 265.685 ;
        RECT 124.770 265.515 132.770 265.685 ;
        RECT 133.060 265.515 141.060 265.685 ;
        RECT 150.770 265.515 158.770 265.685 ;
        RECT 159.060 265.515 167.060 265.685 ;
        RECT 176.770 265.515 184.770 265.685 ;
        RECT 185.060 265.515 193.060 265.685 ;
        RECT 202.770 265.515 210.770 265.685 ;
        RECT 211.060 265.515 219.060 265.685 ;
        RECT 228.770 265.515 236.770 265.685 ;
        RECT 237.060 265.515 245.060 265.685 ;
        RECT 254.770 265.515 262.770 265.685 ;
        RECT 263.060 265.515 271.060 265.685 ;
        RECT 280.770 265.515 288.770 265.685 ;
        RECT 289.060 265.515 297.060 265.685 ;
        RECT 46.770 257.875 54.770 258.045 ;
        RECT 55.060 257.875 63.060 258.045 ;
        RECT 72.770 257.875 80.770 258.045 ;
        RECT 81.060 257.875 89.060 258.045 ;
        RECT 98.770 257.875 106.770 258.045 ;
        RECT 107.060 257.875 115.060 258.045 ;
        RECT 124.770 257.875 132.770 258.045 ;
        RECT 133.060 257.875 141.060 258.045 ;
        RECT 150.770 257.875 158.770 258.045 ;
        RECT 159.060 257.875 167.060 258.045 ;
        RECT 176.770 257.875 184.770 258.045 ;
        RECT 185.060 257.875 193.060 258.045 ;
        RECT 202.770 257.875 210.770 258.045 ;
        RECT 211.060 257.875 219.060 258.045 ;
        RECT 228.770 257.875 236.770 258.045 ;
        RECT 237.060 257.875 245.060 258.045 ;
        RECT 254.770 257.875 262.770 258.045 ;
        RECT 263.060 257.875 271.060 258.045 ;
        RECT 280.770 257.875 288.770 258.045 ;
        RECT 289.060 257.875 297.060 258.045 ;
        RECT 46.770 257.335 54.770 257.505 ;
        RECT 55.060 257.335 63.060 257.505 ;
        RECT 72.770 257.335 80.770 257.505 ;
        RECT 81.060 257.335 89.060 257.505 ;
        RECT 98.770 257.335 106.770 257.505 ;
        RECT 107.060 257.335 115.060 257.505 ;
        RECT 124.770 257.335 132.770 257.505 ;
        RECT 133.060 257.335 141.060 257.505 ;
        RECT 150.770 257.335 158.770 257.505 ;
        RECT 159.060 257.335 167.060 257.505 ;
        RECT 176.770 257.335 184.770 257.505 ;
        RECT 185.060 257.335 193.060 257.505 ;
        RECT 202.770 257.335 210.770 257.505 ;
        RECT 211.060 257.335 219.060 257.505 ;
        RECT 228.770 257.335 236.770 257.505 ;
        RECT 237.060 257.335 245.060 257.505 ;
        RECT 254.770 257.335 262.770 257.505 ;
        RECT 263.060 257.335 271.060 257.505 ;
        RECT 280.770 257.335 288.770 257.505 ;
        RECT 289.060 257.335 297.060 257.505 ;
        RECT 46.770 249.695 54.770 249.865 ;
        RECT 55.060 249.695 63.060 249.865 ;
        RECT 72.770 249.695 80.770 249.865 ;
        RECT 81.060 249.695 89.060 249.865 ;
        RECT 98.770 249.695 106.770 249.865 ;
        RECT 107.060 249.695 115.060 249.865 ;
        RECT 124.770 249.695 132.770 249.865 ;
        RECT 133.060 249.695 141.060 249.865 ;
        RECT 150.770 249.695 158.770 249.865 ;
        RECT 159.060 249.695 167.060 249.865 ;
        RECT 176.770 249.695 184.770 249.865 ;
        RECT 185.060 249.695 193.060 249.865 ;
        RECT 202.770 249.695 210.770 249.865 ;
        RECT 211.060 249.695 219.060 249.865 ;
        RECT 228.770 249.695 236.770 249.865 ;
        RECT 237.060 249.695 245.060 249.865 ;
        RECT 254.770 249.695 262.770 249.865 ;
        RECT 263.060 249.695 271.060 249.865 ;
        RECT 280.770 249.695 288.770 249.865 ;
        RECT 289.060 249.695 297.060 249.865 ;
        RECT 46.770 249.155 54.770 249.325 ;
        RECT 55.060 249.155 63.060 249.325 ;
        RECT 72.770 249.155 80.770 249.325 ;
        RECT 81.060 249.155 89.060 249.325 ;
        RECT 98.770 249.155 106.770 249.325 ;
        RECT 107.060 249.155 115.060 249.325 ;
        RECT 124.770 249.155 132.770 249.325 ;
        RECT 133.060 249.155 141.060 249.325 ;
        RECT 150.770 249.155 158.770 249.325 ;
        RECT 159.060 249.155 167.060 249.325 ;
        RECT 176.770 249.155 184.770 249.325 ;
        RECT 185.060 249.155 193.060 249.325 ;
        RECT 202.770 249.155 210.770 249.325 ;
        RECT 211.060 249.155 219.060 249.325 ;
        RECT 228.770 249.155 236.770 249.325 ;
        RECT 237.060 249.155 245.060 249.325 ;
        RECT 254.770 249.155 262.770 249.325 ;
        RECT 263.060 249.155 271.060 249.325 ;
        RECT 280.770 249.155 288.770 249.325 ;
        RECT 289.060 249.155 297.060 249.325 ;
        RECT 46.770 241.515 54.770 241.685 ;
        RECT 55.060 241.515 63.060 241.685 ;
        RECT 72.770 241.515 80.770 241.685 ;
        RECT 81.060 241.515 89.060 241.685 ;
        RECT 98.770 241.515 106.770 241.685 ;
        RECT 107.060 241.515 115.060 241.685 ;
        RECT 124.770 241.515 132.770 241.685 ;
        RECT 133.060 241.515 141.060 241.685 ;
        RECT 150.770 241.515 158.770 241.685 ;
        RECT 159.060 241.515 167.060 241.685 ;
        RECT 176.770 241.515 184.770 241.685 ;
        RECT 185.060 241.515 193.060 241.685 ;
        RECT 202.770 241.515 210.770 241.685 ;
        RECT 211.060 241.515 219.060 241.685 ;
        RECT 228.770 241.515 236.770 241.685 ;
        RECT 237.060 241.515 245.060 241.685 ;
        RECT 254.770 241.515 262.770 241.685 ;
        RECT 263.060 241.515 271.060 241.685 ;
        RECT 280.770 241.515 288.770 241.685 ;
        RECT 289.060 241.515 297.060 241.685 ;
        RECT 46.770 240.975 54.770 241.145 ;
        RECT 55.060 240.975 63.060 241.145 ;
        RECT 72.770 240.975 80.770 241.145 ;
        RECT 81.060 240.975 89.060 241.145 ;
        RECT 98.770 240.975 106.770 241.145 ;
        RECT 107.060 240.975 115.060 241.145 ;
        RECT 124.770 240.975 132.770 241.145 ;
        RECT 133.060 240.975 141.060 241.145 ;
        RECT 150.770 240.975 158.770 241.145 ;
        RECT 159.060 240.975 167.060 241.145 ;
        RECT 176.770 240.975 184.770 241.145 ;
        RECT 185.060 240.975 193.060 241.145 ;
        RECT 202.770 240.975 210.770 241.145 ;
        RECT 211.060 240.975 219.060 241.145 ;
        RECT 228.770 240.975 236.770 241.145 ;
        RECT 237.060 240.975 245.060 241.145 ;
        RECT 254.770 240.975 262.770 241.145 ;
        RECT 263.060 240.975 271.060 241.145 ;
        RECT 280.770 240.975 288.770 241.145 ;
        RECT 289.060 240.975 297.060 241.145 ;
        RECT 46.770 233.335 54.770 233.505 ;
        RECT 55.060 233.335 63.060 233.505 ;
        RECT 72.770 233.335 80.770 233.505 ;
        RECT 81.060 233.335 89.060 233.505 ;
        RECT 98.770 233.335 106.770 233.505 ;
        RECT 107.060 233.335 115.060 233.505 ;
        RECT 124.770 233.335 132.770 233.505 ;
        RECT 133.060 233.335 141.060 233.505 ;
        RECT 150.770 233.335 158.770 233.505 ;
        RECT 159.060 233.335 167.060 233.505 ;
        RECT 176.770 233.335 184.770 233.505 ;
        RECT 185.060 233.335 193.060 233.505 ;
        RECT 202.770 233.335 210.770 233.505 ;
        RECT 211.060 233.335 219.060 233.505 ;
        RECT 228.770 233.335 236.770 233.505 ;
        RECT 237.060 233.335 245.060 233.505 ;
        RECT 254.770 233.335 262.770 233.505 ;
        RECT 263.060 233.335 271.060 233.505 ;
        RECT 280.770 233.335 288.770 233.505 ;
        RECT 289.060 233.335 297.060 233.505 ;
        RECT 46.770 232.795 54.770 232.965 ;
        RECT 55.060 232.795 63.060 232.965 ;
        RECT 72.770 232.795 80.770 232.965 ;
        RECT 81.060 232.795 89.060 232.965 ;
        RECT 98.770 232.795 106.770 232.965 ;
        RECT 107.060 232.795 115.060 232.965 ;
        RECT 124.770 232.795 132.770 232.965 ;
        RECT 133.060 232.795 141.060 232.965 ;
        RECT 150.770 232.795 158.770 232.965 ;
        RECT 159.060 232.795 167.060 232.965 ;
        RECT 176.770 232.795 184.770 232.965 ;
        RECT 185.060 232.795 193.060 232.965 ;
        RECT 202.770 232.795 210.770 232.965 ;
        RECT 211.060 232.795 219.060 232.965 ;
        RECT 228.770 232.795 236.770 232.965 ;
        RECT 237.060 232.795 245.060 232.965 ;
        RECT 254.770 232.795 262.770 232.965 ;
        RECT 263.060 232.795 271.060 232.965 ;
        RECT 280.770 232.795 288.770 232.965 ;
        RECT 289.060 232.795 297.060 232.965 ;
        RECT 46.770 225.155 54.770 225.325 ;
        RECT 55.060 225.155 63.060 225.325 ;
        RECT 72.770 225.155 80.770 225.325 ;
        RECT 81.060 225.155 89.060 225.325 ;
        RECT 98.770 225.155 106.770 225.325 ;
        RECT 107.060 225.155 115.060 225.325 ;
        RECT 124.770 225.155 132.770 225.325 ;
        RECT 133.060 225.155 141.060 225.325 ;
        RECT 150.770 225.155 158.770 225.325 ;
        RECT 159.060 225.155 167.060 225.325 ;
        RECT 176.770 225.155 184.770 225.325 ;
        RECT 185.060 225.155 193.060 225.325 ;
        RECT 202.770 225.155 210.770 225.325 ;
        RECT 211.060 225.155 219.060 225.325 ;
        RECT 228.770 225.155 236.770 225.325 ;
        RECT 237.060 225.155 245.060 225.325 ;
        RECT 254.770 225.155 262.770 225.325 ;
        RECT 263.060 225.155 271.060 225.325 ;
        RECT 280.770 225.155 288.770 225.325 ;
        RECT 289.060 225.155 297.060 225.325 ;
        RECT 46.770 224.615 54.770 224.785 ;
        RECT 55.060 224.615 63.060 224.785 ;
        RECT 72.770 224.615 80.770 224.785 ;
        RECT 81.060 224.615 89.060 224.785 ;
        RECT 98.770 224.615 106.770 224.785 ;
        RECT 107.060 224.615 115.060 224.785 ;
        RECT 124.770 224.615 132.770 224.785 ;
        RECT 133.060 224.615 141.060 224.785 ;
        RECT 150.770 224.615 158.770 224.785 ;
        RECT 159.060 224.615 167.060 224.785 ;
        RECT 176.770 224.615 184.770 224.785 ;
        RECT 185.060 224.615 193.060 224.785 ;
        RECT 202.770 224.615 210.770 224.785 ;
        RECT 211.060 224.615 219.060 224.785 ;
        RECT 228.770 224.615 236.770 224.785 ;
        RECT 237.060 224.615 245.060 224.785 ;
        RECT 254.770 224.615 262.770 224.785 ;
        RECT 263.060 224.615 271.060 224.785 ;
        RECT 280.770 224.615 288.770 224.785 ;
        RECT 289.060 224.615 297.060 224.785 ;
        RECT 46.770 216.975 54.770 217.145 ;
        RECT 55.060 216.975 63.060 217.145 ;
        RECT 72.770 216.975 80.770 217.145 ;
        RECT 81.060 216.975 89.060 217.145 ;
        RECT 98.770 216.975 106.770 217.145 ;
        RECT 107.060 216.975 115.060 217.145 ;
        RECT 124.770 216.975 132.770 217.145 ;
        RECT 133.060 216.975 141.060 217.145 ;
        RECT 150.770 216.975 158.770 217.145 ;
        RECT 159.060 216.975 167.060 217.145 ;
        RECT 176.770 216.975 184.770 217.145 ;
        RECT 185.060 216.975 193.060 217.145 ;
        RECT 202.770 216.975 210.770 217.145 ;
        RECT 211.060 216.975 219.060 217.145 ;
        RECT 228.770 216.975 236.770 217.145 ;
        RECT 237.060 216.975 245.060 217.145 ;
        RECT 254.770 216.975 262.770 217.145 ;
        RECT 263.060 216.975 271.060 217.145 ;
        RECT 280.770 216.975 288.770 217.145 ;
        RECT 289.060 216.975 297.060 217.145 ;
        RECT 46.770 216.435 54.770 216.605 ;
        RECT 55.060 216.435 63.060 216.605 ;
        RECT 72.770 216.435 80.770 216.605 ;
        RECT 81.060 216.435 89.060 216.605 ;
        RECT 98.770 216.435 106.770 216.605 ;
        RECT 107.060 216.435 115.060 216.605 ;
        RECT 124.770 216.435 132.770 216.605 ;
        RECT 133.060 216.435 141.060 216.605 ;
        RECT 150.770 216.435 158.770 216.605 ;
        RECT 159.060 216.435 167.060 216.605 ;
        RECT 176.770 216.435 184.770 216.605 ;
        RECT 185.060 216.435 193.060 216.605 ;
        RECT 202.770 216.435 210.770 216.605 ;
        RECT 211.060 216.435 219.060 216.605 ;
        RECT 228.770 216.435 236.770 216.605 ;
        RECT 237.060 216.435 245.060 216.605 ;
        RECT 254.770 216.435 262.770 216.605 ;
        RECT 263.060 216.435 271.060 216.605 ;
        RECT 280.770 216.435 288.770 216.605 ;
        RECT 289.060 216.435 297.060 216.605 ;
        RECT 46.770 208.795 54.770 208.965 ;
        RECT 55.060 208.795 63.060 208.965 ;
        RECT 72.770 208.795 80.770 208.965 ;
        RECT 81.060 208.795 89.060 208.965 ;
        RECT 98.770 208.795 106.770 208.965 ;
        RECT 107.060 208.795 115.060 208.965 ;
        RECT 124.770 208.795 132.770 208.965 ;
        RECT 133.060 208.795 141.060 208.965 ;
        RECT 150.770 208.795 158.770 208.965 ;
        RECT 159.060 208.795 167.060 208.965 ;
        RECT 176.770 208.795 184.770 208.965 ;
        RECT 185.060 208.795 193.060 208.965 ;
        RECT 202.770 208.795 210.770 208.965 ;
        RECT 211.060 208.795 219.060 208.965 ;
        RECT 228.770 208.795 236.770 208.965 ;
        RECT 237.060 208.795 245.060 208.965 ;
        RECT 254.770 208.795 262.770 208.965 ;
        RECT 263.060 208.795 271.060 208.965 ;
        RECT 280.770 208.795 288.770 208.965 ;
        RECT 289.060 208.795 297.060 208.965 ;
        RECT 46.770 208.255 54.770 208.425 ;
        RECT 55.060 208.255 63.060 208.425 ;
        RECT 72.770 208.255 80.770 208.425 ;
        RECT 81.060 208.255 89.060 208.425 ;
        RECT 98.770 208.255 106.770 208.425 ;
        RECT 107.060 208.255 115.060 208.425 ;
        RECT 124.770 208.255 132.770 208.425 ;
        RECT 133.060 208.255 141.060 208.425 ;
        RECT 150.770 208.255 158.770 208.425 ;
        RECT 159.060 208.255 167.060 208.425 ;
        RECT 176.770 208.255 184.770 208.425 ;
        RECT 185.060 208.255 193.060 208.425 ;
        RECT 202.770 208.255 210.770 208.425 ;
        RECT 211.060 208.255 219.060 208.425 ;
        RECT 228.770 208.255 236.770 208.425 ;
        RECT 237.060 208.255 245.060 208.425 ;
        RECT 254.770 208.255 262.770 208.425 ;
        RECT 263.060 208.255 271.060 208.425 ;
        RECT 280.770 208.255 288.770 208.425 ;
        RECT 289.060 208.255 297.060 208.425 ;
        RECT 46.770 200.615 54.770 200.785 ;
        RECT 55.060 200.615 63.060 200.785 ;
        RECT 72.770 200.615 80.770 200.785 ;
        RECT 81.060 200.615 89.060 200.785 ;
        RECT 98.770 200.615 106.770 200.785 ;
        RECT 107.060 200.615 115.060 200.785 ;
        RECT 124.770 200.615 132.770 200.785 ;
        RECT 133.060 200.615 141.060 200.785 ;
        RECT 150.770 200.615 158.770 200.785 ;
        RECT 159.060 200.615 167.060 200.785 ;
        RECT 176.770 200.615 184.770 200.785 ;
        RECT 185.060 200.615 193.060 200.785 ;
        RECT 202.770 200.615 210.770 200.785 ;
        RECT 211.060 200.615 219.060 200.785 ;
        RECT 228.770 200.615 236.770 200.785 ;
        RECT 237.060 200.615 245.060 200.785 ;
        RECT 254.770 200.615 262.770 200.785 ;
        RECT 263.060 200.615 271.060 200.785 ;
        RECT 280.770 200.615 288.770 200.785 ;
        RECT 289.060 200.615 297.060 200.785 ;
        RECT 46.770 200.075 54.770 200.245 ;
        RECT 55.060 200.075 63.060 200.245 ;
        RECT 72.770 200.075 80.770 200.245 ;
        RECT 81.060 200.075 89.060 200.245 ;
        RECT 98.770 200.075 106.770 200.245 ;
        RECT 107.060 200.075 115.060 200.245 ;
        RECT 124.770 200.075 132.770 200.245 ;
        RECT 133.060 200.075 141.060 200.245 ;
        RECT 150.770 200.075 158.770 200.245 ;
        RECT 159.060 200.075 167.060 200.245 ;
        RECT 176.770 200.075 184.770 200.245 ;
        RECT 185.060 200.075 193.060 200.245 ;
        RECT 202.770 200.075 210.770 200.245 ;
        RECT 211.060 200.075 219.060 200.245 ;
        RECT 228.770 200.075 236.770 200.245 ;
        RECT 237.060 200.075 245.060 200.245 ;
        RECT 254.770 200.075 262.770 200.245 ;
        RECT 263.060 200.075 271.060 200.245 ;
        RECT 280.770 200.075 288.770 200.245 ;
        RECT 289.060 200.075 297.060 200.245 ;
        RECT 46.770 192.435 54.770 192.605 ;
        RECT 55.060 192.435 63.060 192.605 ;
        RECT 72.770 192.435 80.770 192.605 ;
        RECT 81.060 192.435 89.060 192.605 ;
        RECT 98.770 192.435 106.770 192.605 ;
        RECT 107.060 192.435 115.060 192.605 ;
        RECT 124.770 192.435 132.770 192.605 ;
        RECT 133.060 192.435 141.060 192.605 ;
        RECT 150.770 192.435 158.770 192.605 ;
        RECT 159.060 192.435 167.060 192.605 ;
        RECT 176.770 192.435 184.770 192.605 ;
        RECT 185.060 192.435 193.060 192.605 ;
        RECT 202.770 192.435 210.770 192.605 ;
        RECT 211.060 192.435 219.060 192.605 ;
        RECT 228.770 192.435 236.770 192.605 ;
        RECT 237.060 192.435 245.060 192.605 ;
        RECT 254.770 192.435 262.770 192.605 ;
        RECT 263.060 192.435 271.060 192.605 ;
        RECT 280.770 192.435 288.770 192.605 ;
        RECT 289.060 192.435 297.060 192.605 ;
        RECT 46.770 191.895 54.770 192.065 ;
        RECT 55.060 191.895 63.060 192.065 ;
        RECT 72.770 191.895 80.770 192.065 ;
        RECT 81.060 191.895 89.060 192.065 ;
        RECT 98.770 191.895 106.770 192.065 ;
        RECT 107.060 191.895 115.060 192.065 ;
        RECT 124.770 191.895 132.770 192.065 ;
        RECT 133.060 191.895 141.060 192.065 ;
        RECT 150.770 191.895 158.770 192.065 ;
        RECT 159.060 191.895 167.060 192.065 ;
        RECT 176.770 191.895 184.770 192.065 ;
        RECT 185.060 191.895 193.060 192.065 ;
        RECT 202.770 191.895 210.770 192.065 ;
        RECT 211.060 191.895 219.060 192.065 ;
        RECT 228.770 191.895 236.770 192.065 ;
        RECT 237.060 191.895 245.060 192.065 ;
        RECT 254.770 191.895 262.770 192.065 ;
        RECT 263.060 191.895 271.060 192.065 ;
        RECT 280.770 191.895 288.770 192.065 ;
        RECT 289.060 191.895 297.060 192.065 ;
        RECT 46.770 184.255 54.770 184.425 ;
        RECT 55.060 184.255 63.060 184.425 ;
        RECT 72.770 184.255 80.770 184.425 ;
        RECT 81.060 184.255 89.060 184.425 ;
        RECT 98.770 184.255 106.770 184.425 ;
        RECT 107.060 184.255 115.060 184.425 ;
        RECT 124.770 184.255 132.770 184.425 ;
        RECT 133.060 184.255 141.060 184.425 ;
        RECT 150.770 184.255 158.770 184.425 ;
        RECT 159.060 184.255 167.060 184.425 ;
        RECT 176.770 184.255 184.770 184.425 ;
        RECT 185.060 184.255 193.060 184.425 ;
        RECT 202.770 184.255 210.770 184.425 ;
        RECT 211.060 184.255 219.060 184.425 ;
        RECT 228.770 184.255 236.770 184.425 ;
        RECT 237.060 184.255 245.060 184.425 ;
        RECT 254.770 184.255 262.770 184.425 ;
        RECT 263.060 184.255 271.060 184.425 ;
        RECT 280.770 184.255 288.770 184.425 ;
        RECT 289.060 184.255 297.060 184.425 ;
        RECT 46.770 183.715 54.770 183.885 ;
        RECT 55.060 183.715 63.060 183.885 ;
        RECT 72.770 183.715 80.770 183.885 ;
        RECT 81.060 183.715 89.060 183.885 ;
        RECT 98.770 183.715 106.770 183.885 ;
        RECT 107.060 183.715 115.060 183.885 ;
        RECT 124.770 183.715 132.770 183.885 ;
        RECT 133.060 183.715 141.060 183.885 ;
        RECT 150.770 183.715 158.770 183.885 ;
        RECT 159.060 183.715 167.060 183.885 ;
        RECT 176.770 183.715 184.770 183.885 ;
        RECT 185.060 183.715 193.060 183.885 ;
        RECT 202.770 183.715 210.770 183.885 ;
        RECT 211.060 183.715 219.060 183.885 ;
        RECT 228.770 183.715 236.770 183.885 ;
        RECT 237.060 183.715 245.060 183.885 ;
        RECT 254.770 183.715 262.770 183.885 ;
        RECT 263.060 183.715 271.060 183.885 ;
        RECT 280.770 183.715 288.770 183.885 ;
        RECT 289.060 183.715 297.060 183.885 ;
        RECT 46.770 176.075 54.770 176.245 ;
        RECT 55.060 176.075 63.060 176.245 ;
        RECT 72.770 176.075 80.770 176.245 ;
        RECT 81.060 176.075 89.060 176.245 ;
        RECT 98.770 176.075 106.770 176.245 ;
        RECT 107.060 176.075 115.060 176.245 ;
        RECT 124.770 176.075 132.770 176.245 ;
        RECT 133.060 176.075 141.060 176.245 ;
        RECT 150.770 176.075 158.770 176.245 ;
        RECT 159.060 176.075 167.060 176.245 ;
        RECT 176.770 176.075 184.770 176.245 ;
        RECT 185.060 176.075 193.060 176.245 ;
        RECT 202.770 176.075 210.770 176.245 ;
        RECT 211.060 176.075 219.060 176.245 ;
        RECT 228.770 176.075 236.770 176.245 ;
        RECT 237.060 176.075 245.060 176.245 ;
        RECT 254.770 176.075 262.770 176.245 ;
        RECT 263.060 176.075 271.060 176.245 ;
        RECT 280.770 176.075 288.770 176.245 ;
        RECT 289.060 176.075 297.060 176.245 ;
        RECT 46.770 175.535 54.770 175.705 ;
        RECT 55.060 175.535 63.060 175.705 ;
        RECT 72.770 175.535 80.770 175.705 ;
        RECT 81.060 175.535 89.060 175.705 ;
        RECT 98.770 175.535 106.770 175.705 ;
        RECT 107.060 175.535 115.060 175.705 ;
        RECT 124.770 175.535 132.770 175.705 ;
        RECT 133.060 175.535 141.060 175.705 ;
        RECT 150.770 175.535 158.770 175.705 ;
        RECT 159.060 175.535 167.060 175.705 ;
        RECT 176.770 175.535 184.770 175.705 ;
        RECT 185.060 175.535 193.060 175.705 ;
        RECT 202.770 175.535 210.770 175.705 ;
        RECT 211.060 175.535 219.060 175.705 ;
        RECT 228.770 175.535 236.770 175.705 ;
        RECT 237.060 175.535 245.060 175.705 ;
        RECT 254.770 175.535 262.770 175.705 ;
        RECT 263.060 175.535 271.060 175.705 ;
        RECT 280.770 175.535 288.770 175.705 ;
        RECT 289.060 175.535 297.060 175.705 ;
        RECT 46.770 167.895 54.770 168.065 ;
        RECT 55.060 167.895 63.060 168.065 ;
        RECT 72.770 167.895 80.770 168.065 ;
        RECT 81.060 167.895 89.060 168.065 ;
        RECT 98.770 167.895 106.770 168.065 ;
        RECT 107.060 167.895 115.060 168.065 ;
        RECT 124.770 167.895 132.770 168.065 ;
        RECT 133.060 167.895 141.060 168.065 ;
        RECT 150.770 167.895 158.770 168.065 ;
        RECT 159.060 167.895 167.060 168.065 ;
        RECT 176.770 167.895 184.770 168.065 ;
        RECT 185.060 167.895 193.060 168.065 ;
        RECT 202.770 167.895 210.770 168.065 ;
        RECT 211.060 167.895 219.060 168.065 ;
        RECT 228.770 167.895 236.770 168.065 ;
        RECT 237.060 167.895 245.060 168.065 ;
        RECT 254.770 167.895 262.770 168.065 ;
        RECT 263.060 167.895 271.060 168.065 ;
        RECT 280.770 167.895 288.770 168.065 ;
        RECT 289.060 167.895 297.060 168.065 ;
        RECT 168.270 160.670 169.000 160.900 ;
        RECT 174.360 160.720 174.890 160.870 ;
        RECT 168.280 160.470 168.750 160.670 ;
        RECT 169.760 160.665 174.890 160.720 ;
        RECT 169.740 160.495 174.890 160.665 ;
        RECT 169.760 160.470 174.890 160.495 ;
        RECT 168.280 160.130 168.710 160.470 ;
        RECT 171.540 160.460 174.890 160.470 ;
        RECT 169.100 158.320 169.270 160.200 ;
        RECT 169.580 158.320 169.750 160.200 ;
        RECT 170.060 158.320 170.230 160.200 ;
        RECT 170.540 158.320 170.710 160.200 ;
        RECT 171.020 158.320 171.190 160.200 ;
        RECT 171.540 158.220 171.780 160.460 ;
        RECT 174.360 160.360 174.890 160.460 ;
        RECT 171.540 158.200 171.790 158.220 ;
        RECT 168.460 158.025 170.540 158.070 ;
        RECT 168.460 157.855 170.550 158.025 ;
        RECT 168.460 157.760 170.540 157.855 ;
        RECT 168.460 155.890 168.650 157.760 ;
        RECT 171.550 157.470 171.790 158.200 ;
        RECT 171.150 157.460 171.790 157.470 ;
        RECT 169.480 157.200 171.790 157.460 ;
        RECT 169.480 157.190 171.180 157.200 ;
        RECT 171.550 157.190 171.790 157.200 ;
        RECT 168.860 156.100 169.030 156.980 ;
        RECT 169.340 156.100 169.510 156.980 ;
        RECT 169.820 156.100 169.990 156.980 ;
        RECT 170.300 156.100 170.470 156.980 ;
        RECT 170.780 156.100 170.950 156.980 ;
        RECT 168.460 155.850 170.320 155.890 ;
        RECT 173.020 155.850 173.540 156.010 ;
        RECT 168.460 155.640 173.540 155.850 ;
        RECT 168.460 155.630 170.320 155.640 ;
        RECT 173.020 155.500 173.540 155.640 ;
        RECT 386.380 148.990 386.750 151.150 ;
        RECT 387.990 149.000 388.350 151.160 ;
        RECT 387.990 148.990 388.340 149.000 ;
        RECT 129.260 137.285 129.590 137.455 ;
        RECT 151.160 136.845 151.490 137.015 ;
        RECT 120.790 136.395 124.870 136.565 ;
        RECT 126.790 135.610 127.100 136.090 ;
        RECT 129.560 135.740 129.730 136.680 ;
        RECT 171.950 136.615 172.280 136.785 ;
        RECT 142.690 135.955 146.770 136.125 ;
        RECT 148.730 135.190 149.040 135.670 ;
        RECT 151.460 135.300 151.630 136.240 ;
        RECT 163.480 135.725 167.560 135.895 ;
        RECT 169.480 134.970 169.790 135.450 ;
        RECT 172.250 135.070 172.420 136.010 ;
        RECT 121.810 132.830 122.140 133.000 ;
        RECT 129.180 132.780 129.510 132.950 ;
        RECT 129.480 132.215 129.650 132.545 ;
        RECT 143.710 132.390 144.040 132.560 ;
        RECT 309.310 132.545 309.570 133.230 ;
        RECT 310.240 132.545 310.570 133.230 ;
        RECT 151.080 132.340 151.410 132.510 ;
        RECT 164.500 132.160 164.830 132.330 ;
        RECT 171.870 132.110 172.200 132.280 ;
        RECT 129.180 131.810 129.510 131.980 ;
        RECT 151.380 131.775 151.550 132.105 ;
        RECT 172.170 131.545 172.340 131.875 ;
        RECT 151.080 131.370 151.410 131.540 ;
        RECT 309.310 131.465 309.545 132.545 ;
        RECT 310.300 132.515 310.570 132.545 ;
        RECT 310.740 132.705 310.940 132.945 ;
        RECT 311.750 132.705 312.555 132.945 ;
        RECT 310.740 132.535 312.555 132.705 ;
        RECT 312.725 132.680 313.175 132.945 ;
        RECT 314.060 132.680 314.305 132.945 ;
        RECT 312.725 132.580 314.305 132.680 ;
        RECT 310.400 132.365 310.570 132.515 ;
        RECT 312.000 132.510 312.555 132.535 ;
        RECT 312.985 132.510 314.305 132.580 ;
        RECT 310.400 132.145 310.605 132.365 ;
        RECT 171.870 131.140 172.200 131.310 ;
        RECT 309.310 131.135 310.245 131.465 ;
        RECT 310.425 131.250 310.605 132.145 ;
        RECT 311.250 131.420 311.830 132.365 ;
        RECT 312.000 132.325 312.360 132.510 ;
        RECT 122.060 127.330 122.400 131.040 ;
        RECT 309.310 130.635 309.590 131.135 ;
        RECT 310.425 131.080 311.505 131.250 ;
        RECT 312.000 131.190 312.225 132.325 ;
        RECT 312.395 131.825 312.815 132.155 ;
        RECT 310.425 130.965 310.595 131.080 ;
        RECT 310.190 130.605 310.595 130.965 ;
        RECT 311.265 131.010 311.505 131.080 ;
        RECT 312.395 131.010 312.565 131.825 ;
        RECT 312.985 131.510 313.155 132.510 ;
        RECT 315.140 132.280 315.355 133.120 ;
        RECT 313.325 131.820 313.495 132.240 ;
        RECT 314.280 132.110 315.355 132.280 ;
        RECT 315.710 132.250 316.030 133.125 ;
        RECT 314.280 131.820 314.450 132.110 ;
        RECT 313.325 131.650 314.450 131.820 ;
        RECT 312.735 131.470 313.155 131.510 ;
        RECT 314.620 131.470 314.810 131.930 ;
        RECT 315.140 131.530 315.310 132.110 ;
        RECT 312.735 131.270 314.810 131.470 ;
        RECT 314.980 131.270 315.310 131.530 ;
        RECT 312.735 131.180 313.425 131.270 ;
        RECT 315.480 131.100 315.660 131.930 ;
        RECT 313.750 131.010 315.660 131.100 ;
        RECT 311.265 130.930 315.660 131.010 ;
        RECT 315.830 131.640 316.030 132.250 ;
        RECT 316.410 131.990 316.740 132.480 ;
        RECT 317.410 131.990 317.680 133.065 ;
        RECT 316.410 131.980 317.680 131.990 ;
        RECT 316.410 131.810 318.215 131.980 ;
        RECT 315.830 131.450 317.755 131.640 ;
        RECT 311.265 130.840 313.965 130.930 ;
        RECT 315.830 130.840 316.030 131.450 ;
        RECT 317.935 131.280 318.215 131.810 ;
        RECT 317.435 131.030 318.215 131.280 ;
        RECT 318.385 131.030 318.645 133.130 ;
        RECT 143.960 126.890 144.300 130.600 ;
        RECT 318.455 130.465 318.645 131.030 ;
        RECT 319.315 131.835 319.620 132.695 ;
        RECT 319.315 131.505 320.205 131.835 ;
        RECT 319.315 130.595 319.680 131.505 ;
        RECT 320.375 130.545 320.600 133.285 ;
        RECT 323.000 132.580 323.260 133.265 ;
        RECT 323.930 132.580 324.260 133.265 ;
        RECT 323.000 131.500 323.235 132.580 ;
        RECT 323.990 132.550 324.260 132.580 ;
        RECT 324.430 132.740 324.630 132.980 ;
        RECT 325.440 132.740 326.245 132.980 ;
        RECT 324.430 132.570 326.245 132.740 ;
        RECT 326.415 132.715 326.865 132.980 ;
        RECT 327.750 132.715 327.995 132.980 ;
        RECT 326.415 132.615 327.995 132.715 ;
        RECT 323.405 131.740 323.785 132.410 ;
        RECT 324.090 132.400 324.260 132.550 ;
        RECT 325.690 132.545 326.245 132.570 ;
        RECT 326.675 132.545 327.995 132.615 ;
        RECT 324.090 132.180 324.295 132.400 ;
        RECT 323.000 131.170 323.935 131.500 ;
        RECT 324.115 131.285 324.295 132.180 ;
        RECT 324.940 131.455 325.520 132.400 ;
        RECT 325.690 132.360 326.050 132.545 ;
        RECT 323.000 130.670 323.280 131.170 ;
        RECT 324.115 131.115 325.195 131.285 ;
        RECT 325.690 131.225 325.915 132.360 ;
        RECT 326.085 131.860 326.505 132.190 ;
        RECT 324.115 131.000 324.285 131.115 ;
        RECT 323.880 130.640 324.285 131.000 ;
        RECT 324.955 131.045 325.195 131.115 ;
        RECT 326.085 131.045 326.255 131.860 ;
        RECT 326.675 131.545 326.845 132.545 ;
        RECT 328.830 132.315 329.045 133.155 ;
        RECT 327.015 131.855 327.185 132.275 ;
        RECT 327.970 132.145 329.045 132.315 ;
        RECT 329.400 132.285 329.720 133.160 ;
        RECT 327.970 131.855 328.140 132.145 ;
        RECT 327.015 131.685 328.140 131.855 ;
        RECT 326.425 131.505 326.845 131.545 ;
        RECT 328.310 131.505 328.500 131.965 ;
        RECT 328.830 131.565 329.000 132.145 ;
        RECT 326.425 131.305 328.500 131.505 ;
        RECT 328.670 131.305 329.000 131.565 ;
        RECT 326.425 131.215 327.115 131.305 ;
        RECT 329.170 131.135 329.350 131.965 ;
        RECT 327.440 131.045 329.350 131.135 ;
        RECT 324.955 130.965 329.350 131.045 ;
        RECT 329.520 131.675 329.720 132.285 ;
        RECT 330.100 132.025 330.430 132.515 ;
        RECT 331.100 132.025 331.370 133.100 ;
        RECT 330.100 132.015 331.370 132.025 ;
        RECT 330.100 131.845 331.905 132.015 ;
        RECT 329.520 131.485 331.445 131.675 ;
        RECT 324.955 130.875 327.655 130.965 ;
        RECT 329.520 130.875 329.720 131.485 ;
        RECT 331.625 131.315 331.905 131.845 ;
        RECT 331.125 131.065 331.905 131.315 ;
        RECT 332.075 131.065 332.335 133.165 ;
        RECT 332.145 130.500 332.335 131.065 ;
        RECT 333.005 131.870 333.310 132.730 ;
        RECT 333.005 131.540 333.895 131.870 ;
        RECT 333.005 130.630 333.370 131.540 ;
        RECT 334.065 130.580 334.290 133.320 ;
        RECT 164.750 126.660 165.090 130.370 ;
        RECT 321.110 126.480 321.370 127.165 ;
        RECT 322.040 126.480 322.370 127.165 ;
        RECT 121.810 125.280 122.140 125.450 ;
        RECT 321.110 125.400 321.345 126.480 ;
        RECT 322.100 126.450 322.370 126.480 ;
        RECT 322.540 126.640 322.740 126.880 ;
        RECT 323.550 126.640 324.355 126.880 ;
        RECT 322.540 126.470 324.355 126.640 ;
        RECT 324.525 126.615 324.975 126.880 ;
        RECT 325.860 126.615 326.105 126.880 ;
        RECT 324.525 126.515 326.105 126.615 ;
        RECT 321.515 125.640 321.895 126.310 ;
        RECT 322.200 126.300 322.370 126.450 ;
        RECT 323.800 126.445 324.355 126.470 ;
        RECT 324.785 126.445 326.105 126.515 ;
        RECT 322.200 126.080 322.405 126.300 ;
        RECT 321.110 125.070 322.045 125.400 ;
        RECT 322.225 125.185 322.405 126.080 ;
        RECT 323.050 125.355 323.630 126.300 ;
        RECT 323.800 126.260 324.160 126.445 ;
        RECT 143.710 124.840 144.040 125.010 ;
        RECT 164.500 124.610 164.830 124.780 ;
        RECT 321.110 124.570 321.390 125.070 ;
        RECT 322.225 125.015 323.305 125.185 ;
        RECT 323.800 125.125 324.025 126.260 ;
        RECT 324.195 125.760 324.615 126.090 ;
        RECT 322.225 124.900 322.395 125.015 ;
        RECT 321.990 124.540 322.395 124.900 ;
        RECT 323.065 124.945 323.305 125.015 ;
        RECT 324.195 124.945 324.365 125.760 ;
        RECT 324.785 125.445 324.955 126.445 ;
        RECT 326.940 126.215 327.155 127.055 ;
        RECT 325.125 125.755 325.295 126.175 ;
        RECT 326.080 126.045 327.155 126.215 ;
        RECT 327.510 126.185 327.830 127.060 ;
        RECT 326.080 125.755 326.250 126.045 ;
        RECT 325.125 125.585 326.250 125.755 ;
        RECT 324.535 125.405 324.955 125.445 ;
        RECT 326.420 125.405 326.610 125.865 ;
        RECT 326.940 125.465 327.110 126.045 ;
        RECT 324.535 125.205 326.610 125.405 ;
        RECT 326.780 125.205 327.110 125.465 ;
        RECT 324.535 125.115 325.225 125.205 ;
        RECT 327.280 125.035 327.460 125.865 ;
        RECT 325.550 124.945 327.460 125.035 ;
        RECT 323.065 124.865 327.460 124.945 ;
        RECT 327.630 125.575 327.830 126.185 ;
        RECT 328.210 125.925 328.540 126.415 ;
        RECT 329.210 125.925 329.480 127.000 ;
        RECT 328.210 125.915 329.480 125.925 ;
        RECT 328.210 125.745 330.015 125.915 ;
        RECT 327.630 125.385 329.555 125.575 ;
        RECT 323.065 124.775 325.765 124.865 ;
        RECT 327.630 124.775 327.830 125.385 ;
        RECT 329.735 125.215 330.015 125.745 ;
        RECT 329.235 124.965 330.015 125.215 ;
        RECT 330.185 124.965 330.445 127.065 ;
        RECT 330.255 124.400 330.445 124.965 ;
        RECT 331.115 125.770 331.420 126.630 ;
        RECT 331.115 125.440 332.005 125.770 ;
        RECT 331.115 124.530 331.480 125.440 ;
        RECT 332.175 124.480 332.400 127.220 ;
        RECT 386.390 123.200 386.750 125.360 ;
        RECT 387.990 125.340 388.340 125.360 ;
        RECT 387.980 123.180 388.340 125.340 ;
        RECT 114.860 116.530 117.020 116.880 ;
        RECT 117.520 116.530 119.680 116.880 ;
        RECT 121.010 116.510 123.170 116.860 ;
        RECT 386.260 116.680 386.620 118.840 ;
        RECT 387.860 116.680 388.220 118.840 ;
        RECT 118.190 114.790 120.350 115.140 ;
        RECT 88.710 111.590 172.565 112.750 ;
        RECT 88.710 111.450 172.570 111.590 ;
        RECT 88.725 110.240 104.465 111.450 ;
        RECT 88.725 110.050 95.330 110.240 ;
        RECT 96.440 110.230 96.690 110.240 ;
        RECT 88.425 109.880 95.330 110.050 ;
        RECT 88.725 102.500 95.330 109.880 ;
        RECT 88.425 102.330 95.330 102.500 ;
        RECT 88.725 94.950 95.330 102.330 ;
        RECT 88.425 94.780 95.330 94.950 ;
        RECT 88.725 87.400 95.330 94.780 ;
        RECT 88.425 87.230 95.330 87.400 ;
        RECT 88.725 79.850 95.330 87.230 ;
        RECT 88.425 79.680 95.330 79.850 ;
        RECT 88.725 72.300 95.330 79.680 ;
        RECT 44.460 71.930 44.980 72.240 ;
        RECT 81.370 72.055 81.700 72.225 ;
        RECT 88.425 72.130 95.330 72.300 ;
        RECT 44.460 71.650 45.080 71.930 ;
        RECT 44.810 71.430 45.080 71.650 ;
        RECT 47.100 71.430 47.720 71.840 ;
        RECT 44.620 71.250 47.820 71.430 ;
        RECT 43.320 70.690 43.490 70.740 ;
        RECT 43.050 70.410 43.490 70.690 ;
        RECT 43.900 70.420 44.130 70.500 ;
        RECT 43.050 69.600 43.220 70.410 ;
        RECT 43.660 70.250 44.440 70.420 ;
        RECT 44.620 70.260 44.790 71.250 ;
        RECT 47.650 70.760 47.820 71.250 ;
        RECT 72.900 71.165 76.980 71.335 ;
        RECT 45.710 70.290 47.430 70.460 ;
        RECT 47.645 70.430 47.820 70.760 ;
        RECT 78.910 70.410 79.220 70.890 ;
        RECT 81.670 70.510 81.840 71.450 ;
        RECT 43.900 70.170 44.130 70.250 ;
        RECT 44.610 69.950 44.790 70.260 ;
        RECT 43.660 69.770 44.440 69.940 ;
        RECT 44.610 69.930 44.780 69.950 ;
        RECT 45.515 69.600 45.685 69.740 ;
        RECT 27.245 69.200 27.415 69.530 ;
        RECT 29.565 69.200 29.735 69.530 ;
        RECT 43.050 69.430 45.690 69.600 ;
        RECT 43.050 69.420 45.685 69.430 ;
        RECT 44.970 68.370 45.230 69.420 ;
        RECT 45.515 69.410 45.685 69.420 ;
        RECT 45.900 69.270 47.620 69.440 ;
        RECT 47.000 68.370 47.630 68.760 ;
        RECT 44.660 68.190 47.860 68.370 ;
        RECT 43.360 67.630 43.530 67.680 ;
        RECT 43.090 67.350 43.530 67.630 ;
        RECT 43.780 67.360 44.040 67.420 ;
        RECT 27.275 66.670 27.445 67.000 ;
        RECT 29.595 66.670 29.765 67.000 ;
        RECT 43.090 66.540 43.260 67.350 ;
        RECT 43.700 67.190 44.480 67.360 ;
        RECT 44.660 67.200 44.830 68.190 ;
        RECT 47.690 67.700 47.860 68.190 ;
        RECT 45.750 67.230 47.470 67.400 ;
        RECT 47.685 67.370 47.860 67.700 ;
        RECT 73.920 67.600 74.250 67.770 ;
        RECT 81.290 67.550 81.620 67.720 ;
        RECT 43.780 67.130 44.040 67.190 ;
        RECT 44.650 66.890 44.830 67.200 ;
        RECT 81.590 66.985 81.760 67.315 ;
        RECT 43.700 66.710 44.480 66.880 ;
        RECT 44.650 66.870 44.820 66.890 ;
        RECT 45.555 66.540 45.725 66.680 ;
        RECT 81.290 66.580 81.620 66.750 ;
        RECT 43.090 66.370 45.730 66.540 ;
        RECT 43.090 66.360 45.725 66.370 ;
        RECT 44.960 65.480 45.130 66.360 ;
        RECT 45.555 66.350 45.725 66.360 ;
        RECT 45.940 66.210 47.660 66.380 ;
        RECT 47.030 65.480 47.640 65.860 ;
        RECT 44.640 65.300 47.840 65.480 ;
        RECT 43.340 64.740 43.510 64.790 ;
        RECT 43.070 64.460 43.510 64.740 ;
        RECT 43.880 64.470 44.070 64.550 ;
        RECT 27.265 64.080 27.435 64.410 ;
        RECT 29.585 64.080 29.755 64.410 ;
        RECT 43.070 63.650 43.240 64.460 ;
        RECT 43.680 64.300 44.460 64.470 ;
        RECT 44.640 64.310 44.810 65.300 ;
        RECT 47.670 64.810 47.840 65.300 ;
        RECT 45.730 64.490 47.450 64.510 ;
        RECT 45.730 64.340 47.460 64.490 ;
        RECT 47.665 64.480 47.840 64.810 ;
        RECT 43.880 64.230 44.070 64.300 ;
        RECT 44.630 64.000 44.810 64.310 ;
        RECT 45.920 64.280 47.460 64.340 ;
        RECT 43.680 63.820 44.460 63.990 ;
        RECT 44.630 63.980 44.800 64.000 ;
        RECT 45.535 63.650 45.705 63.790 ;
        RECT 43.070 63.480 45.710 63.650 ;
        RECT 43.070 63.470 45.705 63.480 ;
        RECT 44.990 62.610 45.170 63.470 ;
        RECT 45.535 63.460 45.705 63.470 ;
        RECT 45.920 63.320 47.640 63.490 ;
        RECT 47.060 62.610 47.670 62.990 ;
        RECT 44.680 62.430 47.880 62.610 ;
        RECT 43.380 61.870 43.550 61.920 ;
        RECT 27.265 61.530 27.435 61.860 ;
        RECT 29.585 61.530 29.755 61.860 ;
        RECT 43.110 61.590 43.550 61.870 ;
        RECT 43.910 61.600 44.240 61.680 ;
        RECT 21.210 60.940 21.380 61.270 ;
        RECT 21.550 60.780 24.830 60.950 ;
        RECT 21.210 59.980 21.380 60.310 ;
        RECT 21.550 60.300 24.830 60.470 ;
        RECT 25.000 60.460 25.170 60.790 ;
        RECT 43.110 60.780 43.280 61.590 ;
        RECT 43.720 61.430 44.500 61.600 ;
        RECT 44.680 61.440 44.850 62.430 ;
        RECT 47.710 61.940 47.880 62.430 ;
        RECT 74.170 62.100 74.510 65.810 ;
        RECT 88.725 64.750 95.330 72.130 ;
        RECT 88.425 64.580 95.330 64.750 ;
        RECT 45.770 61.620 47.490 61.640 ;
        RECT 45.770 61.470 47.500 61.620 ;
        RECT 47.705 61.610 47.880 61.940 ;
        RECT 43.910 61.360 44.240 61.430 ;
        RECT 43.960 61.340 44.240 61.360 ;
        RECT 44.670 61.130 44.850 61.440 ;
        RECT 45.920 61.410 47.500 61.470 ;
        RECT 43.720 60.950 44.500 61.120 ;
        RECT 44.670 61.110 44.840 61.130 ;
        RECT 45.575 60.780 45.745 60.920 ;
        RECT 43.110 60.610 45.750 60.780 ;
        RECT 43.110 60.600 45.745 60.610 ;
        RECT 21.550 59.820 24.830 59.990 ;
        RECT 21.210 59.020 21.380 59.350 ;
        RECT 21.550 59.340 24.830 59.510 ;
        RECT 25.000 59.500 25.170 59.830 ;
        RECT 45.020 59.720 45.200 60.600 ;
        RECT 45.575 60.590 45.745 60.600 ;
        RECT 45.960 60.450 47.680 60.620 ;
        RECT 47.050 59.720 47.660 60.100 ;
        RECT 73.920 60.050 74.250 60.220 ;
        RECT 44.680 59.540 47.880 59.720 ;
        RECT 21.550 58.860 24.830 59.030 ;
        RECT 27.265 58.980 27.435 59.310 ;
        RECT 29.585 58.980 29.755 59.310 ;
        RECT 43.380 58.980 43.550 59.030 ;
        RECT 21.200 58.060 21.380 58.390 ;
        RECT 21.550 58.380 24.830 58.550 ;
        RECT 25.000 58.540 25.170 58.870 ;
        RECT 43.110 58.700 43.550 58.980 ;
        RECT 43.920 58.710 44.190 58.780 ;
        RECT 21.550 57.900 24.830 58.070 ;
        RECT 21.200 57.100 21.380 57.430 ;
        RECT 21.550 57.420 24.830 57.590 ;
        RECT 25.000 57.580 25.170 57.910 ;
        RECT 43.110 57.890 43.280 58.700 ;
        RECT 43.720 58.540 44.500 58.710 ;
        RECT 44.680 58.550 44.850 59.540 ;
        RECT 47.710 59.050 47.880 59.540 ;
        RECT 45.770 58.580 47.490 58.750 ;
        RECT 47.705 58.720 47.880 59.050 ;
        RECT 43.920 58.460 44.190 58.540 ;
        RECT 44.010 58.450 44.190 58.460 ;
        RECT 44.670 58.240 44.850 58.550 ;
        RECT 43.720 58.060 44.500 58.230 ;
        RECT 44.670 58.220 44.840 58.240 ;
        RECT 45.575 57.890 45.745 58.030 ;
        RECT 43.110 57.720 45.750 57.890 ;
        RECT 43.110 57.710 45.745 57.720 ;
        RECT 45.040 56.830 45.220 57.710 ;
        RECT 45.575 57.700 45.745 57.710 ;
        RECT 45.960 57.560 47.680 57.730 ;
        RECT 47.040 56.830 47.650 57.210 ;
        RECT 88.725 57.200 95.330 64.580 ;
        RECT 88.425 57.030 95.330 57.200 ;
        RECT 27.265 56.430 27.435 56.760 ;
        RECT 29.585 56.430 29.755 56.760 ;
        RECT 44.680 56.650 47.880 56.830 ;
        RECT 43.380 56.090 43.550 56.140 ;
        RECT 43.110 55.810 43.550 56.090 ;
        RECT 43.910 55.820 44.190 55.900 ;
        RECT 43.110 55.000 43.280 55.810 ;
        RECT 43.720 55.650 44.500 55.820 ;
        RECT 44.680 55.660 44.850 56.650 ;
        RECT 47.710 56.160 47.880 56.650 ;
        RECT 45.770 55.690 47.490 55.860 ;
        RECT 47.705 55.830 47.880 56.160 ;
        RECT 43.910 55.580 44.190 55.650 ;
        RECT 43.980 55.560 44.190 55.580 ;
        RECT 44.670 55.350 44.850 55.660 ;
        RECT 43.720 55.170 44.500 55.340 ;
        RECT 44.670 55.330 44.840 55.350 ;
        RECT 45.575 55.000 45.745 55.140 ;
        RECT 43.110 54.830 45.750 55.000 ;
        RECT 43.110 54.820 45.745 54.830 ;
        RECT 27.265 53.880 27.435 54.210 ;
        RECT 29.585 53.880 29.755 54.210 ;
        RECT 45.070 53.920 45.250 54.820 ;
        RECT 45.575 54.810 45.745 54.820 ;
        RECT 45.960 54.670 47.680 54.840 ;
        RECT 47.150 53.920 47.760 54.290 ;
        RECT 44.700 53.740 47.900 53.920 ;
        RECT 43.400 53.180 43.570 53.230 ;
        RECT 43.130 52.900 43.570 53.180 ;
        RECT 43.950 52.910 44.220 52.990 ;
        RECT 43.130 52.090 43.300 52.900 ;
        RECT 43.740 52.740 44.520 52.910 ;
        RECT 44.700 52.750 44.870 53.740 ;
        RECT 47.150 53.730 47.900 53.740 ;
        RECT 47.730 53.250 47.900 53.730 ;
        RECT 45.790 52.780 47.510 52.950 ;
        RECT 47.725 52.920 47.900 53.250 ;
        RECT 43.950 52.670 44.220 52.740 ;
        RECT 44.010 52.660 44.220 52.670 ;
        RECT 44.690 52.440 44.870 52.750 ;
        RECT 43.740 52.260 44.520 52.430 ;
        RECT 44.690 52.420 44.860 52.440 ;
        RECT 45.595 52.090 45.765 52.230 ;
        RECT 43.130 51.920 45.770 52.090 ;
        RECT 43.130 51.910 45.765 51.920 ;
        RECT 27.265 51.330 27.435 51.660 ;
        RECT 29.585 51.330 29.755 51.660 ;
        RECT 45.070 51.040 45.250 51.910 ;
        RECT 45.595 51.900 45.765 51.910 ;
        RECT 45.980 51.760 47.700 51.930 ;
        RECT 47.130 51.040 47.740 51.420 ;
        RECT 44.680 50.860 47.880 51.040 ;
        RECT 43.910 50.030 44.170 50.110 ;
        RECT 43.720 49.860 44.500 50.030 ;
        RECT 44.680 49.870 44.850 50.860 ;
        RECT 45.070 50.850 45.250 50.860 ;
        RECT 47.710 50.370 47.880 50.860 ;
        RECT 45.770 49.900 47.490 50.070 ;
        RECT 47.705 50.040 47.880 50.370 ;
        RECT 43.910 49.790 44.170 49.860 ;
        RECT 44.670 49.560 44.850 49.870 ;
        RECT 88.725 49.650 95.330 57.030 ;
        RECT 43.720 49.380 44.500 49.550 ;
        RECT 44.670 49.540 44.840 49.560 ;
        RECT 88.425 49.480 95.330 49.650 ;
        RECT 27.265 48.780 27.435 49.110 ;
        RECT 29.585 48.780 29.755 49.110 ;
        RECT 45.960 48.880 47.680 49.050 ;
        RECT 43.370 48.720 43.840 48.800 ;
        RECT 43.270 48.340 43.840 48.720 ;
        RECT 43.270 47.450 43.530 48.340 ;
        RECT 43.090 47.160 43.530 47.450 ;
        RECT 43.920 47.180 44.180 47.250 ;
        RECT 43.090 46.360 43.260 47.160 ;
        RECT 43.700 47.010 44.480 47.180 ;
        RECT 45.750 47.050 47.470 47.220 ;
        RECT 43.920 46.930 44.180 47.010 ;
        RECT 43.700 46.530 44.480 46.700 ;
        RECT 45.555 46.360 45.725 46.500 ;
        RECT 43.090 46.190 45.730 46.360 ;
        RECT 81.760 46.305 82.090 46.475 ;
        RECT 43.090 46.180 45.725 46.190 ;
        RECT 45.555 46.170 45.725 46.180 ;
        RECT 45.940 46.030 47.660 46.200 ;
        RECT 73.290 45.415 77.370 45.585 ;
        RECT 79.280 44.680 79.590 45.160 ;
        RECT 82.060 44.760 82.230 45.700 ;
        RECT 88.725 42.100 95.330 49.480 ;
        RECT 74.310 41.850 74.640 42.020 ;
        RECT 81.680 41.800 82.010 41.970 ;
        RECT 88.425 41.930 95.330 42.100 ;
        RECT 81.980 41.235 82.150 41.565 ;
        RECT 81.680 40.830 82.010 41.000 ;
        RECT 74.560 36.350 74.900 40.060 ;
        RECT 88.725 34.550 95.330 41.930 ;
        RECT 74.310 34.300 74.640 34.470 ;
        RECT 88.425 34.380 95.330 34.550 ;
        RECT 88.725 27.000 95.330 34.380 ;
        RECT 88.425 26.830 95.330 27.000 ;
        RECT 88.725 19.450 95.330 26.830 ;
        RECT 88.425 19.280 95.330 19.450 ;
        RECT 88.725 19.200 95.330 19.280 ;
        RECT 97.800 110.050 104.465 110.240 ;
        RECT 97.800 109.880 104.715 110.050 ;
        RECT 97.800 109.450 104.465 109.880 ;
        RECT 97.800 102.500 104.445 109.450 ;
        RECT 108.700 107.200 110.310 111.450 ;
        RECT 116.100 110.260 116.380 111.260 ;
        RECT 116.090 108.610 116.380 110.260 ;
        RECT 116.880 109.735 117.960 109.905 ;
        RECT 119.170 109.735 120.250 109.905 ;
        RECT 121.460 109.735 122.540 109.905 ;
        RECT 118.480 108.700 118.650 109.300 ;
        RECT 120.770 108.700 120.940 109.300 ;
        RECT 116.880 108.095 117.960 108.265 ;
        RECT 119.170 108.095 120.250 108.265 ;
        RECT 121.460 108.095 122.540 108.265 ;
        RECT 118.000 107.210 118.250 107.280 ;
        RECT 117.850 107.200 118.250 107.210 ;
        RECT 122.980 107.200 123.310 109.420 ;
        RECT 134.130 109.220 134.300 109.240 ;
        RECT 127.480 107.200 127.890 107.740 ;
        RECT 134.070 107.620 134.460 109.220 ;
        RECT 132.270 107.200 137.690 107.620 ;
        RECT 150.440 107.200 152.050 111.450 ;
        RECT 156.830 110.280 172.570 111.450 ;
        RECT 156.830 110.055 163.450 110.280 ;
        RECT 156.530 109.885 163.450 110.055 ;
        RECT 108.700 107.190 148.750 107.200 ;
        RECT 148.930 107.190 152.050 107.200 ;
        RECT 108.700 106.190 152.050 107.190 ;
        RECT 108.700 106.160 114.530 106.190 ;
        RECT 117.250 106.160 152.050 106.190 ;
        RECT 108.700 106.150 110.310 106.160 ;
        RECT 108.750 105.200 109.560 106.150 ;
        RECT 108.745 105.130 109.560 105.200 ;
        RECT 114.250 105.570 114.530 106.160 ;
        RECT 128.010 105.910 128.330 106.160 ;
        RECT 127.970 105.900 128.330 105.910 ;
        RECT 127.970 105.660 128.360 105.900 ;
        RECT 108.745 103.510 109.555 105.130 ;
        RECT 114.250 103.600 114.560 105.570 ;
        RECT 115.500 104.685 117.580 104.855 ;
        RECT 130.090 104.320 130.420 106.160 ;
        RECT 141.340 105.800 141.660 106.160 ;
        RECT 146.660 106.150 152.050 106.160 ;
        RECT 146.660 106.140 148.220 106.150 ;
        RECT 150.440 106.120 152.050 106.150 ;
        RECT 131.340 105.465 133.420 105.635 ;
        RECT 97.800 102.330 104.715 102.500 ;
        RECT 97.800 94.950 104.445 102.330 ;
        RECT 108.770 100.970 109.520 103.510 ;
        RECT 115.500 103.045 117.580 103.215 ;
        RECT 118.490 102.850 118.810 104.270 ;
        RECT 131.340 103.825 133.420 103.995 ;
        RECT 118.490 102.580 119.380 102.850 ;
        RECT 108.745 100.425 109.520 100.970 ;
        RECT 119.080 101.030 119.380 102.580 ;
        RECT 134.260 101.030 134.860 105.140 ;
        RECT 141.010 103.970 141.670 105.800 ;
        RECT 142.260 105.055 144.340 105.225 ;
        RECT 151.260 105.160 152.040 106.120 ;
        RECT 151.260 104.970 152.045 105.160 ;
        RECT 142.260 103.415 144.340 103.585 ;
        RECT 145.170 102.850 145.980 104.650 ;
        RECT 151.265 103.015 152.045 104.970 ;
        RECT 119.080 100.960 130.795 101.030 ;
        RECT 119.090 100.520 130.795 100.960 ;
        RECT 119.090 100.495 122.100 100.520 ;
        RECT 122.540 100.505 130.795 100.520 ;
        RECT 122.870 100.440 123.300 100.505 ;
        RECT 129.480 100.500 130.795 100.505 ;
        RECT 134.240 100.505 144.085 101.030 ;
        RECT 134.240 100.495 136.170 100.505 ;
        RECT 142.845 100.500 144.085 100.505 ;
        RECT 145.170 101.025 145.985 102.850 ;
        RECT 151.285 102.190 152.035 103.015 ;
        RECT 156.830 102.505 163.450 109.885 ;
        RECT 156.530 102.335 163.450 102.505 ;
        RECT 149.550 101.025 150.620 101.770 ;
        RECT 145.170 100.530 150.620 101.025 ;
        RECT 145.170 100.500 148.730 100.530 ;
        RECT 149.170 100.500 150.620 100.530 ;
        RECT 134.260 100.440 134.860 100.495 ;
        RECT 97.800 94.780 104.715 94.950 ;
        RECT 97.800 87.400 104.445 94.780 ;
        RECT 97.800 87.230 104.715 87.400 ;
        RECT 97.800 79.850 104.445 87.230 ;
        RECT 108.770 80.940 109.520 100.425 ;
        RECT 135.420 100.330 136.170 100.495 ;
        RECT 151.280 100.360 152.040 102.190 ;
        RECT 112.480 99.815 112.810 99.985 ;
        RECT 113.770 99.815 114.100 99.985 ;
        RECT 115.060 99.815 115.390 99.985 ;
        RECT 116.350 99.815 116.680 99.985 ;
        RECT 117.640 99.815 117.970 99.985 ;
        RECT 118.930 99.815 119.260 99.985 ;
        RECT 120.220 99.815 120.550 99.985 ;
        RECT 121.510 99.815 121.840 99.985 ;
        RECT 112.480 98.265 112.810 98.435 ;
        RECT 112.480 97.725 112.810 97.895 ;
        RECT 112.480 96.175 112.810 96.345 ;
        RECT 112.480 95.635 112.810 95.805 ;
        RECT 112.480 94.085 112.810 94.255 ;
        RECT 112.480 93.545 112.810 93.715 ;
        RECT 112.480 91.995 112.810 92.165 ;
        RECT 112.480 91.455 112.810 91.625 ;
        RECT 112.480 89.905 112.810 90.075 ;
        RECT 112.480 89.365 112.810 89.535 ;
        RECT 112.480 87.815 112.810 87.985 ;
        RECT 112.480 87.275 112.810 87.445 ;
        RECT 112.480 85.725 112.810 85.895 ;
        RECT 113.175 85.555 113.400 99.785 ;
        RECT 113.770 98.265 114.100 98.435 ;
        RECT 113.770 97.725 114.100 97.895 ;
        RECT 113.770 96.175 114.100 96.345 ;
        RECT 113.770 95.635 114.100 95.805 ;
        RECT 113.770 94.085 114.100 94.255 ;
        RECT 113.770 93.545 114.100 93.715 ;
        RECT 113.770 91.995 114.100 92.165 ;
        RECT 113.770 91.455 114.100 91.625 ;
        RECT 113.770 89.905 114.100 90.075 ;
        RECT 113.770 89.365 114.100 89.535 ;
        RECT 113.770 87.815 114.100 87.985 ;
        RECT 113.770 87.275 114.100 87.445 ;
        RECT 113.770 85.725 114.100 85.895 ;
        RECT 114.460 85.555 114.685 99.785 ;
        RECT 115.060 98.265 115.390 98.435 ;
        RECT 115.060 97.725 115.390 97.895 ;
        RECT 115.060 96.175 115.390 96.345 ;
        RECT 115.060 95.635 115.390 95.805 ;
        RECT 115.060 94.085 115.390 94.255 ;
        RECT 115.060 93.545 115.390 93.715 ;
        RECT 115.060 91.995 115.390 92.165 ;
        RECT 115.060 91.455 115.390 91.625 ;
        RECT 115.060 89.905 115.390 90.075 ;
        RECT 115.060 89.365 115.390 89.535 ;
        RECT 115.060 87.815 115.390 87.985 ;
        RECT 115.060 87.275 115.390 87.445 ;
        RECT 115.060 85.725 115.390 85.895 ;
        RECT 115.760 85.555 115.985 99.785 ;
        RECT 116.350 98.265 116.680 98.435 ;
        RECT 116.350 97.725 116.680 97.895 ;
        RECT 116.350 96.175 116.680 96.345 ;
        RECT 116.350 95.635 116.680 95.805 ;
        RECT 116.350 94.085 116.680 94.255 ;
        RECT 116.350 93.545 116.680 93.715 ;
        RECT 116.350 91.995 116.680 92.165 ;
        RECT 116.350 91.455 116.680 91.625 ;
        RECT 116.350 89.905 116.680 90.075 ;
        RECT 116.350 89.365 116.680 89.535 ;
        RECT 116.350 87.815 116.680 87.985 ;
        RECT 116.350 87.275 116.680 87.445 ;
        RECT 116.350 85.725 116.680 85.895 ;
        RECT 117.050 85.555 117.275 99.785 ;
        RECT 117.640 98.265 117.970 98.435 ;
        RECT 117.640 97.725 117.970 97.895 ;
        RECT 117.640 96.175 117.970 96.345 ;
        RECT 117.640 95.635 117.970 95.805 ;
        RECT 117.640 94.085 117.970 94.255 ;
        RECT 117.640 93.545 117.970 93.715 ;
        RECT 117.640 91.995 117.970 92.165 ;
        RECT 117.640 91.455 117.970 91.625 ;
        RECT 117.640 89.905 117.970 90.075 ;
        RECT 117.640 89.365 117.970 89.535 ;
        RECT 117.640 87.815 117.970 87.985 ;
        RECT 117.640 87.275 117.970 87.445 ;
        RECT 117.640 85.725 117.970 85.895 ;
        RECT 118.335 85.555 118.560 99.785 ;
        RECT 118.930 98.265 119.260 98.435 ;
        RECT 118.930 97.725 119.260 97.895 ;
        RECT 118.930 96.175 119.260 96.345 ;
        RECT 118.930 95.635 119.260 95.805 ;
        RECT 118.930 94.085 119.260 94.255 ;
        RECT 118.930 93.545 119.260 93.715 ;
        RECT 118.930 91.995 119.260 92.165 ;
        RECT 118.930 91.455 119.260 91.625 ;
        RECT 118.930 89.905 119.260 90.075 ;
        RECT 118.930 89.365 119.260 89.535 ;
        RECT 118.930 87.815 119.260 87.985 ;
        RECT 118.930 87.275 119.260 87.445 ;
        RECT 118.930 85.725 119.260 85.895 ;
        RECT 119.620 85.555 119.845 99.785 ;
        RECT 120.220 98.265 120.550 98.435 ;
        RECT 120.220 97.725 120.550 97.895 ;
        RECT 120.220 96.175 120.550 96.345 ;
        RECT 120.220 95.635 120.550 95.805 ;
        RECT 120.220 94.085 120.550 94.255 ;
        RECT 120.220 93.545 120.550 93.715 ;
        RECT 120.220 91.995 120.550 92.165 ;
        RECT 120.220 91.455 120.550 91.625 ;
        RECT 120.220 89.905 120.550 90.075 ;
        RECT 120.220 89.365 120.550 89.535 ;
        RECT 120.220 87.815 120.550 87.985 ;
        RECT 120.220 87.275 120.550 87.445 ;
        RECT 120.220 85.725 120.550 85.895 ;
        RECT 120.915 85.555 121.140 99.785 ;
        RECT 121.510 98.265 121.840 98.435 ;
        RECT 121.510 97.725 121.840 97.895 ;
        RECT 121.510 96.175 121.840 96.345 ;
        RECT 121.510 95.635 121.840 95.805 ;
        RECT 121.510 94.085 121.840 94.255 ;
        RECT 121.510 93.545 121.840 93.715 ;
        RECT 121.510 91.995 121.840 92.165 ;
        RECT 121.510 91.455 121.840 91.625 ;
        RECT 121.510 89.905 121.840 90.075 ;
        RECT 121.510 89.365 121.840 89.535 ;
        RECT 121.510 87.815 121.840 87.985 ;
        RECT 121.510 87.275 121.840 87.445 ;
        RECT 121.510 85.725 121.840 85.895 ;
        RECT 122.205 85.800 122.430 99.850 ;
        RECT 125.830 99.815 126.160 99.985 ;
        RECT 127.120 99.815 127.450 99.985 ;
        RECT 128.410 99.815 128.740 99.985 ;
        RECT 129.700 99.815 130.030 99.985 ;
        RECT 130.990 99.815 131.320 99.985 ;
        RECT 132.280 99.815 132.610 99.985 ;
        RECT 133.570 99.815 133.900 99.985 ;
        RECT 134.860 99.815 135.190 99.985 ;
        RECT 125.830 98.265 126.160 98.435 ;
        RECT 125.830 97.725 126.160 97.895 ;
        RECT 125.830 96.175 126.160 96.345 ;
        RECT 125.830 95.635 126.160 95.805 ;
        RECT 125.830 94.085 126.160 94.255 ;
        RECT 125.830 93.545 126.160 93.715 ;
        RECT 125.830 91.995 126.160 92.165 ;
        RECT 125.830 91.455 126.160 91.625 ;
        RECT 125.830 89.905 126.160 90.075 ;
        RECT 125.830 89.365 126.160 89.535 ;
        RECT 125.830 87.815 126.160 87.985 ;
        RECT 125.830 87.275 126.160 87.445 ;
        RECT 122.170 85.270 122.460 85.800 ;
        RECT 125.830 85.725 126.160 85.895 ;
        RECT 126.525 85.555 126.750 99.785 ;
        RECT 127.120 98.265 127.450 98.435 ;
        RECT 127.120 97.725 127.450 97.895 ;
        RECT 127.120 96.175 127.450 96.345 ;
        RECT 127.120 95.635 127.450 95.805 ;
        RECT 127.120 94.085 127.450 94.255 ;
        RECT 127.120 93.545 127.450 93.715 ;
        RECT 127.120 91.995 127.450 92.165 ;
        RECT 127.120 91.455 127.450 91.625 ;
        RECT 127.120 89.905 127.450 90.075 ;
        RECT 127.120 89.365 127.450 89.535 ;
        RECT 127.120 87.815 127.450 87.985 ;
        RECT 127.120 87.275 127.450 87.445 ;
        RECT 127.120 85.725 127.450 85.895 ;
        RECT 127.810 85.555 128.035 99.785 ;
        RECT 128.410 98.265 128.740 98.435 ;
        RECT 128.410 97.725 128.740 97.895 ;
        RECT 128.410 96.175 128.740 96.345 ;
        RECT 128.410 95.635 128.740 95.805 ;
        RECT 128.410 94.085 128.740 94.255 ;
        RECT 128.410 93.545 128.740 93.715 ;
        RECT 128.410 91.995 128.740 92.165 ;
        RECT 128.410 91.455 128.740 91.625 ;
        RECT 128.410 89.905 128.740 90.075 ;
        RECT 128.410 89.365 128.740 89.535 ;
        RECT 128.410 87.815 128.740 87.985 ;
        RECT 128.410 87.275 128.740 87.445 ;
        RECT 128.410 85.725 128.740 85.895 ;
        RECT 129.110 85.555 129.335 99.785 ;
        RECT 129.700 98.265 130.030 98.435 ;
        RECT 129.700 97.725 130.030 97.895 ;
        RECT 129.700 96.175 130.030 96.345 ;
        RECT 129.700 95.635 130.030 95.805 ;
        RECT 129.700 94.085 130.030 94.255 ;
        RECT 129.700 93.545 130.030 93.715 ;
        RECT 129.700 91.995 130.030 92.165 ;
        RECT 129.700 91.455 130.030 91.625 ;
        RECT 129.700 89.905 130.030 90.075 ;
        RECT 129.700 89.365 130.030 89.535 ;
        RECT 129.700 87.815 130.030 87.985 ;
        RECT 129.700 87.275 130.030 87.445 ;
        RECT 129.700 85.725 130.030 85.895 ;
        RECT 130.400 85.555 130.625 99.785 ;
        RECT 130.990 98.265 131.320 98.435 ;
        RECT 130.990 97.725 131.320 97.895 ;
        RECT 130.990 96.175 131.320 96.345 ;
        RECT 130.990 95.635 131.320 95.805 ;
        RECT 130.990 94.085 131.320 94.255 ;
        RECT 130.990 93.545 131.320 93.715 ;
        RECT 130.990 91.995 131.320 92.165 ;
        RECT 130.990 91.455 131.320 91.625 ;
        RECT 130.990 89.905 131.320 90.075 ;
        RECT 130.990 89.365 131.320 89.535 ;
        RECT 130.990 87.815 131.320 87.985 ;
        RECT 130.990 87.275 131.320 87.445 ;
        RECT 130.990 85.725 131.320 85.895 ;
        RECT 131.685 85.555 131.910 99.785 ;
        RECT 132.280 98.265 132.610 98.435 ;
        RECT 132.280 97.725 132.610 97.895 ;
        RECT 132.280 96.175 132.610 96.345 ;
        RECT 132.280 95.635 132.610 95.805 ;
        RECT 132.280 94.085 132.610 94.255 ;
        RECT 132.280 93.545 132.610 93.715 ;
        RECT 132.280 91.995 132.610 92.165 ;
        RECT 132.280 91.455 132.610 91.625 ;
        RECT 132.280 89.905 132.610 90.075 ;
        RECT 132.280 89.365 132.610 89.535 ;
        RECT 132.280 87.815 132.610 87.985 ;
        RECT 132.280 87.275 132.610 87.445 ;
        RECT 132.280 85.725 132.610 85.895 ;
        RECT 132.970 85.555 133.195 99.785 ;
        RECT 133.570 98.265 133.900 98.435 ;
        RECT 133.570 97.725 133.900 97.895 ;
        RECT 133.570 96.175 133.900 96.345 ;
        RECT 133.570 95.635 133.900 95.805 ;
        RECT 133.570 94.085 133.900 94.255 ;
        RECT 133.570 93.545 133.900 93.715 ;
        RECT 133.570 91.995 133.900 92.165 ;
        RECT 133.570 91.455 133.900 91.625 ;
        RECT 133.570 89.905 133.900 90.075 ;
        RECT 133.570 89.365 133.900 89.535 ;
        RECT 133.570 87.815 133.900 87.985 ;
        RECT 133.570 87.275 133.900 87.445 ;
        RECT 133.570 85.725 133.900 85.895 ;
        RECT 134.265 85.555 134.490 99.785 ;
        RECT 134.860 98.265 135.190 98.435 ;
        RECT 134.860 97.725 135.190 97.895 ;
        RECT 134.860 96.175 135.190 96.345 ;
        RECT 134.860 95.635 135.190 95.805 ;
        RECT 134.860 94.085 135.190 94.255 ;
        RECT 134.860 93.545 135.190 93.715 ;
        RECT 134.860 91.995 135.190 92.165 ;
        RECT 134.860 91.455 135.190 91.625 ;
        RECT 134.860 89.905 135.190 90.075 ;
        RECT 134.860 89.365 135.190 89.535 ;
        RECT 134.860 87.815 135.190 87.985 ;
        RECT 134.860 87.275 135.190 87.445 ;
        RECT 134.860 85.725 135.190 85.895 ;
        RECT 135.555 85.790 135.780 99.860 ;
        RECT 139.145 99.820 139.475 99.990 ;
        RECT 140.435 99.820 140.765 99.990 ;
        RECT 141.725 99.820 142.055 99.990 ;
        RECT 143.015 99.820 143.345 99.990 ;
        RECT 144.305 99.820 144.635 99.990 ;
        RECT 145.595 99.820 145.925 99.990 ;
        RECT 146.885 99.820 147.215 99.990 ;
        RECT 148.175 99.820 148.505 99.990 ;
        RECT 139.145 98.270 139.475 98.440 ;
        RECT 139.145 97.730 139.475 97.900 ;
        RECT 139.145 96.180 139.475 96.350 ;
        RECT 139.145 95.640 139.475 95.810 ;
        RECT 139.145 94.090 139.475 94.260 ;
        RECT 139.145 93.550 139.475 93.720 ;
        RECT 139.145 92.000 139.475 92.170 ;
        RECT 139.145 91.460 139.475 91.630 ;
        RECT 139.145 89.910 139.475 90.080 ;
        RECT 139.145 89.370 139.475 89.540 ;
        RECT 139.145 87.820 139.475 87.990 ;
        RECT 139.145 87.280 139.475 87.450 ;
        RECT 115.840 84.860 122.550 85.270 ;
        RECT 135.550 85.260 135.800 85.790 ;
        RECT 139.145 85.730 139.475 85.900 ;
        RECT 139.840 85.560 140.065 99.790 ;
        RECT 140.435 98.270 140.765 98.440 ;
        RECT 140.435 97.730 140.765 97.900 ;
        RECT 140.435 96.180 140.765 96.350 ;
        RECT 140.435 95.640 140.765 95.810 ;
        RECT 140.435 94.090 140.765 94.260 ;
        RECT 140.435 93.550 140.765 93.720 ;
        RECT 140.435 92.000 140.765 92.170 ;
        RECT 140.435 91.460 140.765 91.630 ;
        RECT 140.435 89.910 140.765 90.080 ;
        RECT 140.435 89.370 140.765 89.540 ;
        RECT 140.435 87.820 140.765 87.990 ;
        RECT 140.435 87.280 140.765 87.450 ;
        RECT 140.435 85.730 140.765 85.900 ;
        RECT 141.125 85.560 141.350 99.790 ;
        RECT 141.725 98.270 142.055 98.440 ;
        RECT 141.725 97.730 142.055 97.900 ;
        RECT 141.725 96.180 142.055 96.350 ;
        RECT 141.725 95.640 142.055 95.810 ;
        RECT 141.725 94.090 142.055 94.260 ;
        RECT 141.725 93.550 142.055 93.720 ;
        RECT 141.725 92.000 142.055 92.170 ;
        RECT 141.725 91.460 142.055 91.630 ;
        RECT 141.725 89.910 142.055 90.080 ;
        RECT 141.725 89.370 142.055 89.540 ;
        RECT 141.725 87.820 142.055 87.990 ;
        RECT 141.725 87.280 142.055 87.450 ;
        RECT 141.725 85.730 142.055 85.900 ;
        RECT 142.425 85.560 142.650 99.790 ;
        RECT 143.015 98.270 143.345 98.440 ;
        RECT 143.015 97.730 143.345 97.900 ;
        RECT 143.015 96.180 143.345 96.350 ;
        RECT 143.015 95.640 143.345 95.810 ;
        RECT 143.015 94.090 143.345 94.260 ;
        RECT 143.015 93.550 143.345 93.720 ;
        RECT 143.015 92.000 143.345 92.170 ;
        RECT 143.015 91.460 143.345 91.630 ;
        RECT 143.015 89.910 143.345 90.080 ;
        RECT 143.015 89.370 143.345 89.540 ;
        RECT 143.015 87.820 143.345 87.990 ;
        RECT 143.015 87.280 143.345 87.450 ;
        RECT 143.015 85.730 143.345 85.900 ;
        RECT 143.715 85.560 143.940 99.790 ;
        RECT 144.305 98.270 144.635 98.440 ;
        RECT 144.305 97.730 144.635 97.900 ;
        RECT 144.305 96.180 144.635 96.350 ;
        RECT 144.305 95.640 144.635 95.810 ;
        RECT 144.305 94.090 144.635 94.260 ;
        RECT 144.305 93.550 144.635 93.720 ;
        RECT 144.305 92.000 144.635 92.170 ;
        RECT 144.305 91.460 144.635 91.630 ;
        RECT 144.305 89.910 144.635 90.080 ;
        RECT 144.305 89.370 144.635 89.540 ;
        RECT 144.305 87.820 144.635 87.990 ;
        RECT 144.305 87.280 144.635 87.450 ;
        RECT 144.305 85.730 144.635 85.900 ;
        RECT 145.000 85.560 145.225 99.790 ;
        RECT 145.595 98.270 145.925 98.440 ;
        RECT 145.595 97.730 145.925 97.900 ;
        RECT 145.595 96.180 145.925 96.350 ;
        RECT 145.595 95.640 145.925 95.810 ;
        RECT 145.595 94.090 145.925 94.260 ;
        RECT 145.595 93.550 145.925 93.720 ;
        RECT 145.595 92.000 145.925 92.170 ;
        RECT 145.595 91.460 145.925 91.630 ;
        RECT 145.595 89.910 145.925 90.080 ;
        RECT 145.595 89.370 145.925 89.540 ;
        RECT 145.595 87.820 145.925 87.990 ;
        RECT 145.595 87.280 145.925 87.450 ;
        RECT 145.595 85.730 145.925 85.900 ;
        RECT 146.285 85.560 146.510 99.790 ;
        RECT 146.885 98.270 147.215 98.440 ;
        RECT 146.885 97.730 147.215 97.900 ;
        RECT 146.885 96.180 147.215 96.350 ;
        RECT 146.885 95.640 147.215 95.810 ;
        RECT 146.885 94.090 147.215 94.260 ;
        RECT 146.885 93.550 147.215 93.720 ;
        RECT 146.885 92.000 147.215 92.170 ;
        RECT 146.885 91.460 147.215 91.630 ;
        RECT 146.885 89.910 147.215 90.080 ;
        RECT 146.885 89.370 147.215 89.540 ;
        RECT 146.885 87.820 147.215 87.990 ;
        RECT 146.885 87.280 147.215 87.450 ;
        RECT 146.885 85.730 147.215 85.900 ;
        RECT 147.580 85.560 147.805 99.790 ;
        RECT 148.175 98.270 148.505 98.440 ;
        RECT 148.175 97.730 148.505 97.900 ;
        RECT 148.175 96.180 148.505 96.350 ;
        RECT 148.175 95.640 148.505 95.810 ;
        RECT 148.175 94.090 148.505 94.260 ;
        RECT 148.175 93.550 148.505 93.720 ;
        RECT 148.175 92.000 148.505 92.170 ;
        RECT 148.175 91.460 148.505 91.630 ;
        RECT 148.175 89.910 148.505 90.080 ;
        RECT 148.175 89.370 148.505 89.540 ;
        RECT 148.175 87.820 148.505 87.990 ;
        RECT 148.175 87.280 148.505 87.450 ;
        RECT 148.175 85.730 148.505 85.900 ;
        RECT 148.870 85.730 149.095 99.860 ;
        RECT 130.540 85.140 135.800 85.260 ;
        RECT 148.860 85.150 149.110 85.730 ;
        RECT 115.860 83.140 116.200 84.860 ;
        RECT 130.520 84.780 135.800 85.140 ;
        RECT 116.390 83.830 116.970 84.000 ;
        RECT 117.170 83.230 117.490 83.610 ;
        RECT 130.520 83.260 130.840 84.780 ;
        RECT 143.130 84.670 149.130 85.150 ;
        RECT 143.080 84.450 149.130 84.670 ;
        RECT 131.050 83.870 131.630 84.040 ;
        RECT 143.080 84.030 143.380 84.450 ;
        RECT 131.790 83.270 132.190 83.670 ;
        RECT 143.100 83.240 143.350 84.030 ;
        RECT 143.610 83.870 144.190 84.040 ;
        RECT 144.460 83.610 144.630 83.635 ;
        RECT 144.420 83.260 144.700 83.610 ;
        RECT 116.390 82.860 116.970 83.030 ;
        RECT 131.050 82.900 131.630 83.070 ;
        RECT 143.610 82.900 144.190 83.070 ;
        RECT 108.770 80.935 150.415 80.940 ;
        RECT 151.285 80.935 152.035 100.360 ;
        RECT 156.830 94.955 163.450 102.335 ;
        RECT 156.530 94.785 163.450 94.955 ;
        RECT 156.830 87.405 163.450 94.785 ;
        RECT 156.530 87.235 163.450 87.405 ;
        RECT 108.770 80.340 152.035 80.935 ;
        RECT 97.800 79.680 104.715 79.850 ;
        RECT 97.800 72.300 104.445 79.680 ;
        RECT 108.770 78.810 109.520 80.340 ;
        RECT 108.770 77.140 109.530 78.810 ;
        RECT 114.670 77.690 114.990 80.340 ;
        RECT 128.020 77.830 128.340 80.340 ;
        RECT 97.800 72.130 104.715 72.300 ;
        RECT 97.800 64.750 104.445 72.130 ;
        RECT 97.800 64.580 104.715 64.750 ;
        RECT 97.800 57.200 104.445 64.580 ;
        RECT 97.800 57.030 104.715 57.200 ;
        RECT 97.800 49.650 104.445 57.030 ;
        RECT 108.770 52.050 109.520 77.140 ;
        RECT 114.590 75.650 115.060 77.690 ;
        RECT 115.870 76.715 117.950 76.885 ;
        RECT 118.900 75.430 119.370 76.360 ;
        RECT 127.930 75.760 128.700 77.830 ;
        RECT 141.330 77.670 141.650 80.340 ;
        RECT 149.050 80.335 152.035 80.340 ;
        RECT 151.285 78.890 152.035 80.335 ;
        RECT 156.830 79.855 163.450 87.235 ;
        RECT 156.530 79.685 163.450 79.855 ;
        RECT 129.580 76.835 131.660 77.005 ;
        RECT 132.400 76.400 132.950 76.440 ;
        RECT 132.400 75.790 135.150 76.400 ;
        RECT 115.870 75.075 117.950 75.245 ;
        RECT 118.890 74.360 120.320 75.430 ;
        RECT 129.580 75.195 131.660 75.365 ;
        RECT 118.900 74.320 119.390 74.360 ;
        RECT 119.030 72.960 119.390 74.320 ;
        RECT 132.400 74.230 132.950 75.790 ;
        RECT 141.130 75.600 141.900 77.670 ;
        RECT 142.760 76.875 144.840 77.045 ;
        RECT 151.280 76.980 152.040 78.890 ;
        RECT 145.600 76.450 146.200 76.460 ;
        RECT 142.760 75.235 144.840 75.405 ;
        RECT 145.510 74.380 146.280 76.450 ;
        RECT 110.500 72.780 122.440 72.960 ;
        RECT 110.470 72.365 122.440 72.780 ;
        RECT 132.430 72.670 132.790 74.230 ;
        RECT 132.430 72.640 135.790 72.670 ;
        RECT 145.740 72.640 146.020 74.380 ;
        RECT 110.465 71.910 122.440 72.365 ;
        RECT 110.470 71.870 122.440 71.910 ;
        RECT 110.500 71.860 122.440 71.870 ;
        RECT 111.540 71.800 122.440 71.860 ;
        RECT 122.200 71.710 122.430 71.800 ;
        RECT 123.990 71.690 135.790 72.640 ;
        RECT 137.160 71.750 149.690 72.640 ;
        RECT 137.160 71.740 148.800 71.750 ;
        RECT 149.220 71.740 149.690 71.750 ;
        RECT 145.740 71.710 148.800 71.740 ;
        RECT 123.990 71.680 135.780 71.690 ;
        RECT 112.480 71.230 112.810 71.400 ;
        RECT 113.770 71.230 114.100 71.400 ;
        RECT 115.060 71.230 115.390 71.400 ;
        RECT 116.350 71.230 116.680 71.400 ;
        RECT 117.640 71.230 117.970 71.400 ;
        RECT 118.930 71.230 119.260 71.400 ;
        RECT 120.220 71.230 120.550 71.400 ;
        RECT 121.510 71.230 121.840 71.400 ;
        RECT 112.480 69.680 112.810 69.850 ;
        RECT 112.480 69.140 112.810 69.310 ;
        RECT 112.480 67.590 112.810 67.760 ;
        RECT 112.480 67.050 112.810 67.220 ;
        RECT 112.480 65.500 112.810 65.670 ;
        RECT 112.480 64.960 112.810 65.130 ;
        RECT 112.480 63.410 112.810 63.580 ;
        RECT 112.480 62.870 112.810 63.040 ;
        RECT 112.480 61.320 112.810 61.490 ;
        RECT 112.480 60.780 112.810 60.950 ;
        RECT 112.480 59.230 112.810 59.400 ;
        RECT 112.480 58.690 112.810 58.860 ;
        RECT 112.480 57.140 112.810 57.310 ;
        RECT 113.175 56.970 113.400 71.200 ;
        RECT 113.770 69.680 114.100 69.850 ;
        RECT 113.770 69.140 114.100 69.310 ;
        RECT 113.770 67.590 114.100 67.760 ;
        RECT 113.770 67.050 114.100 67.220 ;
        RECT 113.770 65.500 114.100 65.670 ;
        RECT 113.770 64.960 114.100 65.130 ;
        RECT 113.770 63.410 114.100 63.580 ;
        RECT 113.770 62.870 114.100 63.040 ;
        RECT 113.770 61.320 114.100 61.490 ;
        RECT 113.770 60.780 114.100 60.950 ;
        RECT 113.770 59.230 114.100 59.400 ;
        RECT 113.770 58.690 114.100 58.860 ;
        RECT 113.770 57.140 114.100 57.310 ;
        RECT 114.460 56.970 114.685 71.200 ;
        RECT 115.060 69.680 115.390 69.850 ;
        RECT 115.060 69.140 115.390 69.310 ;
        RECT 115.060 67.590 115.390 67.760 ;
        RECT 115.060 67.050 115.390 67.220 ;
        RECT 115.060 65.500 115.390 65.670 ;
        RECT 115.060 64.960 115.390 65.130 ;
        RECT 115.060 63.410 115.390 63.580 ;
        RECT 115.060 62.870 115.390 63.040 ;
        RECT 115.060 61.320 115.390 61.490 ;
        RECT 115.060 60.780 115.390 60.950 ;
        RECT 115.060 59.230 115.390 59.400 ;
        RECT 115.060 58.690 115.390 58.860 ;
        RECT 115.060 57.140 115.390 57.310 ;
        RECT 115.760 56.970 115.985 71.200 ;
        RECT 116.350 69.680 116.680 69.850 ;
        RECT 116.350 69.140 116.680 69.310 ;
        RECT 116.350 67.590 116.680 67.760 ;
        RECT 116.350 67.050 116.680 67.220 ;
        RECT 116.350 65.500 116.680 65.670 ;
        RECT 116.350 64.960 116.680 65.130 ;
        RECT 116.350 63.410 116.680 63.580 ;
        RECT 116.350 62.870 116.680 63.040 ;
        RECT 116.350 61.320 116.680 61.490 ;
        RECT 116.350 60.780 116.680 60.950 ;
        RECT 116.350 59.230 116.680 59.400 ;
        RECT 116.350 58.690 116.680 58.860 ;
        RECT 116.350 57.140 116.680 57.310 ;
        RECT 117.050 56.970 117.275 71.200 ;
        RECT 117.640 69.680 117.970 69.850 ;
        RECT 117.640 69.140 117.970 69.310 ;
        RECT 117.640 67.590 117.970 67.760 ;
        RECT 117.640 67.050 117.970 67.220 ;
        RECT 117.640 65.500 117.970 65.670 ;
        RECT 117.640 64.960 117.970 65.130 ;
        RECT 117.640 63.410 117.970 63.580 ;
        RECT 117.640 62.870 117.970 63.040 ;
        RECT 117.640 61.320 117.970 61.490 ;
        RECT 117.640 60.780 117.970 60.950 ;
        RECT 117.640 59.230 117.970 59.400 ;
        RECT 117.640 58.690 117.970 58.860 ;
        RECT 117.640 57.140 117.970 57.310 ;
        RECT 118.335 56.970 118.560 71.200 ;
        RECT 118.930 69.680 119.260 69.850 ;
        RECT 118.930 69.140 119.260 69.310 ;
        RECT 118.930 67.590 119.260 67.760 ;
        RECT 118.930 67.050 119.260 67.220 ;
        RECT 118.930 65.500 119.260 65.670 ;
        RECT 118.930 64.960 119.260 65.130 ;
        RECT 118.930 63.410 119.260 63.580 ;
        RECT 118.930 62.870 119.260 63.040 ;
        RECT 118.930 61.320 119.260 61.490 ;
        RECT 118.930 60.780 119.260 60.950 ;
        RECT 118.930 59.230 119.260 59.400 ;
        RECT 118.930 58.690 119.260 58.860 ;
        RECT 118.930 57.140 119.260 57.310 ;
        RECT 119.620 56.970 119.845 71.200 ;
        RECT 120.220 69.680 120.550 69.850 ;
        RECT 120.220 69.140 120.550 69.310 ;
        RECT 120.220 67.590 120.550 67.760 ;
        RECT 120.220 67.050 120.550 67.220 ;
        RECT 120.220 65.500 120.550 65.670 ;
        RECT 120.220 64.960 120.550 65.130 ;
        RECT 120.220 63.410 120.550 63.580 ;
        RECT 120.220 62.870 120.550 63.040 ;
        RECT 120.220 61.320 120.550 61.490 ;
        RECT 120.220 60.780 120.550 60.950 ;
        RECT 120.220 59.230 120.550 59.400 ;
        RECT 120.220 58.690 120.550 58.860 ;
        RECT 120.220 57.140 120.550 57.310 ;
        RECT 120.915 56.970 121.140 71.200 ;
        RECT 122.200 71.020 122.430 71.370 ;
        RECT 125.830 71.230 126.160 71.400 ;
        RECT 127.120 71.230 127.450 71.400 ;
        RECT 128.410 71.230 128.740 71.400 ;
        RECT 129.700 71.230 130.030 71.400 ;
        RECT 130.990 71.230 131.320 71.400 ;
        RECT 132.280 71.230 132.610 71.400 ;
        RECT 133.570 71.230 133.900 71.400 ;
        RECT 134.860 71.230 135.190 71.400 ;
        RECT 121.510 69.680 121.840 69.850 ;
        RECT 121.510 69.140 121.840 69.310 ;
        RECT 121.510 67.590 121.840 67.760 ;
        RECT 121.510 67.050 121.840 67.220 ;
        RECT 121.510 65.500 121.840 65.670 ;
        RECT 121.510 64.960 121.840 65.130 ;
        RECT 121.510 63.410 121.840 63.580 ;
        RECT 121.510 62.870 121.840 63.040 ;
        RECT 121.510 61.320 121.840 61.490 ;
        RECT 121.510 60.780 121.840 60.950 ;
        RECT 121.510 59.230 121.840 59.400 ;
        RECT 121.510 58.690 121.840 58.860 ;
        RECT 122.205 58.320 122.430 71.020 ;
        RECT 125.830 69.680 126.160 69.850 ;
        RECT 125.830 69.140 126.160 69.310 ;
        RECT 125.830 67.590 126.160 67.760 ;
        RECT 125.830 67.050 126.160 67.220 ;
        RECT 125.830 65.500 126.160 65.670 ;
        RECT 125.830 64.960 126.160 65.130 ;
        RECT 125.830 63.410 126.160 63.580 ;
        RECT 125.830 62.870 126.160 63.040 ;
        RECT 125.830 61.320 126.160 61.490 ;
        RECT 125.830 60.780 126.160 60.950 ;
        RECT 125.830 59.230 126.160 59.400 ;
        RECT 125.830 58.690 126.160 58.860 ;
        RECT 121.510 57.140 121.840 57.310 ;
        RECT 122.160 56.640 122.550 58.320 ;
        RECT 125.830 57.140 126.160 57.310 ;
        RECT 126.525 56.970 126.750 71.200 ;
        RECT 127.120 69.680 127.450 69.850 ;
        RECT 127.120 69.140 127.450 69.310 ;
        RECT 127.120 67.590 127.450 67.760 ;
        RECT 127.120 67.050 127.450 67.220 ;
        RECT 127.120 65.500 127.450 65.670 ;
        RECT 127.120 64.960 127.450 65.130 ;
        RECT 127.120 63.410 127.450 63.580 ;
        RECT 127.120 62.870 127.450 63.040 ;
        RECT 127.120 61.320 127.450 61.490 ;
        RECT 127.120 60.780 127.450 60.950 ;
        RECT 127.120 59.230 127.450 59.400 ;
        RECT 127.120 58.690 127.450 58.860 ;
        RECT 127.120 57.140 127.450 57.310 ;
        RECT 127.810 56.970 128.035 71.200 ;
        RECT 128.410 69.680 128.740 69.850 ;
        RECT 128.410 69.140 128.740 69.310 ;
        RECT 128.410 67.590 128.740 67.760 ;
        RECT 128.410 67.050 128.740 67.220 ;
        RECT 128.410 65.500 128.740 65.670 ;
        RECT 128.410 64.960 128.740 65.130 ;
        RECT 128.410 63.410 128.740 63.580 ;
        RECT 128.410 62.870 128.740 63.040 ;
        RECT 128.410 61.320 128.740 61.490 ;
        RECT 128.410 60.780 128.740 60.950 ;
        RECT 128.410 59.230 128.740 59.400 ;
        RECT 128.410 58.690 128.740 58.860 ;
        RECT 128.410 57.140 128.740 57.310 ;
        RECT 129.110 56.970 129.335 71.200 ;
        RECT 129.700 69.680 130.030 69.850 ;
        RECT 129.700 69.140 130.030 69.310 ;
        RECT 129.700 67.590 130.030 67.760 ;
        RECT 129.700 67.050 130.030 67.220 ;
        RECT 129.700 65.500 130.030 65.670 ;
        RECT 129.700 64.960 130.030 65.130 ;
        RECT 129.700 63.410 130.030 63.580 ;
        RECT 129.700 62.870 130.030 63.040 ;
        RECT 129.700 61.320 130.030 61.490 ;
        RECT 129.700 60.780 130.030 60.950 ;
        RECT 129.700 59.230 130.030 59.400 ;
        RECT 129.700 58.690 130.030 58.860 ;
        RECT 129.700 57.140 130.030 57.310 ;
        RECT 130.400 56.970 130.625 71.200 ;
        RECT 130.990 69.680 131.320 69.850 ;
        RECT 130.990 69.140 131.320 69.310 ;
        RECT 130.990 67.590 131.320 67.760 ;
        RECT 130.990 67.050 131.320 67.220 ;
        RECT 130.990 65.500 131.320 65.670 ;
        RECT 130.990 64.960 131.320 65.130 ;
        RECT 130.990 63.410 131.320 63.580 ;
        RECT 130.990 62.870 131.320 63.040 ;
        RECT 130.990 61.320 131.320 61.490 ;
        RECT 130.990 60.780 131.320 60.950 ;
        RECT 130.990 59.230 131.320 59.400 ;
        RECT 130.990 58.690 131.320 58.860 ;
        RECT 130.990 57.140 131.320 57.310 ;
        RECT 131.685 56.970 131.910 71.200 ;
        RECT 132.280 69.680 132.610 69.850 ;
        RECT 132.280 69.140 132.610 69.310 ;
        RECT 132.280 67.590 132.610 67.760 ;
        RECT 132.280 67.050 132.610 67.220 ;
        RECT 132.280 65.500 132.610 65.670 ;
        RECT 132.280 64.960 132.610 65.130 ;
        RECT 132.280 63.410 132.610 63.580 ;
        RECT 132.280 62.870 132.610 63.040 ;
        RECT 132.280 61.320 132.610 61.490 ;
        RECT 132.280 60.780 132.610 60.950 ;
        RECT 132.280 59.230 132.610 59.400 ;
        RECT 132.280 58.690 132.610 58.860 ;
        RECT 132.280 57.140 132.610 57.310 ;
        RECT 132.970 56.970 133.195 71.200 ;
        RECT 133.570 69.680 133.900 69.850 ;
        RECT 133.570 69.140 133.900 69.310 ;
        RECT 133.570 67.590 133.900 67.760 ;
        RECT 133.570 67.050 133.900 67.220 ;
        RECT 133.570 65.500 133.900 65.670 ;
        RECT 133.570 64.960 133.900 65.130 ;
        RECT 133.570 63.410 133.900 63.580 ;
        RECT 133.570 62.870 133.900 63.040 ;
        RECT 133.570 61.320 133.900 61.490 ;
        RECT 133.570 60.780 133.900 60.950 ;
        RECT 133.570 59.230 133.900 59.400 ;
        RECT 133.570 58.690 133.900 58.860 ;
        RECT 133.570 57.140 133.900 57.310 ;
        RECT 134.265 56.970 134.490 71.200 ;
        RECT 135.560 71.080 135.780 71.260 ;
        RECT 139.145 71.235 139.475 71.405 ;
        RECT 140.435 71.235 140.765 71.405 ;
        RECT 141.725 71.235 142.055 71.405 ;
        RECT 143.015 71.235 143.345 71.405 ;
        RECT 144.305 71.235 144.635 71.405 ;
        RECT 145.595 71.235 145.925 71.405 ;
        RECT 146.885 71.235 147.215 71.405 ;
        RECT 148.175 71.235 148.505 71.405 ;
        RECT 148.870 71.230 149.060 71.270 ;
        RECT 134.860 69.680 135.190 69.850 ;
        RECT 134.860 69.140 135.190 69.310 ;
        RECT 134.860 67.590 135.190 67.760 ;
        RECT 134.860 67.050 135.190 67.220 ;
        RECT 134.860 65.500 135.190 65.670 ;
        RECT 134.860 64.960 135.190 65.130 ;
        RECT 134.860 63.410 135.190 63.580 ;
        RECT 134.860 62.870 135.190 63.040 ;
        RECT 134.860 61.320 135.190 61.490 ;
        RECT 134.860 60.780 135.190 60.950 ;
        RECT 134.860 59.230 135.190 59.400 ;
        RECT 134.860 58.690 135.190 58.860 ;
        RECT 135.555 57.790 135.780 71.080 ;
        RECT 139.145 69.685 139.475 69.855 ;
        RECT 139.145 69.145 139.475 69.315 ;
        RECT 139.145 67.595 139.475 67.765 ;
        RECT 139.145 67.055 139.475 67.225 ;
        RECT 139.145 65.505 139.475 65.675 ;
        RECT 139.145 64.965 139.475 65.135 ;
        RECT 139.145 63.415 139.475 63.585 ;
        RECT 139.145 62.875 139.475 63.045 ;
        RECT 139.145 61.325 139.475 61.495 ;
        RECT 139.145 60.785 139.475 60.955 ;
        RECT 139.145 59.235 139.475 59.405 ;
        RECT 139.145 58.695 139.475 58.865 ;
        RECT 134.860 57.140 135.190 57.310 ;
        RECT 115.820 56.320 122.650 56.640 ;
        RECT 115.820 55.080 116.060 56.320 ;
        RECT 129.970 56.210 130.360 56.280 ;
        RECT 135.510 56.210 135.900 57.790 ;
        RECT 139.145 57.145 139.475 57.315 ;
        RECT 139.840 56.975 140.065 71.205 ;
        RECT 140.435 69.685 140.765 69.855 ;
        RECT 140.435 69.145 140.765 69.315 ;
        RECT 140.435 67.595 140.765 67.765 ;
        RECT 140.435 67.055 140.765 67.225 ;
        RECT 140.435 65.505 140.765 65.675 ;
        RECT 140.435 64.965 140.765 65.135 ;
        RECT 140.435 63.415 140.765 63.585 ;
        RECT 140.435 62.875 140.765 63.045 ;
        RECT 140.435 61.325 140.765 61.495 ;
        RECT 140.435 60.785 140.765 60.955 ;
        RECT 140.435 59.235 140.765 59.405 ;
        RECT 140.435 58.695 140.765 58.865 ;
        RECT 140.435 57.145 140.765 57.315 ;
        RECT 141.125 56.975 141.350 71.205 ;
        RECT 141.725 69.685 142.055 69.855 ;
        RECT 141.725 69.145 142.055 69.315 ;
        RECT 141.725 67.595 142.055 67.765 ;
        RECT 141.725 67.055 142.055 67.225 ;
        RECT 141.725 65.505 142.055 65.675 ;
        RECT 141.725 64.965 142.055 65.135 ;
        RECT 141.725 63.415 142.055 63.585 ;
        RECT 141.725 62.875 142.055 63.045 ;
        RECT 141.725 61.325 142.055 61.495 ;
        RECT 141.725 60.785 142.055 60.955 ;
        RECT 141.725 59.235 142.055 59.405 ;
        RECT 141.725 58.695 142.055 58.865 ;
        RECT 141.725 57.145 142.055 57.315 ;
        RECT 142.425 56.975 142.650 71.205 ;
        RECT 143.015 69.685 143.345 69.855 ;
        RECT 143.015 69.145 143.345 69.315 ;
        RECT 143.015 67.595 143.345 67.765 ;
        RECT 143.015 67.055 143.345 67.225 ;
        RECT 143.015 65.505 143.345 65.675 ;
        RECT 143.015 64.965 143.345 65.135 ;
        RECT 143.015 63.415 143.345 63.585 ;
        RECT 143.015 62.875 143.345 63.045 ;
        RECT 143.015 61.325 143.345 61.495 ;
        RECT 143.015 60.785 143.345 60.955 ;
        RECT 143.015 59.235 143.345 59.405 ;
        RECT 143.015 58.695 143.345 58.865 ;
        RECT 143.015 57.145 143.345 57.315 ;
        RECT 143.715 56.975 143.940 71.205 ;
        RECT 144.305 69.685 144.635 69.855 ;
        RECT 144.305 69.145 144.635 69.315 ;
        RECT 144.305 67.595 144.635 67.765 ;
        RECT 144.305 67.055 144.635 67.225 ;
        RECT 144.305 65.505 144.635 65.675 ;
        RECT 144.305 64.965 144.635 65.135 ;
        RECT 144.305 63.415 144.635 63.585 ;
        RECT 144.305 62.875 144.635 63.045 ;
        RECT 144.305 61.325 144.635 61.495 ;
        RECT 144.305 60.785 144.635 60.955 ;
        RECT 144.305 59.235 144.635 59.405 ;
        RECT 144.305 58.695 144.635 58.865 ;
        RECT 144.305 57.145 144.635 57.315 ;
        RECT 145.000 56.975 145.225 71.205 ;
        RECT 145.595 69.685 145.925 69.855 ;
        RECT 145.595 69.145 145.925 69.315 ;
        RECT 145.595 67.595 145.925 67.765 ;
        RECT 145.595 67.055 145.925 67.225 ;
        RECT 145.595 65.505 145.925 65.675 ;
        RECT 145.595 64.965 145.925 65.135 ;
        RECT 145.595 63.415 145.925 63.585 ;
        RECT 145.595 62.875 145.925 63.045 ;
        RECT 145.595 61.325 145.925 61.495 ;
        RECT 145.595 60.785 145.925 60.955 ;
        RECT 145.595 59.235 145.925 59.405 ;
        RECT 145.595 58.695 145.925 58.865 ;
        RECT 145.595 57.145 145.925 57.315 ;
        RECT 146.285 56.975 146.510 71.205 ;
        RECT 146.885 69.685 147.215 69.855 ;
        RECT 146.885 69.145 147.215 69.315 ;
        RECT 146.885 67.595 147.215 67.765 ;
        RECT 146.885 67.055 147.215 67.225 ;
        RECT 146.885 65.505 147.215 65.675 ;
        RECT 146.885 64.965 147.215 65.135 ;
        RECT 146.885 63.415 147.215 63.585 ;
        RECT 146.885 62.875 147.215 63.045 ;
        RECT 146.885 61.325 147.215 61.495 ;
        RECT 146.885 60.785 147.215 60.955 ;
        RECT 146.885 59.235 147.215 59.405 ;
        RECT 146.885 58.695 147.215 58.865 ;
        RECT 146.885 57.145 147.215 57.315 ;
        RECT 147.580 56.975 147.805 71.205 ;
        RECT 148.870 71.060 149.100 71.230 ;
        RECT 148.175 69.685 148.505 69.855 ;
        RECT 148.175 69.145 148.505 69.315 ;
        RECT 148.175 67.595 148.505 67.765 ;
        RECT 148.175 67.055 148.505 67.225 ;
        RECT 148.175 65.505 148.505 65.675 ;
        RECT 148.175 64.965 148.505 65.135 ;
        RECT 148.175 63.415 148.505 63.585 ;
        RECT 148.175 62.875 148.505 63.045 ;
        RECT 148.175 61.325 148.505 61.495 ;
        RECT 148.175 60.785 148.505 60.955 ;
        RECT 148.175 59.235 148.505 59.405 ;
        RECT 148.175 58.695 148.505 58.865 ;
        RECT 148.870 57.900 149.095 71.060 ;
        RECT 148.175 57.145 148.505 57.315 ;
        RECT 142.120 56.300 142.510 56.320 ;
        RECT 148.850 56.300 149.240 57.900 ;
        RECT 151.285 57.660 152.035 76.980 ;
        RECT 156.830 72.305 163.450 79.685 ;
        RECT 156.530 72.135 163.450 72.305 ;
        RECT 156.830 64.755 163.450 72.135 ;
        RECT 156.530 64.585 163.450 64.755 ;
        RECT 129.970 55.820 135.970 56.210 ;
        RECT 142.120 55.930 149.240 56.300 ;
        RECT 142.120 55.900 149.220 55.930 ;
        RECT 116.300 55.290 116.880 55.460 ;
        RECT 115.780 54.670 116.160 55.080 ;
        RECT 117.070 54.550 117.380 55.080 ;
        RECT 116.300 54.320 116.880 54.490 ;
        RECT 129.970 54.310 130.360 55.820 ;
        RECT 130.580 55.000 131.160 55.170 ;
        RECT 131.380 54.280 131.690 54.810 ;
        RECT 142.120 54.350 142.510 55.900 ;
        RECT 142.690 54.980 143.270 55.150 ;
        RECT 143.480 54.310 143.790 54.840 ;
        RECT 130.580 54.030 131.160 54.200 ;
        RECT 142.690 54.010 143.270 54.180 ;
        RECT 151.280 52.050 152.040 57.660 ;
        RECT 156.830 57.205 163.450 64.585 ;
        RECT 156.530 57.035 163.450 57.205 ;
        RECT 108.770 51.430 152.040 52.050 ;
        RECT 97.800 49.480 104.715 49.650 ;
        RECT 97.800 42.100 104.445 49.480 ;
        RECT 114.670 47.880 114.990 51.430 ;
        RECT 128.010 48.410 128.330 51.430 ;
        RECT 114.670 47.610 115.180 47.880 ;
        RECT 114.680 46.170 115.180 47.610 ;
        RECT 116.150 47.245 118.230 47.415 ;
        RECT 127.950 47.080 128.460 48.410 ;
        RECT 141.340 48.290 141.660 51.430 ;
        RECT 156.830 49.655 163.450 57.035 ;
        RECT 156.530 49.485 163.450 49.655 ;
        RECT 129.850 47.485 131.930 47.655 ;
        RECT 132.750 47.090 133.260 47.150 ;
        RECT 118.880 45.880 119.860 46.980 ;
        RECT 127.950 46.440 128.900 47.080 ;
        RECT 116.150 45.605 118.230 45.775 ;
        RECT 119.160 45.390 119.590 45.880 ;
        RECT 129.850 45.845 131.930 46.015 ;
        RECT 132.730 45.390 133.260 47.090 ;
        RECT 141.190 46.220 141.960 48.290 ;
        RECT 142.530 47.255 144.610 47.425 ;
        RECT 142.530 45.615 144.610 45.785 ;
        RECT 145.400 45.440 146.170 47.070 ;
        RECT 119.160 45.140 119.670 45.390 ;
        RECT 132.390 45.340 133.260 45.390 ;
        RECT 132.380 45.180 133.260 45.340 ;
        RECT 132.380 45.170 133.240 45.180 ;
        RECT 119.290 42.925 119.670 45.140 ;
        RECT 132.390 45.120 133.240 45.170 ;
        RECT 132.390 45.110 132.900 45.120 ;
        RECT 132.440 43.110 132.670 45.110 ;
        RECT 132.440 42.925 132.665 43.110 ;
        RECT 119.290 42.400 130.795 42.925 ;
        RECT 119.290 42.390 122.445 42.400 ;
        RECT 129.480 42.395 130.795 42.400 ;
        RECT 132.440 42.400 144.085 42.925 ;
        RECT 132.440 42.390 135.520 42.400 ;
        RECT 142.845 42.395 144.085 42.400 ;
        RECT 145.380 42.920 146.170 45.440 ;
        RECT 148.830 44.310 150.300 44.320 ;
        RECT 148.830 42.920 150.560 44.310 ;
        RECT 145.380 42.400 150.560 42.920 ;
        RECT 152.170 42.640 153.420 44.090 ;
        RECT 145.380 42.395 150.415 42.400 ;
        RECT 119.290 42.360 119.670 42.390 ;
        RECT 145.380 42.380 146.170 42.395 ;
        RECT 148.850 42.390 149.095 42.395 ;
        RECT 156.830 42.105 163.450 49.485 ;
        RECT 97.800 41.930 104.715 42.100 ;
        RECT 97.800 34.550 104.445 41.930 ;
        RECT 112.480 41.710 112.810 41.880 ;
        RECT 113.770 41.710 114.100 41.880 ;
        RECT 115.060 41.710 115.390 41.880 ;
        RECT 116.350 41.710 116.680 41.880 ;
        RECT 117.640 41.710 117.970 41.880 ;
        RECT 118.930 41.710 119.260 41.880 ;
        RECT 120.220 41.710 120.550 41.880 ;
        RECT 121.510 41.710 121.840 41.880 ;
        RECT 112.480 40.160 112.810 40.330 ;
        RECT 112.480 39.620 112.810 39.790 ;
        RECT 112.480 38.070 112.810 38.240 ;
        RECT 112.480 37.530 112.810 37.700 ;
        RECT 112.480 35.980 112.810 36.150 ;
        RECT 112.480 35.440 112.810 35.610 ;
        RECT 97.800 34.380 104.715 34.550 ;
        RECT 97.800 27.000 104.445 34.380 ;
        RECT 112.480 33.890 112.810 34.060 ;
        RECT 112.480 33.350 112.810 33.520 ;
        RECT 112.480 31.800 112.810 31.970 ;
        RECT 112.480 31.260 112.810 31.430 ;
        RECT 112.480 29.710 112.810 29.880 ;
        RECT 112.480 29.170 112.810 29.340 ;
        RECT 112.480 27.620 112.810 27.790 ;
        RECT 113.175 27.450 113.400 41.680 ;
        RECT 113.770 40.160 114.100 40.330 ;
        RECT 113.770 39.620 114.100 39.790 ;
        RECT 113.770 38.070 114.100 38.240 ;
        RECT 113.770 37.530 114.100 37.700 ;
        RECT 113.770 35.980 114.100 36.150 ;
        RECT 113.770 35.440 114.100 35.610 ;
        RECT 113.770 33.890 114.100 34.060 ;
        RECT 113.770 33.350 114.100 33.520 ;
        RECT 113.770 31.800 114.100 31.970 ;
        RECT 113.770 31.260 114.100 31.430 ;
        RECT 113.770 29.710 114.100 29.880 ;
        RECT 113.770 29.170 114.100 29.340 ;
        RECT 113.770 27.620 114.100 27.790 ;
        RECT 114.460 27.450 114.685 41.680 ;
        RECT 115.060 40.160 115.390 40.330 ;
        RECT 115.060 39.620 115.390 39.790 ;
        RECT 115.060 38.070 115.390 38.240 ;
        RECT 115.060 37.530 115.390 37.700 ;
        RECT 115.060 35.980 115.390 36.150 ;
        RECT 115.060 35.440 115.390 35.610 ;
        RECT 115.060 33.890 115.390 34.060 ;
        RECT 115.060 33.350 115.390 33.520 ;
        RECT 115.060 31.800 115.390 31.970 ;
        RECT 115.060 31.260 115.390 31.430 ;
        RECT 115.060 29.710 115.390 29.880 ;
        RECT 115.060 29.170 115.390 29.340 ;
        RECT 115.060 27.620 115.390 27.790 ;
        RECT 115.760 27.450 115.985 41.680 ;
        RECT 116.350 40.160 116.680 40.330 ;
        RECT 116.350 39.620 116.680 39.790 ;
        RECT 116.350 38.070 116.680 38.240 ;
        RECT 116.350 37.530 116.680 37.700 ;
        RECT 116.350 35.980 116.680 36.150 ;
        RECT 116.350 35.440 116.680 35.610 ;
        RECT 116.350 33.890 116.680 34.060 ;
        RECT 116.350 33.350 116.680 33.520 ;
        RECT 116.350 31.800 116.680 31.970 ;
        RECT 116.350 31.260 116.680 31.430 ;
        RECT 116.350 29.710 116.680 29.880 ;
        RECT 116.350 29.170 116.680 29.340 ;
        RECT 116.350 27.620 116.680 27.790 ;
        RECT 117.050 27.450 117.275 41.680 ;
        RECT 117.640 40.160 117.970 40.330 ;
        RECT 117.640 39.620 117.970 39.790 ;
        RECT 117.640 38.070 117.970 38.240 ;
        RECT 117.640 37.530 117.970 37.700 ;
        RECT 117.640 35.980 117.970 36.150 ;
        RECT 117.640 35.440 117.970 35.610 ;
        RECT 117.640 33.890 117.970 34.060 ;
        RECT 117.640 33.350 117.970 33.520 ;
        RECT 117.640 31.800 117.970 31.970 ;
        RECT 117.640 31.260 117.970 31.430 ;
        RECT 117.640 29.710 117.970 29.880 ;
        RECT 117.640 29.170 117.970 29.340 ;
        RECT 117.640 27.620 117.970 27.790 ;
        RECT 118.335 27.450 118.560 41.680 ;
        RECT 118.930 40.160 119.260 40.330 ;
        RECT 118.930 39.620 119.260 39.790 ;
        RECT 118.930 38.070 119.260 38.240 ;
        RECT 118.930 37.530 119.260 37.700 ;
        RECT 118.930 35.980 119.260 36.150 ;
        RECT 118.930 35.440 119.260 35.610 ;
        RECT 118.930 33.890 119.260 34.060 ;
        RECT 118.930 33.350 119.260 33.520 ;
        RECT 118.930 31.800 119.260 31.970 ;
        RECT 118.930 31.260 119.260 31.430 ;
        RECT 118.930 29.710 119.260 29.880 ;
        RECT 118.930 29.170 119.260 29.340 ;
        RECT 118.930 27.620 119.260 27.790 ;
        RECT 119.620 27.450 119.845 41.680 ;
        RECT 120.220 40.160 120.550 40.330 ;
        RECT 120.220 39.620 120.550 39.790 ;
        RECT 120.220 38.070 120.550 38.240 ;
        RECT 120.220 37.530 120.550 37.700 ;
        RECT 120.220 35.980 120.550 36.150 ;
        RECT 120.220 35.440 120.550 35.610 ;
        RECT 120.220 33.890 120.550 34.060 ;
        RECT 120.220 33.350 120.550 33.520 ;
        RECT 120.220 31.800 120.550 31.970 ;
        RECT 120.220 31.260 120.550 31.430 ;
        RECT 120.220 29.710 120.550 29.880 ;
        RECT 120.220 29.170 120.550 29.340 ;
        RECT 120.220 27.620 120.550 27.790 ;
        RECT 120.915 27.450 121.140 41.680 ;
        RECT 121.510 40.160 121.840 40.330 ;
        RECT 121.510 39.620 121.840 39.790 ;
        RECT 121.510 38.070 121.840 38.240 ;
        RECT 121.510 37.530 121.840 37.700 ;
        RECT 121.510 35.980 121.840 36.150 ;
        RECT 121.510 35.440 121.840 35.610 ;
        RECT 121.510 33.890 121.840 34.060 ;
        RECT 121.510 33.350 121.840 33.520 ;
        RECT 121.510 31.800 121.840 31.970 ;
        RECT 121.510 31.260 121.840 31.430 ;
        RECT 121.510 29.710 121.840 29.880 ;
        RECT 121.510 29.170 121.840 29.340 ;
        RECT 121.510 27.620 121.840 27.790 ;
        RECT 122.205 27.710 122.430 42.070 ;
        RECT 156.530 41.935 163.450 42.105 ;
        RECT 125.830 41.710 126.160 41.880 ;
        RECT 127.120 41.710 127.450 41.880 ;
        RECT 128.410 41.710 128.740 41.880 ;
        RECT 129.700 41.710 130.030 41.880 ;
        RECT 130.990 41.710 131.320 41.880 ;
        RECT 132.280 41.710 132.610 41.880 ;
        RECT 133.570 41.710 133.900 41.880 ;
        RECT 134.860 41.710 135.190 41.880 ;
        RECT 125.830 40.160 126.160 40.330 ;
        RECT 125.830 39.620 126.160 39.790 ;
        RECT 125.830 38.070 126.160 38.240 ;
        RECT 125.830 37.530 126.160 37.700 ;
        RECT 125.830 35.980 126.160 36.150 ;
        RECT 125.830 35.440 126.160 35.610 ;
        RECT 125.830 33.890 126.160 34.060 ;
        RECT 125.830 33.350 126.160 33.520 ;
        RECT 125.830 31.800 126.160 31.970 ;
        RECT 125.830 31.260 126.160 31.430 ;
        RECT 125.830 29.710 126.160 29.880 ;
        RECT 125.830 29.170 126.160 29.340 ;
        RECT 97.800 26.830 104.715 27.000 ;
        RECT 115.750 26.850 116.080 26.880 ;
        RECT 122.170 26.850 122.470 27.710 ;
        RECT 125.830 27.620 126.160 27.790 ;
        RECT 126.525 27.450 126.750 41.680 ;
        RECT 127.120 40.160 127.450 40.330 ;
        RECT 127.120 39.620 127.450 39.790 ;
        RECT 127.120 38.070 127.450 38.240 ;
        RECT 127.120 37.530 127.450 37.700 ;
        RECT 127.120 35.980 127.450 36.150 ;
        RECT 127.120 35.440 127.450 35.610 ;
        RECT 127.120 33.890 127.450 34.060 ;
        RECT 127.120 33.350 127.450 33.520 ;
        RECT 127.120 31.800 127.450 31.970 ;
        RECT 127.120 31.260 127.450 31.430 ;
        RECT 127.120 29.710 127.450 29.880 ;
        RECT 127.120 29.170 127.450 29.340 ;
        RECT 127.120 27.620 127.450 27.790 ;
        RECT 127.810 27.450 128.035 41.680 ;
        RECT 128.410 40.160 128.740 40.330 ;
        RECT 128.410 39.620 128.740 39.790 ;
        RECT 128.410 38.070 128.740 38.240 ;
        RECT 128.410 37.530 128.740 37.700 ;
        RECT 128.410 35.980 128.740 36.150 ;
        RECT 128.410 35.440 128.740 35.610 ;
        RECT 128.410 33.890 128.740 34.060 ;
        RECT 128.410 33.350 128.740 33.520 ;
        RECT 128.410 31.800 128.740 31.970 ;
        RECT 128.410 31.260 128.740 31.430 ;
        RECT 128.410 29.710 128.740 29.880 ;
        RECT 128.410 29.170 128.740 29.340 ;
        RECT 128.410 27.620 128.740 27.790 ;
        RECT 129.110 27.450 129.335 41.680 ;
        RECT 129.700 40.160 130.030 40.330 ;
        RECT 129.700 39.620 130.030 39.790 ;
        RECT 129.700 38.070 130.030 38.240 ;
        RECT 129.700 37.530 130.030 37.700 ;
        RECT 129.700 35.980 130.030 36.150 ;
        RECT 129.700 35.440 130.030 35.610 ;
        RECT 129.700 33.890 130.030 34.060 ;
        RECT 129.700 33.350 130.030 33.520 ;
        RECT 129.700 31.800 130.030 31.970 ;
        RECT 129.700 31.260 130.030 31.430 ;
        RECT 129.700 29.710 130.030 29.880 ;
        RECT 129.700 29.170 130.030 29.340 ;
        RECT 129.700 27.620 130.030 27.790 ;
        RECT 130.400 27.450 130.625 41.680 ;
        RECT 130.990 40.160 131.320 40.330 ;
        RECT 130.990 39.620 131.320 39.790 ;
        RECT 130.990 38.070 131.320 38.240 ;
        RECT 130.990 37.530 131.320 37.700 ;
        RECT 130.990 35.980 131.320 36.150 ;
        RECT 130.990 35.440 131.320 35.610 ;
        RECT 130.990 33.890 131.320 34.060 ;
        RECT 130.990 33.350 131.320 33.520 ;
        RECT 130.990 31.800 131.320 31.970 ;
        RECT 130.990 31.260 131.320 31.430 ;
        RECT 130.990 29.710 131.320 29.880 ;
        RECT 130.990 29.170 131.320 29.340 ;
        RECT 130.990 27.620 131.320 27.790 ;
        RECT 131.685 27.450 131.910 41.680 ;
        RECT 132.280 40.160 132.610 40.330 ;
        RECT 132.280 39.620 132.610 39.790 ;
        RECT 132.280 38.070 132.610 38.240 ;
        RECT 132.280 37.530 132.610 37.700 ;
        RECT 132.280 35.980 132.610 36.150 ;
        RECT 132.280 35.440 132.610 35.610 ;
        RECT 132.280 33.890 132.610 34.060 ;
        RECT 132.280 33.350 132.610 33.520 ;
        RECT 132.280 31.800 132.610 31.970 ;
        RECT 132.280 31.260 132.610 31.430 ;
        RECT 132.280 29.710 132.610 29.880 ;
        RECT 132.280 29.170 132.610 29.340 ;
        RECT 132.280 27.620 132.610 27.790 ;
        RECT 132.970 27.450 133.195 41.680 ;
        RECT 133.570 40.160 133.900 40.330 ;
        RECT 133.570 39.620 133.900 39.790 ;
        RECT 133.570 38.070 133.900 38.240 ;
        RECT 133.570 37.530 133.900 37.700 ;
        RECT 133.570 35.980 133.900 36.150 ;
        RECT 133.570 35.440 133.900 35.610 ;
        RECT 133.570 33.890 133.900 34.060 ;
        RECT 133.570 33.350 133.900 33.520 ;
        RECT 133.570 31.800 133.900 31.970 ;
        RECT 133.570 31.260 133.900 31.430 ;
        RECT 133.570 29.710 133.900 29.880 ;
        RECT 133.570 29.170 133.900 29.340 ;
        RECT 133.570 27.620 133.900 27.790 ;
        RECT 134.265 27.450 134.490 41.680 ;
        RECT 134.860 40.160 135.190 40.330 ;
        RECT 134.860 39.620 135.190 39.790 ;
        RECT 134.860 38.070 135.190 38.240 ;
        RECT 134.860 37.530 135.190 37.700 ;
        RECT 134.860 35.980 135.190 36.150 ;
        RECT 134.860 35.440 135.190 35.610 ;
        RECT 134.860 33.890 135.190 34.060 ;
        RECT 134.860 33.350 135.190 33.520 ;
        RECT 134.860 31.800 135.190 31.970 ;
        RECT 134.860 31.260 135.190 31.430 ;
        RECT 134.860 29.710 135.190 29.880 ;
        RECT 134.860 29.170 135.190 29.340 ;
        RECT 135.555 27.810 135.780 41.880 ;
        RECT 139.145 41.715 139.475 41.885 ;
        RECT 140.435 41.715 140.765 41.885 ;
        RECT 141.725 41.715 142.055 41.885 ;
        RECT 143.015 41.715 143.345 41.885 ;
        RECT 144.305 41.715 144.635 41.885 ;
        RECT 145.595 41.715 145.925 41.885 ;
        RECT 146.885 41.715 147.215 41.885 ;
        RECT 148.175 41.715 148.505 41.885 ;
        RECT 139.145 40.165 139.475 40.335 ;
        RECT 139.145 39.625 139.475 39.795 ;
        RECT 139.145 38.075 139.475 38.245 ;
        RECT 139.145 37.535 139.475 37.705 ;
        RECT 139.145 35.985 139.475 36.155 ;
        RECT 139.145 35.445 139.475 35.615 ;
        RECT 139.145 33.895 139.475 34.065 ;
        RECT 139.145 33.355 139.475 33.525 ;
        RECT 139.145 31.805 139.475 31.975 ;
        RECT 139.145 31.265 139.475 31.435 ;
        RECT 139.145 29.715 139.475 29.885 ;
        RECT 139.145 29.175 139.475 29.345 ;
        RECT 134.860 27.620 135.190 27.790 ;
        RECT 97.800 19.450 104.445 26.830 ;
        RECT 115.750 26.490 122.470 26.850 ;
        RECT 135.480 26.660 135.800 27.810 ;
        RECT 139.145 27.625 139.475 27.795 ;
        RECT 139.840 27.455 140.065 41.685 ;
        RECT 140.435 40.165 140.765 40.335 ;
        RECT 140.435 39.625 140.765 39.795 ;
        RECT 140.435 38.075 140.765 38.245 ;
        RECT 140.435 37.535 140.765 37.705 ;
        RECT 140.435 35.985 140.765 36.155 ;
        RECT 140.435 35.445 140.765 35.615 ;
        RECT 140.435 33.895 140.765 34.065 ;
        RECT 140.435 33.355 140.765 33.525 ;
        RECT 140.435 31.805 140.765 31.975 ;
        RECT 140.435 31.265 140.765 31.435 ;
        RECT 140.435 29.715 140.765 29.885 ;
        RECT 140.435 29.175 140.765 29.345 ;
        RECT 140.435 27.625 140.765 27.795 ;
        RECT 141.125 27.455 141.350 41.685 ;
        RECT 141.725 40.165 142.055 40.335 ;
        RECT 141.725 39.625 142.055 39.795 ;
        RECT 141.725 38.075 142.055 38.245 ;
        RECT 141.725 37.535 142.055 37.705 ;
        RECT 141.725 35.985 142.055 36.155 ;
        RECT 141.725 35.445 142.055 35.615 ;
        RECT 141.725 33.895 142.055 34.065 ;
        RECT 141.725 33.355 142.055 33.525 ;
        RECT 141.725 31.805 142.055 31.975 ;
        RECT 141.725 31.265 142.055 31.435 ;
        RECT 141.725 29.715 142.055 29.885 ;
        RECT 141.725 29.175 142.055 29.345 ;
        RECT 141.725 27.625 142.055 27.795 ;
        RECT 142.425 27.455 142.650 41.685 ;
        RECT 143.015 40.165 143.345 40.335 ;
        RECT 143.015 39.625 143.345 39.795 ;
        RECT 143.015 38.075 143.345 38.245 ;
        RECT 143.015 37.535 143.345 37.705 ;
        RECT 143.015 35.985 143.345 36.155 ;
        RECT 143.015 35.445 143.345 35.615 ;
        RECT 143.015 33.895 143.345 34.065 ;
        RECT 143.015 33.355 143.345 33.525 ;
        RECT 143.015 31.805 143.345 31.975 ;
        RECT 143.015 31.265 143.345 31.435 ;
        RECT 143.015 29.715 143.345 29.885 ;
        RECT 143.015 29.175 143.345 29.345 ;
        RECT 143.015 27.625 143.345 27.795 ;
        RECT 143.715 27.455 143.940 41.685 ;
        RECT 144.305 40.165 144.635 40.335 ;
        RECT 144.305 39.625 144.635 39.795 ;
        RECT 144.305 38.075 144.635 38.245 ;
        RECT 144.305 37.535 144.635 37.705 ;
        RECT 144.305 35.985 144.635 36.155 ;
        RECT 144.305 35.445 144.635 35.615 ;
        RECT 144.305 33.895 144.635 34.065 ;
        RECT 144.305 33.355 144.635 33.525 ;
        RECT 144.305 31.805 144.635 31.975 ;
        RECT 144.305 31.265 144.635 31.435 ;
        RECT 144.305 29.715 144.635 29.885 ;
        RECT 144.305 29.175 144.635 29.345 ;
        RECT 144.305 27.625 144.635 27.795 ;
        RECT 145.000 27.455 145.225 41.685 ;
        RECT 145.595 40.165 145.925 40.335 ;
        RECT 145.595 39.625 145.925 39.795 ;
        RECT 145.595 38.075 145.925 38.245 ;
        RECT 145.595 37.535 145.925 37.705 ;
        RECT 145.595 35.985 145.925 36.155 ;
        RECT 145.595 35.445 145.925 35.615 ;
        RECT 145.595 33.895 145.925 34.065 ;
        RECT 145.595 33.355 145.925 33.525 ;
        RECT 145.595 31.805 145.925 31.975 ;
        RECT 145.595 31.265 145.925 31.435 ;
        RECT 145.595 29.715 145.925 29.885 ;
        RECT 145.595 29.175 145.925 29.345 ;
        RECT 145.595 27.625 145.925 27.795 ;
        RECT 146.285 27.455 146.510 41.685 ;
        RECT 146.885 40.165 147.215 40.335 ;
        RECT 146.885 39.625 147.215 39.795 ;
        RECT 146.885 38.075 147.215 38.245 ;
        RECT 146.885 37.535 147.215 37.705 ;
        RECT 146.885 35.985 147.215 36.155 ;
        RECT 146.885 35.445 147.215 35.615 ;
        RECT 146.885 33.895 147.215 34.065 ;
        RECT 146.885 33.355 147.215 33.525 ;
        RECT 146.885 31.805 147.215 31.975 ;
        RECT 146.885 31.265 147.215 31.435 ;
        RECT 146.885 29.715 147.215 29.885 ;
        RECT 146.885 29.175 147.215 29.345 ;
        RECT 146.885 27.625 147.215 27.795 ;
        RECT 147.580 27.455 147.805 41.685 ;
        RECT 148.175 40.165 148.505 40.335 ;
        RECT 148.175 39.625 148.505 39.795 ;
        RECT 148.175 38.075 148.505 38.245 ;
        RECT 148.175 37.535 148.505 37.705 ;
        RECT 148.175 35.985 148.505 36.155 ;
        RECT 148.175 35.445 148.505 35.615 ;
        RECT 148.175 33.895 148.505 34.065 ;
        RECT 148.175 33.355 148.505 33.525 ;
        RECT 148.175 31.805 148.505 31.975 ;
        RECT 148.175 31.265 148.505 31.435 ;
        RECT 148.175 29.715 148.505 29.885 ;
        RECT 148.175 29.175 148.505 29.345 ;
        RECT 148.175 27.625 148.505 27.795 ;
        RECT 148.870 27.780 149.095 41.870 ;
        RECT 156.830 34.555 163.450 41.935 ;
        RECT 156.530 34.385 163.450 34.555 ;
        RECT 142.830 26.820 143.140 26.840 ;
        RECT 148.800 26.820 149.230 27.780 ;
        RECT 156.830 27.005 163.450 34.385 ;
        RECT 156.530 26.835 163.450 27.005 ;
        RECT 115.750 25.090 116.080 26.490 ;
        RECT 122.170 26.430 122.470 26.490 ;
        RECT 128.910 26.220 135.890 26.660 ;
        RECT 142.780 26.290 149.230 26.820 ;
        RECT 142.780 26.260 149.220 26.290 ;
        RECT 116.280 25.770 116.860 25.940 ;
        RECT 118.040 25.570 119.070 25.790 ;
        RECT 117.060 25.170 119.070 25.570 ;
        RECT 116.280 24.800 116.860 24.970 ;
        RECT 118.040 24.930 119.070 25.170 ;
        RECT 128.910 24.930 129.220 26.220 ;
        RECT 129.390 25.550 129.970 25.720 ;
        RECT 131.130 25.340 132.160 25.560 ;
        RECT 130.120 24.940 132.160 25.340 ;
        RECT 142.830 25.120 143.140 26.260 ;
        RECT 143.390 25.680 143.970 25.850 ;
        RECT 145.000 25.490 146.030 25.700 ;
        RECT 142.950 25.115 143.120 25.120 ;
        RECT 144.140 25.040 146.030 25.490 ;
        RECT 129.390 24.580 129.970 24.750 ;
        RECT 131.130 24.700 132.160 24.940 ;
        RECT 143.390 24.710 143.970 24.880 ;
        RECT 145.000 24.840 146.030 25.040 ;
        RECT 156.830 19.455 163.450 26.835 ;
        RECT 97.800 19.280 104.715 19.450 ;
        RECT 156.530 19.285 163.450 19.455 ;
        RECT 97.800 19.200 104.445 19.280 ;
        RECT 156.830 19.205 163.450 19.285 ;
        RECT 165.915 110.055 172.570 110.280 ;
        RECT 165.915 109.885 172.820 110.055 ;
        RECT 165.915 109.455 172.570 109.885 ;
        RECT 165.915 102.505 172.550 109.455 ;
        RECT 234.280 107.470 236.440 107.820 ;
        RECT 255.690 107.470 257.850 107.820 ;
        RECT 281.670 107.480 283.830 107.830 ;
        RECT 234.280 105.880 236.440 106.230 ;
        RECT 255.690 105.880 257.850 106.230 ;
        RECT 281.670 105.890 283.830 106.240 ;
        RECT 255.690 104.290 257.850 104.640 ;
        RECT 260.260 104.300 262.420 104.650 ;
        RECT 281.670 104.300 283.830 104.650 ;
        RECT 255.690 102.700 257.850 103.050 ;
        RECT 260.260 102.710 262.420 103.060 ;
        RECT 281.670 102.710 283.830 103.060 ;
        RECT 165.915 102.335 172.820 102.505 ;
        RECT 165.915 94.955 172.550 102.335 ;
        RECT 255.690 101.110 257.850 101.460 ;
        RECT 260.260 101.120 262.420 101.470 ;
        RECT 281.670 101.120 283.830 101.470 ;
        RECT 234.280 99.520 236.440 99.870 ;
        RECT 255.690 99.520 257.850 99.870 ;
        RECT 281.670 99.530 283.830 99.880 ;
        RECT 234.280 97.930 236.440 98.280 ;
        RECT 260.260 97.940 262.420 98.290 ;
        RECT 234.280 96.340 236.440 96.690 ;
        RECT 260.260 96.350 262.420 96.700 ;
        RECT 165.915 94.785 172.820 94.955 ;
        RECT 165.915 87.405 172.550 94.785 ;
        RECT 255.690 94.750 257.850 95.100 ;
        RECT 260.260 94.760 262.420 95.110 ;
        RECT 386.260 90.880 386.630 93.050 ;
        RECT 387.850 90.880 388.220 93.050 ;
        RECT 244.060 89.360 244.760 89.520 ;
        RECT 236.610 89.330 244.760 89.360 ;
        RECT 225.000 89.150 244.760 89.330 ;
        RECT 225.000 89.140 236.880 89.150 ;
        RECT 165.915 87.235 172.820 87.405 ;
        RECT 225.040 87.290 225.230 89.140 ;
        RECT 236.770 88.950 236.990 88.960 ;
        RECT 230.110 88.760 236.990 88.950 ;
        RECT 244.060 88.900 244.760 89.150 ;
        RECT 230.110 87.290 230.300 88.760 ;
        RECT 165.915 79.855 172.550 87.235 ;
        RECT 224.190 86.920 226.240 87.290 ;
        RECT 227.070 86.660 227.690 87.120 ;
        RECT 229.230 86.920 231.280 87.290 ;
        RECT 227.230 86.500 227.570 86.660 ;
        RECT 223.150 86.280 225.290 86.290 ;
        RECT 223.150 85.960 225.300 86.280 ;
        RECT 210.980 83.060 213.210 83.120 ;
        RECT 210.980 82.940 215.530 83.060 ;
        RECT 165.915 79.685 172.820 79.855 ;
        RECT 165.915 72.305 172.550 79.685 ;
        RECT 210.980 75.010 211.210 82.940 ;
        RECT 213.030 82.890 215.530 82.940 ;
        RECT 213.030 82.715 213.310 82.890 ;
        RECT 212.950 82.690 213.310 82.715 ;
        RECT 215.260 82.800 215.530 82.890 ;
        RECT 212.950 82.545 213.280 82.690 ;
        RECT 214.110 82.535 214.440 82.705 ;
        RECT 215.260 82.695 215.580 82.800 ;
        RECT 215.250 82.525 215.580 82.695 ;
        RECT 216.340 82.535 216.670 82.705 ;
        RECT 215.310 82.510 215.520 82.525 ;
        RECT 212.810 80.370 212.980 82.250 ;
        RECT 213.250 80.370 213.420 82.250 ;
        RECT 213.970 80.360 214.140 82.240 ;
        RECT 214.410 80.360 214.580 82.240 ;
        RECT 215.110 80.350 215.280 82.230 ;
        RECT 215.550 80.350 215.720 82.230 ;
        RECT 216.200 80.360 216.370 82.240 ;
        RECT 216.640 80.360 216.810 82.240 ;
        RECT 212.990 80.075 213.230 80.090 ;
        RECT 212.950 79.905 213.280 80.075 ;
        RECT 213.670 80.065 214.390 80.100 ;
        RECT 214.780 80.090 215.090 80.100 ;
        RECT 212.990 79.750 213.230 79.905 ;
        RECT 213.670 79.900 214.440 80.065 ;
        RECT 212.090 79.510 213.440 79.520 ;
        RECT 213.670 79.510 213.850 79.900 ;
        RECT 214.110 79.895 214.440 79.900 ;
        RECT 214.780 80.055 215.530 80.090 ;
        RECT 215.910 80.065 216.600 80.080 ;
        RECT 212.080 79.310 213.850 79.510 ;
        RECT 214.780 79.885 215.580 80.055 ;
        RECT 215.910 79.895 216.670 80.065 ;
        RECT 215.910 79.890 216.600 79.895 ;
        RECT 214.780 79.840 215.530 79.885 ;
        RECT 214.780 79.770 215.090 79.840 ;
        RECT 214.780 79.490 214.970 79.770 ;
        RECT 215.910 79.490 216.090 79.890 ;
        RECT 214.150 79.320 214.970 79.490 ;
        RECT 215.240 79.320 216.090 79.490 ;
        RECT 216.350 79.310 216.680 79.480 ;
        RECT 212.080 79.290 213.440 79.310 ;
        RECT 212.080 75.550 212.290 79.290 ;
        RECT 212.930 78.180 213.100 79.060 ;
        RECT 213.370 78.180 213.540 79.060 ;
        RECT 214.010 78.190 214.180 79.070 ;
        RECT 214.450 78.190 214.620 79.070 ;
        RECT 215.100 78.190 215.270 79.070 ;
        RECT 215.540 78.190 215.710 79.070 ;
        RECT 216.210 78.180 216.380 79.060 ;
        RECT 216.650 78.180 216.820 79.060 ;
        RECT 223.160 78.910 223.370 85.960 ;
        RECT 225.080 85.900 225.300 85.960 ;
        RECT 225.090 85.790 225.300 85.900 ;
        RECT 227.240 85.900 227.570 86.500 ;
        RECT 223.820 83.310 223.990 85.540 ;
        RECT 225.090 85.340 225.310 85.790 ;
        RECT 223.770 82.360 224.030 83.310 ;
        RECT 225.110 82.940 225.280 85.340 ;
        RECT 226.400 83.290 226.570 85.540 ;
        RECT 226.360 82.420 226.620 83.290 ;
        RECT 227.240 82.420 227.550 85.900 ;
        RECT 230.080 85.780 232.270 86.280 ;
        RECT 228.820 83.130 228.990 85.540 ;
        RECT 230.090 85.350 230.310 85.780 ;
        RECT 225.430 82.360 227.550 82.420 ;
        RECT 223.770 82.320 227.550 82.360 ;
        RECT 228.790 82.470 229.020 83.130 ;
        RECT 230.110 82.940 230.280 85.350 ;
        RECT 231.400 83.190 231.570 85.540 ;
        RECT 231.370 82.470 231.600 83.190 ;
        RECT 228.790 82.320 231.600 82.470 ;
        RECT 223.770 82.000 231.600 82.320 ;
        RECT 223.770 81.990 226.630 82.000 ;
        RECT 227.160 81.990 231.600 82.000 ;
        RECT 225.010 81.980 225.380 81.990 ;
        RECT 226.360 81.980 226.620 81.990 ;
        RECT 228.790 81.980 231.600 81.990 ;
        RECT 228.810 81.940 231.600 81.980 ;
        RECT 232.080 80.590 232.270 85.780 ;
        RECT 231.950 80.410 232.280 80.590 ;
        RECT 223.160 78.720 227.410 78.910 ;
        RECT 225.780 78.030 226.750 78.350 ;
        RECT 227.190 78.030 227.390 78.720 ;
        RECT 213.150 77.930 213.330 77.950 ;
        RECT 214.420 77.940 214.870 77.980 ;
        RECT 213.070 77.760 213.400 77.930 ;
        RECT 214.150 77.770 214.870 77.940 ;
        RECT 215.240 77.770 215.570 77.950 ;
        RECT 215.910 77.930 216.350 77.980 ;
        RECT 213.150 77.580 213.330 77.760 ;
        RECT 214.420 77.750 214.870 77.770 ;
        RECT 215.330 77.580 215.500 77.770 ;
        RECT 215.910 77.760 216.680 77.930 ;
        RECT 225.780 77.790 227.420 78.030 ;
        RECT 215.910 77.750 216.350 77.760 ;
        RECT 215.910 77.720 216.190 77.750 ;
        RECT 213.150 77.380 215.500 77.580 ;
        RECT 225.780 77.470 226.750 77.790 ;
        RECT 212.020 75.200 212.400 75.550 ;
        RECT 210.760 74.420 211.370 75.010 ;
        RECT 227.190 74.300 227.390 77.790 ;
        RECT 230.850 76.640 231.820 76.950 ;
        RECT 232.060 76.640 232.280 80.410 ;
        RECT 236.770 77.250 236.990 88.760 ;
        RECT 245.530 88.550 245.910 89.250 ;
        RECT 246.410 88.590 246.840 89.250 ;
        RECT 250.050 88.590 250.550 89.340 ;
        RECT 258.930 88.620 259.520 89.510 ;
        RECT 238.920 84.380 239.410 84.690 ;
        RECT 243.120 84.680 243.590 84.770 ;
        RECT 244.890 84.680 245.360 84.770 ;
        RECT 243.120 84.460 245.360 84.680 ;
        RECT 238.970 83.190 239.280 84.380 ;
        RECT 243.120 84.370 243.590 84.460 ;
        RECT 244.890 84.370 245.360 84.460 ;
        RECT 238.080 83.180 239.280 83.190 ;
        RECT 237.690 83.150 239.280 83.180 ;
        RECT 237.680 83.010 241.460 83.150 ;
        RECT 236.710 76.910 237.020 77.250 ;
        RECT 236.770 76.900 236.990 76.910 ;
        RECT 230.850 76.400 232.310 76.640 ;
        RECT 230.850 76.070 231.820 76.400 ;
        RECT 227.180 74.060 227.400 74.300 ;
        RECT 232.060 74.210 232.280 76.400 ;
        RECT 237.680 75.800 237.890 83.010 ;
        RECT 238.960 82.980 241.460 83.010 ;
        RECT 238.960 82.805 239.240 82.980 ;
        RECT 238.880 82.780 239.240 82.805 ;
        RECT 241.190 82.890 241.460 82.980 ;
        RECT 238.880 82.635 239.210 82.780 ;
        RECT 240.040 82.625 240.370 82.795 ;
        RECT 241.190 82.785 241.510 82.890 ;
        RECT 241.180 82.615 241.510 82.785 ;
        RECT 242.270 82.625 242.600 82.795 ;
        RECT 241.240 82.600 241.450 82.615 ;
        RECT 238.740 80.460 238.910 82.340 ;
        RECT 239.180 80.460 239.350 82.340 ;
        RECT 239.900 80.450 240.070 82.330 ;
        RECT 240.340 80.450 240.510 82.330 ;
        RECT 241.040 80.440 241.210 82.320 ;
        RECT 241.480 80.440 241.650 82.320 ;
        RECT 242.130 80.450 242.300 82.330 ;
        RECT 242.570 80.450 242.740 82.330 ;
        RECT 238.920 80.165 239.160 80.180 ;
        RECT 238.880 79.995 239.210 80.165 ;
        RECT 239.600 80.155 240.320 80.190 ;
        RECT 240.710 80.180 241.020 80.190 ;
        RECT 238.920 79.840 239.160 79.995 ;
        RECT 239.600 79.990 240.370 80.155 ;
        RECT 239.600 79.610 239.780 79.990 ;
        RECT 240.040 79.985 240.370 79.990 ;
        RECT 240.710 80.145 241.460 80.180 ;
        RECT 241.840 80.155 242.530 80.170 ;
        RECT 238.130 79.400 239.780 79.610 ;
        RECT 240.710 79.975 241.510 80.145 ;
        RECT 241.840 79.985 242.600 80.155 ;
        RECT 241.840 79.980 242.530 79.985 ;
        RECT 240.710 79.930 241.460 79.975 ;
        RECT 240.710 79.860 241.020 79.930 ;
        RECT 240.710 79.580 240.900 79.860 ;
        RECT 241.840 79.580 242.020 79.980 ;
        RECT 240.080 79.410 240.900 79.580 ;
        RECT 241.170 79.410 242.020 79.580 ;
        RECT 242.280 79.400 242.610 79.570 ;
        RECT 238.130 79.380 239.640 79.400 ;
        RECT 237.680 74.600 237.880 75.800 ;
        RECT 238.150 75.560 238.350 79.380 ;
        RECT 238.860 78.270 239.030 79.150 ;
        RECT 239.300 78.270 239.470 79.150 ;
        RECT 239.940 78.280 240.110 79.160 ;
        RECT 240.380 78.280 240.550 79.160 ;
        RECT 241.030 78.280 241.200 79.160 ;
        RECT 241.470 78.280 241.640 79.160 ;
        RECT 242.140 78.270 242.310 79.150 ;
        RECT 242.580 78.270 242.750 79.150 ;
        RECT 239.080 78.020 239.260 78.040 ;
        RECT 240.350 78.030 240.800 78.070 ;
        RECT 239.000 77.850 239.330 78.020 ;
        RECT 240.080 77.860 240.800 78.030 ;
        RECT 241.170 77.860 241.500 78.040 ;
        RECT 241.840 78.020 242.280 78.070 ;
        RECT 239.080 77.670 239.260 77.850 ;
        RECT 240.350 77.840 240.800 77.860 ;
        RECT 241.260 77.670 241.430 77.860 ;
        RECT 241.840 77.850 242.610 78.020 ;
        RECT 241.840 77.840 242.280 77.850 ;
        RECT 241.840 77.810 242.120 77.840 ;
        RECT 239.080 77.470 241.430 77.670 ;
        RECT 240.870 76.420 241.210 77.470 ;
        RECT 240.820 75.970 241.310 76.420 ;
        RECT 238.050 75.230 238.470 75.560 ;
        RECT 237.610 74.380 237.950 74.600 ;
        RECT 165.915 72.135 172.820 72.305 ;
        RECT 165.915 64.755 172.550 72.135 ;
        RECT 227.190 71.300 227.390 74.060 ;
        RECT 232.050 73.910 232.290 74.210 ;
        RECT 232.060 71.300 232.280 73.910 ;
        RECT 227.190 70.870 227.430 71.300 ;
        RECT 232.060 71.110 232.300 71.300 ;
        RECT 227.210 70.720 227.430 70.870 ;
        RECT 224.140 69.980 226.220 70.150 ;
        RECT 227.230 68.940 227.420 70.720 ;
        RECT 232.090 70.700 232.300 71.110 ;
        RECT 229.000 69.980 231.080 70.150 ;
        RECT 232.100 68.970 232.290 70.700 ;
        RECT 165.915 64.585 172.820 64.755 ;
        RECT 165.915 57.205 172.550 64.585 ;
        RECT 245.620 64.090 245.840 88.550 ;
        RECT 246.500 65.270 246.710 88.590 ;
        RECT 250.160 86.380 250.500 88.590 ;
        RECT 253.670 86.760 254.330 87.180 ;
        RECT 256.950 87.060 257.730 87.610 ;
        RECT 250.160 81.620 250.460 86.380 ;
        RECT 253.860 85.910 254.130 86.760 ;
        RECT 256.090 85.920 256.440 85.930 ;
        RECT 257.180 85.920 257.470 87.060 ;
        RECT 259.080 86.510 259.420 88.620 ;
        RECT 271.260 87.560 271.800 88.140 ;
        RECT 278.420 87.640 278.910 88.020 ;
        RECT 280.780 87.640 281.100 87.690 ;
        RECT 288.710 87.640 289.680 87.740 ;
        RECT 250.660 85.635 251.240 85.805 ;
        RECT 253.105 85.765 255.480 85.910 ;
        RECT 253.055 85.595 255.480 85.765 ;
        RECT 253.105 85.550 255.480 85.595 ;
        RECT 256.090 85.570 258.880 85.920 ;
        RECT 256.395 85.560 258.880 85.570 ;
        RECT 250.220 81.600 250.390 81.620 ;
        RECT 251.430 80.040 251.710 84.220 ;
        RECT 253.925 84.160 254.095 84.440 ;
        RECT 257.215 84.170 257.385 84.300 ;
        RECT 252.550 81.590 252.840 84.160 ;
        RECT 253.905 82.610 254.095 84.160 ;
        RECT 255.195 84.150 255.365 84.160 ;
        RECT 253.905 82.020 254.075 82.610 ;
        RECT 252.615 81.560 252.785 81.590 ;
        RECT 253.890 79.910 254.120 82.020 ;
        RECT 255.175 80.410 255.385 84.150 ;
        RECT 255.895 81.620 256.095 84.170 ;
        RECT 257.195 82.940 257.385 84.170 ;
        RECT 257.165 82.170 257.395 82.940 ;
        RECT 255.905 81.570 256.075 81.620 ;
        RECT 253.680 79.470 254.350 79.910 ;
        RECT 255.150 79.010 255.390 80.410 ;
        RECT 257.180 79.850 257.380 82.170 ;
        RECT 258.485 81.940 258.655 84.170 ;
        RECT 258.450 81.570 258.655 81.940 ;
        RECT 258.450 80.210 258.645 81.570 ;
        RECT 259.110 81.510 259.370 86.510 ;
        RECT 259.630 85.505 260.210 85.675 ;
        RECT 260.480 84.060 260.650 84.070 ;
        RECT 259.190 81.470 259.360 81.510 ;
        RECT 258.450 80.200 258.660 80.210 ;
        RECT 255.100 78.460 255.390 79.010 ;
        RECT 255.100 77.110 255.360 78.460 ;
        RECT 250.010 76.910 255.360 77.110 ;
        RECT 250.030 76.820 255.360 76.910 ;
        RECT 257.160 77.120 257.400 79.850 ;
        RECT 258.440 78.750 258.670 80.200 ;
        RECT 260.430 79.700 260.690 84.060 ;
        RECT 262.110 82.990 262.990 83.740 ;
        RECT 264.370 83.640 264.880 84.070 ;
        RECT 264.480 83.210 264.670 83.640 ;
        RECT 264.480 83.040 267.340 83.210 ;
        RECT 262.350 81.570 262.550 82.990 ;
        RECT 264.840 82.865 265.120 83.040 ;
        RECT 264.760 82.840 265.120 82.865 ;
        RECT 267.070 82.950 267.340 83.040 ;
        RECT 264.760 82.695 265.090 82.840 ;
        RECT 265.920 82.685 266.250 82.855 ;
        RECT 267.070 82.845 267.390 82.950 ;
        RECT 267.060 82.675 267.390 82.845 ;
        RECT 268.150 82.685 268.480 82.855 ;
        RECT 267.120 82.660 267.330 82.675 ;
        RECT 262.350 81.370 264.390 81.570 ;
        RECT 258.440 78.610 258.660 78.750 ;
        RECT 260.420 78.440 260.690 79.700 ;
        RECT 263.340 79.560 263.920 80.070 ;
        RECT 260.010 77.830 261.020 78.440 ;
        RECT 257.160 76.930 258.680 77.120 ;
        RECT 250.030 76.690 250.320 76.820 ;
        RECT 257.160 76.780 260.990 76.930 ;
        RECT 257.160 76.770 257.400 76.780 ;
        RECT 250.010 76.620 250.320 76.690 ;
        RECT 258.440 76.660 260.990 76.780 ;
        RECT 250.010 76.035 250.360 76.620 ;
        RECT 260.100 76.500 260.990 76.660 ;
        RECT 253.210 76.040 253.600 76.080 ;
        RECT 258.280 76.040 258.670 76.080 ;
        RECT 249.915 75.345 250.480 76.035 ;
        RECT 253.210 76.030 253.640 76.040 ;
        RECT 255.680 76.030 255.860 76.040 ;
        RECT 258.280 76.030 258.710 76.040 ;
        RECT 251.870 75.900 255.900 76.030 ;
        RECT 256.940 75.970 260.700 76.030 ;
        RECT 261.000 75.970 261.880 76.050 ;
        RECT 256.940 75.900 261.880 75.970 ;
        RECT 251.850 75.730 255.900 75.900 ;
        RECT 256.920 75.730 261.880 75.900 ;
        RECT 251.870 75.700 255.900 75.730 ;
        RECT 256.940 75.700 261.880 75.730 ;
        RECT 250.060 70.020 250.330 75.345 ;
        RECT 251.315 73.640 251.575 75.100 ;
        RECT 251.350 72.190 251.570 73.640 ;
        RECT 251.870 73.120 252.300 75.700 ;
        RECT 252.660 74.990 252.830 74.995 ;
        RECT 252.580 74.030 252.880 74.990 ;
        RECT 253.210 73.120 253.640 75.700 ;
        RECT 251.850 72.950 252.350 73.120 ;
        RECT 253.140 72.950 253.640 73.120 ;
        RECT 251.870 72.880 252.300 72.950 ;
        RECT 253.210 72.930 253.640 72.950 ;
        RECT 251.330 71.290 251.570 72.190 ;
        RECT 252.600 71.300 252.900 72.260 ;
        RECT 253.920 72.010 254.140 75.040 ;
        RECT 254.500 73.120 254.930 75.700 ;
        RECT 255.210 74.110 255.510 75.070 ;
        RECT 255.240 74.085 255.410 74.110 ;
        RECT 254.430 72.950 254.930 73.120 ;
        RECT 254.500 72.920 254.930 72.950 ;
        RECT 253.900 71.340 254.140 72.010 ;
        RECT 251.330 70.850 251.550 71.290 ;
        RECT 253.900 70.850 254.120 71.340 ;
        RECT 255.220 71.330 255.500 72.290 ;
        RECT 255.240 71.305 255.410 71.330 ;
        RECT 251.320 70.460 254.140 70.850 ;
        RECT 250.060 69.700 250.390 70.020 ;
        RECT 253.290 69.070 253.490 70.460 ;
        RECT 255.680 70.120 255.860 75.700 ;
        RECT 256.385 73.640 256.645 75.100 ;
        RECT 256.420 72.190 256.640 73.640 ;
        RECT 256.940 73.120 257.370 75.700 ;
        RECT 257.730 74.990 257.900 74.995 ;
        RECT 257.650 74.030 257.950 74.990 ;
        RECT 258.280 73.120 258.710 75.700 ;
        RECT 256.920 72.950 257.420 73.120 ;
        RECT 258.210 72.950 258.710 73.120 ;
        RECT 256.940 72.880 257.370 72.950 ;
        RECT 258.280 72.930 258.710 72.950 ;
        RECT 256.400 71.290 256.640 72.190 ;
        RECT 257.670 71.300 257.970 72.260 ;
        RECT 258.990 72.010 259.210 75.040 ;
        RECT 259.570 73.120 260.000 75.700 ;
        RECT 261.000 75.610 261.880 75.700 ;
        RECT 260.280 74.110 260.580 75.070 ;
        RECT 260.310 74.085 260.480 74.110 ;
        RECT 259.500 72.950 260.000 73.120 ;
        RECT 259.570 72.920 260.000 72.950 ;
        RECT 258.970 71.340 259.210 72.010 ;
        RECT 256.400 70.850 256.620 71.290 ;
        RECT 258.970 70.850 259.190 71.340 ;
        RECT 260.290 71.330 260.570 72.290 ;
        RECT 260.310 71.305 260.480 71.330 ;
        RECT 256.390 70.520 259.210 70.850 ;
        RECT 256.390 70.460 259.660 70.520 ;
        RECT 258.360 70.340 259.660 70.460 ;
        RECT 255.520 69.440 256.120 70.120 ;
        RECT 259.440 69.680 259.660 70.340 ;
        RECT 259.440 69.670 261.560 69.680 ;
        RECT 262.200 69.670 262.800 69.840 ;
        RECT 259.440 69.460 262.800 69.670 ;
        RECT 261.300 69.450 262.800 69.460 ;
        RECT 262.200 69.380 262.800 69.450 ;
        RECT 263.410 69.070 263.590 79.560 ;
        RECT 253.290 68.880 263.590 69.070 ;
        RECT 264.100 73.810 264.270 81.370 ;
        RECT 264.620 80.520 264.790 82.400 ;
        RECT 265.060 80.520 265.230 82.400 ;
        RECT 265.780 80.510 265.950 82.390 ;
        RECT 266.220 80.510 266.390 82.390 ;
        RECT 266.920 80.500 267.090 82.380 ;
        RECT 267.360 80.500 267.530 82.380 ;
        RECT 268.010 80.510 268.180 82.390 ;
        RECT 268.450 80.510 268.620 82.390 ;
        RECT 264.800 80.225 265.040 80.240 ;
        RECT 264.760 80.055 265.090 80.225 ;
        RECT 265.480 80.215 266.200 80.250 ;
        RECT 266.590 80.240 266.900 80.250 ;
        RECT 264.800 79.900 265.040 80.055 ;
        RECT 265.480 80.050 266.250 80.215 ;
        RECT 265.480 79.660 265.660 80.050 ;
        RECT 265.920 80.045 266.250 80.050 ;
        RECT 266.590 80.205 267.340 80.240 ;
        RECT 267.720 80.215 268.410 80.230 ;
        RECT 264.520 79.460 265.660 79.660 ;
        RECT 266.590 80.035 267.390 80.205 ;
        RECT 267.720 80.045 268.480 80.215 ;
        RECT 267.720 80.040 268.410 80.045 ;
        RECT 266.590 79.990 267.340 80.035 ;
        RECT 266.590 79.920 266.900 79.990 ;
        RECT 266.590 79.640 266.780 79.920 ;
        RECT 267.720 79.640 267.900 80.040 ;
        RECT 265.960 79.470 266.780 79.640 ;
        RECT 267.050 79.470 267.900 79.640 ;
        RECT 268.160 79.460 268.490 79.630 ;
        RECT 264.520 79.430 265.230 79.460 ;
        RECT 264.740 78.330 264.910 79.210 ;
        RECT 265.180 78.330 265.350 79.210 ;
        RECT 265.820 78.340 265.990 79.220 ;
        RECT 266.260 78.340 266.430 79.220 ;
        RECT 266.910 78.340 267.080 79.220 ;
        RECT 267.350 78.340 267.520 79.220 ;
        RECT 268.020 78.330 268.190 79.210 ;
        RECT 268.460 78.330 268.630 79.210 ;
        RECT 264.960 78.080 265.140 78.100 ;
        RECT 266.230 78.090 266.680 78.130 ;
        RECT 264.880 77.910 265.210 78.080 ;
        RECT 265.960 77.920 266.680 78.090 ;
        RECT 267.050 77.920 267.380 78.100 ;
        RECT 267.720 78.080 268.160 78.130 ;
        RECT 264.960 77.730 265.140 77.910 ;
        RECT 266.230 77.900 266.680 77.920 ;
        RECT 267.140 77.730 267.310 77.920 ;
        RECT 267.720 77.910 268.490 78.080 ;
        RECT 267.720 77.900 268.160 77.910 ;
        RECT 267.720 77.870 268.000 77.900 ;
        RECT 264.960 77.530 267.310 77.730 ;
        RECT 265.800 77.090 266.020 77.530 ;
        RECT 265.750 77.010 266.190 77.090 ;
        RECT 270.910 77.010 271.150 77.090 ;
        RECT 265.750 76.760 271.150 77.010 ;
        RECT 265.750 76.670 266.190 76.760 ;
        RECT 270.910 76.700 271.150 76.760 ;
        RECT 270.870 73.810 271.170 74.000 ;
        RECT 264.100 73.580 271.170 73.810 ;
        RECT 264.100 68.570 264.270 73.580 ;
        RECT 270.870 73.480 271.170 73.580 ;
        RECT 265.830 72.610 266.150 72.830 ;
        RECT 255.210 68.330 264.270 68.570 ;
        RECT 265.800 68.720 266.150 72.610 ;
        RECT 265.800 68.500 266.140 68.720 ;
        RECT 255.210 67.050 255.490 68.330 ;
        RECT 268.980 68.030 269.700 68.260 ;
        RECT 261.250 67.990 269.700 68.030 ;
        RECT 258.230 67.760 269.700 67.990 ;
        RECT 258.230 67.050 258.500 67.760 ;
        RECT 261.250 67.750 269.700 67.760 ;
        RECT 268.980 67.600 269.700 67.750 ;
        RECT 253.615 67.005 255.040 67.015 ;
        RECT 253.160 66.695 255.040 67.005 ;
        RECT 253.615 66.665 255.040 66.695 ;
        RECT 255.210 66.600 255.480 67.050 ;
        RECT 256.645 66.910 257.750 67.015 ;
        RECT 256.645 66.900 257.755 66.910 ;
        RECT 256.640 66.730 257.755 66.900 ;
        RECT 256.645 66.720 257.755 66.730 ;
        RECT 256.645 66.665 257.750 66.720 ;
        RECT 252.975 66.325 253.145 66.340 ;
        RECT 252.915 66.285 253.145 66.325 ;
        RECT 252.915 65.690 253.165 66.285 ;
        RECT 255.250 65.785 255.475 66.600 ;
        RECT 255.865 66.290 256.125 66.355 ;
        RECT 258.255 66.340 258.455 67.050 ;
        RECT 255.265 65.740 255.435 65.785 ;
        RECT 252.970 65.270 253.165 65.690 ;
        RECT 255.865 65.735 256.180 66.290 ;
        RECT 258.240 65.810 258.455 66.340 ;
        RECT 258.240 65.740 258.410 65.810 ;
        RECT 255.865 65.270 256.125 65.735 ;
        RECT 246.500 65.040 253.180 65.270 ;
        RECT 252.970 65.020 253.165 65.040 ;
        RECT 255.870 64.090 256.120 65.270 ;
        RECT 245.620 63.890 256.120 64.090 ;
        RECT 271.440 57.350 271.650 87.560 ;
        RECT 278.520 84.040 278.770 87.640 ;
        RECT 280.750 87.470 289.680 87.640 ;
        RECT 279.330 85.075 280.250 85.090 ;
        RECT 279.250 84.905 280.330 85.075 ;
        RECT 279.330 84.900 280.250 84.905 ;
        RECT 278.520 83.190 278.760 84.040 ;
        RECT 280.780 83.200 281.100 87.470 ;
        RECT 288.710 87.420 289.680 87.470 ;
        RECT 289.160 87.130 289.830 87.140 ;
        RECT 283.890 87.110 289.830 87.130 ;
        RECT 283.630 86.930 289.830 87.110 ;
        RECT 281.350 86.040 281.650 86.550 ;
        RECT 281.370 83.880 281.620 86.040 ;
        RECT 282.190 85.075 283.110 85.100 ;
        RECT 282.110 84.905 283.190 85.075 ;
        RECT 281.380 83.200 281.620 83.880 ;
        RECT 283.630 83.250 283.950 86.930 ;
        RECT 289.160 86.890 289.830 86.930 ;
        RECT 278.560 80.870 278.730 83.190 ;
        RECT 280.850 81.240 281.020 83.200 ;
        RECT 280.690 79.130 281.120 81.240 ;
        RECT 281.420 80.870 281.590 83.200 ;
        RECT 283.710 81.140 283.880 83.250 ;
        RECT 295.140 82.880 295.820 83.420 ;
        RECT 291.420 82.170 293.310 82.200 ;
        RECT 295.340 82.170 295.630 82.880 ;
        RECT 291.420 82.020 295.630 82.170 ;
        RECT 283.560 79.180 284.070 81.140 ;
        RECT 280.690 79.090 281.000 79.130 ;
        RECT 280.560 77.410 281.000 79.090 ;
        RECT 283.560 79.070 283.980 79.180 ;
        RECT 280.530 76.840 281.030 77.410 ;
        RECT 283.550 77.360 283.980 79.070 ;
        RECT 287.330 77.620 287.770 77.930 ;
        RECT 283.510 76.910 284.100 77.360 ;
        RECT 280.560 73.900 281.000 76.840 ;
        RECT 280.580 73.890 281.000 73.900 ;
        RECT 283.550 74.070 283.980 76.910 ;
        RECT 287.410 76.690 287.670 77.620 ;
        RECT 291.420 77.170 291.660 82.020 ;
        RECT 293.120 82.000 295.630 82.020 ;
        RECT 293.120 81.825 293.400 82.000 ;
        RECT 293.040 81.800 293.400 81.825 ;
        RECT 295.350 81.830 295.620 82.000 ;
        RECT 293.040 81.655 293.370 81.800 ;
        RECT 294.200 81.645 294.530 81.815 ;
        RECT 295.350 81.805 295.670 81.830 ;
        RECT 295.340 81.635 295.670 81.805 ;
        RECT 296.430 81.645 296.760 81.815 ;
        RECT 295.400 81.620 295.610 81.635 ;
        RECT 292.900 79.480 293.070 81.360 ;
        RECT 293.340 79.480 293.510 81.360 ;
        RECT 294.060 79.470 294.230 81.350 ;
        RECT 294.500 79.470 294.670 81.350 ;
        RECT 295.200 79.460 295.370 81.340 ;
        RECT 295.640 79.460 295.810 81.340 ;
        RECT 296.290 79.470 296.460 81.350 ;
        RECT 296.730 79.470 296.900 81.350 ;
        RECT 482.180 81.300 489.520 82.190 ;
        RECT 482.110 80.710 489.520 81.300 ;
        RECT 481.900 80.570 489.520 80.710 ;
        RECT 536.610 80.570 543.320 82.690 ;
        RECT 293.080 79.185 293.320 79.200 ;
        RECT 293.040 79.015 293.370 79.185 ;
        RECT 293.760 79.175 294.480 79.210 ;
        RECT 294.870 79.200 295.180 79.210 ;
        RECT 293.080 78.860 293.320 79.015 ;
        RECT 293.760 79.010 294.530 79.175 ;
        RECT 293.760 78.620 293.940 79.010 ;
        RECT 294.200 79.005 294.530 79.010 ;
        RECT 294.870 79.165 295.620 79.200 ;
        RECT 296.000 79.175 296.690 79.190 ;
        RECT 292.320 78.420 293.940 78.620 ;
        RECT 294.870 78.995 295.670 79.165 ;
        RECT 296.000 79.005 296.760 79.175 ;
        RECT 296.000 79.000 296.690 79.005 ;
        RECT 294.870 78.950 295.620 78.995 ;
        RECT 294.870 78.880 295.180 78.950 ;
        RECT 294.870 78.600 295.060 78.880 ;
        RECT 296.000 78.600 296.180 79.000 ;
        RECT 294.240 78.430 295.060 78.600 ;
        RECT 295.330 78.430 296.180 78.600 ;
        RECT 296.440 78.420 296.770 78.590 ;
        RECT 481.900 78.210 543.320 80.570 ;
        RECT 293.020 77.290 293.190 78.170 ;
        RECT 293.460 77.290 293.630 78.170 ;
        RECT 294.100 77.300 294.270 78.180 ;
        RECT 294.540 77.300 294.710 78.180 ;
        RECT 295.190 77.300 295.360 78.180 ;
        RECT 295.630 77.300 295.800 78.180 ;
        RECT 296.300 77.290 296.470 78.170 ;
        RECT 296.740 77.290 296.910 78.170 ;
        RECT 291.420 76.830 291.750 77.170 ;
        RECT 293.240 77.040 293.420 77.060 ;
        RECT 294.510 77.050 294.960 77.090 ;
        RECT 293.160 76.870 293.490 77.040 ;
        RECT 294.240 76.880 294.960 77.050 ;
        RECT 295.330 76.880 295.660 77.060 ;
        RECT 296.000 77.040 296.440 77.090 ;
        RECT 291.420 76.810 291.660 76.830 ;
        RECT 293.240 76.690 293.420 76.870 ;
        RECT 294.510 76.860 294.960 76.880 ;
        RECT 295.420 76.690 295.590 76.880 ;
        RECT 296.000 76.870 296.770 77.040 ;
        RECT 296.000 76.860 296.440 76.870 ;
        RECT 296.000 76.830 296.280 76.860 ;
        RECT 481.900 76.810 489.520 78.210 ;
        RECT 536.610 77.580 543.320 78.210 ;
        RECT 287.410 76.650 291.240 76.690 ;
        RECT 291.950 76.660 295.590 76.690 ;
        RECT 304.770 76.660 305.230 76.720 ;
        RECT 482.180 76.710 489.520 76.810 ;
        RECT 287.410 76.630 291.250 76.650 ;
        RECT 291.950 76.630 305.250 76.660 ;
        RECT 287.410 76.490 305.250 76.630 ;
        RECT 287.410 76.480 293.940 76.490 ;
        RECT 295.200 76.480 305.250 76.490 ;
        RECT 291.160 76.430 292.140 76.480 ;
        RECT 304.770 76.450 305.230 76.480 ;
        RECT 291.240 76.420 291.980 76.430 ;
        RECT 277.220 72.210 277.800 72.380 ;
        RECT 278.510 72.210 279.090 72.380 ;
        RECT 279.800 72.210 280.380 72.380 ;
        RECT 280.580 72.010 281.010 73.890 ;
        RECT 283.550 73.880 283.960 74.070 ;
        RECT 283.550 73.640 285.880 73.880 ;
        RECT 285.600 73.120 285.880 73.640 ;
        RECT 282.220 72.210 282.800 72.380 ;
        RECT 283.510 72.210 284.090 72.380 ;
        RECT 284.800 72.210 285.380 72.380 ;
        RECT 278.020 71.660 281.010 72.010 ;
        RECT 285.650 71.990 285.870 73.120 ;
        RECT 283.010 71.980 283.400 71.990 ;
        RECT 284.020 71.980 285.880 71.990 ;
        RECT 276.730 59.620 277.010 71.120 ;
        RECT 277.220 67.430 277.800 67.600 ;
        RECT 277.220 62.650 277.800 62.820 ;
        RECT 276.710 59.460 277.010 59.620 ;
        RECT 276.710 58.980 277.000 59.460 ;
        RECT 278.020 59.300 278.300 71.660 ;
        RECT 279.360 70.980 279.530 71.070 ;
        RECT 278.510 67.430 279.090 67.600 ;
        RECT 278.510 62.650 279.090 62.820 ;
        RECT 279.320 59.650 279.600 70.980 ;
        RECT 280.600 70.960 280.880 71.660 ;
        RECT 283.010 71.640 285.880 71.980 ;
        RECT 281.780 71.020 281.950 71.070 ;
        RECT 283.040 71.040 283.290 71.640 ;
        RECT 285.610 71.610 285.870 71.640 ;
        RECT 284.360 71.060 284.530 71.070 ;
        RECT 280.600 70.710 280.890 70.960 ;
        RECT 279.800 67.430 280.380 67.600 ;
        RECT 279.800 62.650 280.380 62.820 ;
        RECT 279.320 58.980 279.610 59.650 ;
        RECT 280.610 59.300 280.890 70.710 ;
        RECT 281.720 59.600 282.000 71.020 ;
        RECT 282.220 67.430 282.800 67.600 ;
        RECT 282.220 62.650 282.800 62.820 ;
        RECT 281.720 59.360 282.020 59.600 ;
        RECT 283.030 59.380 283.310 71.040 ;
        RECT 283.510 67.430 284.090 67.600 ;
        RECT 283.510 62.650 284.090 62.820 ;
        RECT 284.290 59.600 284.570 71.060 ;
        RECT 285.610 71.040 285.860 71.610 ;
        RECT 284.800 67.430 285.380 67.600 ;
        RECT 284.800 62.650 285.380 62.820 ;
        RECT 284.290 59.400 284.600 59.600 ;
        RECT 281.730 58.980 282.020 59.360 ;
        RECT 284.310 58.980 284.600 59.400 ;
        RECT 285.580 59.380 285.860 71.040 ;
        RECT 276.690 58.440 284.600 58.980 ;
        RECT 281.080 57.350 281.280 58.440 ;
        RECT 165.915 57.035 172.820 57.205 ;
        RECT 271.440 57.130 281.280 57.350 ;
        RECT 271.440 57.120 281.270 57.130 ;
        RECT 165.915 49.655 172.550 57.035 ;
        RECT 501.290 56.630 572.910 59.720 ;
        RECT 197.560 55.905 197.890 56.075 ;
        RECT 189.090 55.015 193.170 55.185 ;
        RECT 195.110 54.260 195.420 54.740 ;
        RECT 197.860 54.360 198.030 55.300 ;
        RECT 190.110 51.450 190.440 51.620 ;
        RECT 197.480 51.400 197.810 51.570 ;
        RECT 197.780 50.835 197.950 51.165 ;
        RECT 197.480 50.430 197.810 50.600 ;
        RECT 165.915 49.485 172.820 49.655 ;
        RECT 165.915 42.105 172.550 49.485 ;
        RECT 190.360 45.950 190.700 49.660 ;
        RECT 190.110 43.900 190.440 44.070 ;
        RECT 165.915 41.935 172.820 42.105 ;
        RECT 165.915 34.555 172.550 41.935 ;
        RECT 271.970 40.160 274.130 40.510 ;
        RECT 250.560 38.480 252.720 38.830 ;
        RECT 271.970 38.480 274.130 38.830 ;
        RECT 250.750 36.810 252.910 37.160 ;
        RECT 272.160 36.810 274.320 37.160 ;
        RECT 272.260 35.220 274.420 35.570 ;
        RECT 165.915 34.385 172.820 34.555 ;
        RECT 165.915 27.005 172.550 34.385 ;
        RECT 293.110 29.165 294.950 29.170 ;
        RECT 293.030 28.995 295.030 29.165 ;
        RECT 293.110 28.990 294.950 28.995 ;
        RECT 165.915 26.835 172.820 27.005 ;
        RECT 165.915 19.455 172.550 26.835 ;
        RECT 270.670 25.725 274.670 25.895 ;
        RECT 275.660 25.885 279.510 25.890 ;
        RECT 270.750 25.720 274.590 25.725 ;
        RECT 275.590 25.715 279.590 25.885 ;
        RECT 249.890 25.245 269.730 25.250 ;
        RECT 249.810 25.075 269.810 25.245 ;
        RECT 249.890 25.070 269.730 25.075 ;
        RECT 269.870 24.780 270.040 24.860 ;
        RECT 269.870 23.900 270.050 24.780 ;
        RECT 269.870 23.820 270.040 23.900 ;
        RECT 274.730 23.810 274.900 25.510 ;
        RECT 279.650 25.420 279.820 25.500 ;
        RECT 279.650 23.870 279.830 25.420 ;
        RECT 281.040 23.910 281.210 28.950 ;
        RECT 282.330 23.910 282.500 28.950 ;
        RECT 292.800 28.710 292.970 28.780 ;
        RECT 288.610 28.300 288.780 28.370 ;
        RECT 288.610 26.690 288.790 28.300 ;
        RECT 288.610 26.610 288.780 26.690 ;
        RECT 284.620 26.395 288.480 26.400 ;
        RECT 284.550 26.225 288.550 26.395 ;
        RECT 284.620 26.220 288.480 26.225 ;
        RECT 284.160 25.525 292.000 25.540 ;
        RECT 284.080 25.355 292.080 25.525 ;
        RECT 284.160 25.350 292.000 25.355 ;
        RECT 292.140 24.560 292.310 25.140 ;
        RECT 279.650 23.800 279.820 23.870 ;
        RECT 292.800 23.820 292.980 28.710 ;
        RECT 292.800 23.740 292.970 23.820 ;
        RECT 295.090 23.740 295.260 28.780 ;
        RECT 281.350 23.695 282.190 23.700 ;
        RECT 281.270 23.525 282.270 23.695 ;
        RECT 249.610 23.120 257.450 23.130 ;
        RECT 249.530 22.950 257.530 23.120 ;
        RECT 257.590 21.460 257.760 22.780 ;
        RECT 266.440 21.750 266.610 23.070 ;
        RECT 274.730 21.750 274.900 23.070 ;
        RECT 283.020 21.750 283.190 23.070 ;
        RECT 294.030 23.010 295.030 23.180 ;
        RECT 290.900 22.920 291.740 22.930 ;
        RECT 289.530 22.750 290.530 22.920 ;
        RECT 290.820 22.750 291.820 22.920 ;
        RECT 284.310 22.410 288.310 22.580 ;
        RECT 290.590 22.500 290.760 22.580 ;
        RECT 258.380 21.410 266.380 21.580 ;
        RECT 266.670 21.410 274.670 21.580 ;
        RECT 274.960 21.410 282.960 21.580 ;
        RECT 288.370 21.200 288.540 22.240 ;
        RECT 258.460 20.620 266.460 20.790 ;
        RECT 266.750 20.620 274.750 20.790 ;
        RECT 275.040 20.620 283.040 20.790 ;
        RECT 249.580 19.920 257.580 20.090 ;
        RECT 249.660 19.910 257.500 19.920 ;
        RECT 165.915 19.285 172.820 19.455 ;
        RECT 165.915 19.205 172.550 19.285 ;
        RECT 249.350 18.430 249.520 19.750 ;
        RECT 257.640 18.430 257.810 19.750 ;
        RECT 123.750 15.655 124.080 15.825 ;
        RECT 140.660 15.565 140.990 15.735 ;
        RECT 159.130 15.655 159.460 15.825 ;
        RECT 266.520 15.580 266.690 20.450 ;
        RECT 274.810 15.580 274.980 20.450 ;
        RECT 283.100 15.580 283.270 20.450 ;
        RECT 290.580 19.620 290.760 22.500 ;
        RECT 295.090 21.780 295.260 22.840 ;
        RECT 294.030 21.440 295.030 21.610 ;
        RECT 290.590 19.540 290.760 19.620 ;
        RECT 289.530 19.200 290.530 19.370 ;
        RECT 290.820 19.200 291.820 19.370 ;
        RECT 115.280 14.765 119.360 14.935 ;
        RECT 132.190 14.675 136.270 14.845 ;
        RECT 121.290 14.010 121.600 14.490 ;
        RECT 138.240 13.930 138.550 14.410 ;
        RECT 140.960 14.020 141.130 14.960 ;
        RECT 150.660 14.765 154.740 14.935 ;
        RECT 156.720 14.020 157.030 14.500 ;
        RECT 159.430 14.110 159.600 15.050 ;
        RECT 258.550 14.520 266.390 14.530 ;
        RECT 275.120 14.520 282.960 14.530 ;
        RECT 258.460 14.350 266.460 14.520 ;
        RECT 266.750 14.350 274.750 14.520 ;
        RECT 275.040 14.350 283.040 14.520 ;
        RECT 258.550 14.330 266.390 14.350 ;
        RECT 266.810 14.340 274.680 14.350 ;
        RECT 266.520 12.640 266.690 14.180 ;
        RECT 274.810 12.640 274.980 14.180 ;
        RECT 283.100 12.640 283.270 14.180 ;
        RECT 116.300 11.200 116.630 11.370 ;
        RECT 123.670 11.150 124.000 11.320 ;
        RECT 133.210 11.110 133.540 11.280 ;
        RECT 140.580 11.060 140.910 11.230 ;
        RECT 151.680 11.200 152.010 11.370 ;
        RECT 159.050 11.150 159.380 11.320 ;
        RECT 140.880 10.495 141.050 10.825 ;
        RECT 159.350 10.585 159.520 10.915 ;
        RECT 123.670 10.180 124.000 10.350 ;
        RECT 140.580 10.090 140.910 10.260 ;
        RECT 159.050 10.180 159.380 10.350 ;
        RECT 116.550 5.700 116.890 9.410 ;
        RECT 133.460 5.610 133.800 9.320 ;
        RECT 151.930 5.700 152.270 9.410 ;
        RECT 116.300 3.650 116.630 3.820 ;
        RECT 133.210 3.560 133.540 3.730 ;
        RECT 151.680 3.650 152.010 3.820 ;
      LAYER mcon ;
        RECT 46.850 330.955 54.690 331.125 ;
        RECT 55.140 330.955 62.980 331.125 ;
        RECT 72.850 330.955 80.690 331.125 ;
        RECT 81.140 330.955 88.980 331.125 ;
        RECT 98.850 330.955 106.690 331.125 ;
        RECT 107.140 330.955 114.980 331.125 ;
        RECT 124.850 330.955 132.690 331.125 ;
        RECT 133.140 330.955 140.980 331.125 ;
        RECT 150.850 330.955 158.690 331.125 ;
        RECT 159.140 330.955 166.980 331.125 ;
        RECT 176.850 330.955 184.690 331.125 ;
        RECT 185.140 330.955 192.980 331.125 ;
        RECT 202.850 330.955 210.690 331.125 ;
        RECT 211.140 330.955 218.980 331.125 ;
        RECT 228.850 330.955 236.690 331.125 ;
        RECT 237.140 330.955 244.980 331.125 ;
        RECT 254.850 330.955 262.690 331.125 ;
        RECT 263.140 330.955 270.980 331.125 ;
        RECT 280.850 330.955 288.690 331.125 ;
        RECT 289.140 330.955 296.980 331.125 ;
        RECT 46.850 323.315 54.690 323.485 ;
        RECT 55.140 323.315 62.980 323.485 ;
        RECT 72.850 323.315 80.690 323.485 ;
        RECT 81.140 323.315 88.980 323.485 ;
        RECT 98.850 323.315 106.690 323.485 ;
        RECT 107.140 323.315 114.980 323.485 ;
        RECT 124.850 323.315 132.690 323.485 ;
        RECT 133.140 323.315 140.980 323.485 ;
        RECT 150.850 323.315 158.690 323.485 ;
        RECT 159.140 323.315 166.980 323.485 ;
        RECT 176.850 323.315 184.690 323.485 ;
        RECT 185.140 323.315 192.980 323.485 ;
        RECT 202.850 323.315 210.690 323.485 ;
        RECT 211.140 323.315 218.980 323.485 ;
        RECT 228.850 323.315 236.690 323.485 ;
        RECT 237.140 323.315 244.980 323.485 ;
        RECT 254.850 323.315 262.690 323.485 ;
        RECT 263.140 323.315 270.980 323.485 ;
        RECT 280.850 323.315 288.690 323.485 ;
        RECT 289.140 323.315 296.980 323.485 ;
        RECT 46.850 322.775 54.690 322.945 ;
        RECT 55.140 322.775 62.980 322.945 ;
        RECT 72.850 322.775 80.690 322.945 ;
        RECT 81.140 322.775 88.980 322.945 ;
        RECT 98.850 322.775 106.690 322.945 ;
        RECT 107.140 322.775 114.980 322.945 ;
        RECT 124.850 322.775 132.690 322.945 ;
        RECT 133.140 322.775 140.980 322.945 ;
        RECT 150.850 322.775 158.690 322.945 ;
        RECT 159.140 322.775 166.980 322.945 ;
        RECT 176.850 322.775 184.690 322.945 ;
        RECT 185.140 322.775 192.980 322.945 ;
        RECT 202.850 322.775 210.690 322.945 ;
        RECT 211.140 322.775 218.980 322.945 ;
        RECT 228.850 322.775 236.690 322.945 ;
        RECT 237.140 322.775 244.980 322.945 ;
        RECT 254.850 322.775 262.690 322.945 ;
        RECT 263.140 322.775 270.980 322.945 ;
        RECT 280.850 322.775 288.690 322.945 ;
        RECT 289.140 322.775 296.980 322.945 ;
        RECT 46.850 315.135 54.690 315.305 ;
        RECT 55.140 315.135 62.980 315.305 ;
        RECT 72.850 315.135 80.690 315.305 ;
        RECT 81.140 315.135 88.980 315.305 ;
        RECT 98.850 315.135 106.690 315.305 ;
        RECT 107.140 315.135 114.980 315.305 ;
        RECT 124.850 315.135 132.690 315.305 ;
        RECT 133.140 315.135 140.980 315.305 ;
        RECT 150.850 315.135 158.690 315.305 ;
        RECT 159.140 315.135 166.980 315.305 ;
        RECT 176.850 315.135 184.690 315.305 ;
        RECT 185.140 315.135 192.980 315.305 ;
        RECT 202.850 315.135 210.690 315.305 ;
        RECT 211.140 315.135 218.980 315.305 ;
        RECT 228.850 315.135 236.690 315.305 ;
        RECT 237.140 315.135 244.980 315.305 ;
        RECT 254.850 315.135 262.690 315.305 ;
        RECT 263.140 315.135 270.980 315.305 ;
        RECT 280.850 315.135 288.690 315.305 ;
        RECT 289.140 315.135 296.980 315.305 ;
        RECT 46.850 314.595 54.690 314.765 ;
        RECT 55.140 314.595 62.980 314.765 ;
        RECT 72.850 314.595 80.690 314.765 ;
        RECT 81.140 314.595 88.980 314.765 ;
        RECT 98.850 314.595 106.690 314.765 ;
        RECT 107.140 314.595 114.980 314.765 ;
        RECT 124.850 314.595 132.690 314.765 ;
        RECT 133.140 314.595 140.980 314.765 ;
        RECT 150.850 314.595 158.690 314.765 ;
        RECT 159.140 314.595 166.980 314.765 ;
        RECT 176.850 314.595 184.690 314.765 ;
        RECT 185.140 314.595 192.980 314.765 ;
        RECT 202.850 314.595 210.690 314.765 ;
        RECT 211.140 314.595 218.980 314.765 ;
        RECT 228.850 314.595 236.690 314.765 ;
        RECT 237.140 314.595 244.980 314.765 ;
        RECT 254.850 314.595 262.690 314.765 ;
        RECT 263.140 314.595 270.980 314.765 ;
        RECT 280.850 314.595 288.690 314.765 ;
        RECT 289.140 314.595 296.980 314.765 ;
        RECT 46.850 306.955 54.690 307.125 ;
        RECT 55.140 306.955 62.980 307.125 ;
        RECT 72.850 306.955 80.690 307.125 ;
        RECT 81.140 306.955 88.980 307.125 ;
        RECT 98.850 306.955 106.690 307.125 ;
        RECT 107.140 306.955 114.980 307.125 ;
        RECT 124.850 306.955 132.690 307.125 ;
        RECT 133.140 306.955 140.980 307.125 ;
        RECT 150.850 306.955 158.690 307.125 ;
        RECT 159.140 306.955 166.980 307.125 ;
        RECT 176.850 306.955 184.690 307.125 ;
        RECT 185.140 306.955 192.980 307.125 ;
        RECT 202.850 306.955 210.690 307.125 ;
        RECT 211.140 306.955 218.980 307.125 ;
        RECT 228.850 306.955 236.690 307.125 ;
        RECT 237.140 306.955 244.980 307.125 ;
        RECT 254.850 306.955 262.690 307.125 ;
        RECT 263.140 306.955 270.980 307.125 ;
        RECT 280.850 306.955 288.690 307.125 ;
        RECT 289.140 306.955 296.980 307.125 ;
        RECT 46.850 306.415 54.690 306.585 ;
        RECT 55.140 306.415 62.980 306.585 ;
        RECT 72.850 306.415 80.690 306.585 ;
        RECT 81.140 306.415 88.980 306.585 ;
        RECT 98.850 306.415 106.690 306.585 ;
        RECT 107.140 306.415 114.980 306.585 ;
        RECT 124.850 306.415 132.690 306.585 ;
        RECT 133.140 306.415 140.980 306.585 ;
        RECT 150.850 306.415 158.690 306.585 ;
        RECT 159.140 306.415 166.980 306.585 ;
        RECT 176.850 306.415 184.690 306.585 ;
        RECT 185.140 306.415 192.980 306.585 ;
        RECT 202.850 306.415 210.690 306.585 ;
        RECT 211.140 306.415 218.980 306.585 ;
        RECT 228.850 306.415 236.690 306.585 ;
        RECT 237.140 306.415 244.980 306.585 ;
        RECT 254.850 306.415 262.690 306.585 ;
        RECT 263.140 306.415 270.980 306.585 ;
        RECT 280.850 306.415 288.690 306.585 ;
        RECT 289.140 306.415 296.980 306.585 ;
        RECT 46.850 298.775 54.690 298.945 ;
        RECT 55.140 298.775 62.980 298.945 ;
        RECT 72.850 298.775 80.690 298.945 ;
        RECT 81.140 298.775 88.980 298.945 ;
        RECT 98.850 298.775 106.690 298.945 ;
        RECT 107.140 298.775 114.980 298.945 ;
        RECT 124.850 298.775 132.690 298.945 ;
        RECT 133.140 298.775 140.980 298.945 ;
        RECT 150.850 298.775 158.690 298.945 ;
        RECT 159.140 298.775 166.980 298.945 ;
        RECT 176.850 298.775 184.690 298.945 ;
        RECT 185.140 298.775 192.980 298.945 ;
        RECT 202.850 298.775 210.690 298.945 ;
        RECT 211.140 298.775 218.980 298.945 ;
        RECT 228.850 298.775 236.690 298.945 ;
        RECT 237.140 298.775 244.980 298.945 ;
        RECT 254.850 298.775 262.690 298.945 ;
        RECT 263.140 298.775 270.980 298.945 ;
        RECT 280.850 298.775 288.690 298.945 ;
        RECT 289.140 298.775 296.980 298.945 ;
        RECT 46.850 298.235 54.690 298.405 ;
        RECT 55.140 298.235 62.980 298.405 ;
        RECT 72.850 298.235 80.690 298.405 ;
        RECT 81.140 298.235 88.980 298.405 ;
        RECT 98.850 298.235 106.690 298.405 ;
        RECT 107.140 298.235 114.980 298.405 ;
        RECT 124.850 298.235 132.690 298.405 ;
        RECT 133.140 298.235 140.980 298.405 ;
        RECT 150.850 298.235 158.690 298.405 ;
        RECT 159.140 298.235 166.980 298.405 ;
        RECT 176.850 298.235 184.690 298.405 ;
        RECT 185.140 298.235 192.980 298.405 ;
        RECT 202.850 298.235 210.690 298.405 ;
        RECT 211.140 298.235 218.980 298.405 ;
        RECT 228.850 298.235 236.690 298.405 ;
        RECT 237.140 298.235 244.980 298.405 ;
        RECT 254.850 298.235 262.690 298.405 ;
        RECT 263.140 298.235 270.980 298.405 ;
        RECT 280.850 298.235 288.690 298.405 ;
        RECT 289.140 298.235 296.980 298.405 ;
        RECT 46.850 290.595 54.690 290.765 ;
        RECT 55.140 290.595 62.980 290.765 ;
        RECT 72.850 290.595 80.690 290.765 ;
        RECT 81.140 290.595 88.980 290.765 ;
        RECT 98.850 290.595 106.690 290.765 ;
        RECT 107.140 290.595 114.980 290.765 ;
        RECT 124.850 290.595 132.690 290.765 ;
        RECT 133.140 290.595 140.980 290.765 ;
        RECT 150.850 290.595 158.690 290.765 ;
        RECT 159.140 290.595 166.980 290.765 ;
        RECT 176.850 290.595 184.690 290.765 ;
        RECT 185.140 290.595 192.980 290.765 ;
        RECT 202.850 290.595 210.690 290.765 ;
        RECT 211.140 290.595 218.980 290.765 ;
        RECT 228.850 290.595 236.690 290.765 ;
        RECT 237.140 290.595 244.980 290.765 ;
        RECT 254.850 290.595 262.690 290.765 ;
        RECT 263.140 290.595 270.980 290.765 ;
        RECT 280.850 290.595 288.690 290.765 ;
        RECT 289.140 290.595 296.980 290.765 ;
        RECT 46.850 290.055 54.690 290.225 ;
        RECT 55.140 290.055 62.980 290.225 ;
        RECT 72.850 290.055 80.690 290.225 ;
        RECT 81.140 290.055 88.980 290.225 ;
        RECT 98.850 290.055 106.690 290.225 ;
        RECT 107.140 290.055 114.980 290.225 ;
        RECT 124.850 290.055 132.690 290.225 ;
        RECT 133.140 290.055 140.980 290.225 ;
        RECT 150.850 290.055 158.690 290.225 ;
        RECT 159.140 290.055 166.980 290.225 ;
        RECT 176.850 290.055 184.690 290.225 ;
        RECT 185.140 290.055 192.980 290.225 ;
        RECT 202.850 290.055 210.690 290.225 ;
        RECT 211.140 290.055 218.980 290.225 ;
        RECT 228.850 290.055 236.690 290.225 ;
        RECT 237.140 290.055 244.980 290.225 ;
        RECT 254.850 290.055 262.690 290.225 ;
        RECT 263.140 290.055 270.980 290.225 ;
        RECT 280.850 290.055 288.690 290.225 ;
        RECT 289.140 290.055 296.980 290.225 ;
        RECT 46.850 282.415 54.690 282.585 ;
        RECT 55.140 282.415 62.980 282.585 ;
        RECT 72.850 282.415 80.690 282.585 ;
        RECT 81.140 282.415 88.980 282.585 ;
        RECT 98.850 282.415 106.690 282.585 ;
        RECT 107.140 282.415 114.980 282.585 ;
        RECT 124.850 282.415 132.690 282.585 ;
        RECT 133.140 282.415 140.980 282.585 ;
        RECT 150.850 282.415 158.690 282.585 ;
        RECT 159.140 282.415 166.980 282.585 ;
        RECT 176.850 282.415 184.690 282.585 ;
        RECT 185.140 282.415 192.980 282.585 ;
        RECT 202.850 282.415 210.690 282.585 ;
        RECT 211.140 282.415 218.980 282.585 ;
        RECT 228.850 282.415 236.690 282.585 ;
        RECT 237.140 282.415 244.980 282.585 ;
        RECT 254.850 282.415 262.690 282.585 ;
        RECT 263.140 282.415 270.980 282.585 ;
        RECT 280.850 282.415 288.690 282.585 ;
        RECT 289.140 282.415 296.980 282.585 ;
        RECT 46.850 281.875 54.690 282.045 ;
        RECT 55.140 281.875 62.980 282.045 ;
        RECT 72.850 281.875 80.690 282.045 ;
        RECT 81.140 281.875 88.980 282.045 ;
        RECT 98.850 281.875 106.690 282.045 ;
        RECT 107.140 281.875 114.980 282.045 ;
        RECT 124.850 281.875 132.690 282.045 ;
        RECT 133.140 281.875 140.980 282.045 ;
        RECT 150.850 281.875 158.690 282.045 ;
        RECT 159.140 281.875 166.980 282.045 ;
        RECT 176.850 281.875 184.690 282.045 ;
        RECT 185.140 281.875 192.980 282.045 ;
        RECT 202.850 281.875 210.690 282.045 ;
        RECT 211.140 281.875 218.980 282.045 ;
        RECT 228.850 281.875 236.690 282.045 ;
        RECT 237.140 281.875 244.980 282.045 ;
        RECT 254.850 281.875 262.690 282.045 ;
        RECT 263.140 281.875 270.980 282.045 ;
        RECT 280.850 281.875 288.690 282.045 ;
        RECT 289.140 281.875 296.980 282.045 ;
        RECT 46.850 274.235 54.690 274.405 ;
        RECT 55.140 274.235 62.980 274.405 ;
        RECT 72.850 274.235 80.690 274.405 ;
        RECT 81.140 274.235 88.980 274.405 ;
        RECT 98.850 274.235 106.690 274.405 ;
        RECT 107.140 274.235 114.980 274.405 ;
        RECT 124.850 274.235 132.690 274.405 ;
        RECT 133.140 274.235 140.980 274.405 ;
        RECT 150.850 274.235 158.690 274.405 ;
        RECT 159.140 274.235 166.980 274.405 ;
        RECT 176.850 274.235 184.690 274.405 ;
        RECT 185.140 274.235 192.980 274.405 ;
        RECT 202.850 274.235 210.690 274.405 ;
        RECT 211.140 274.235 218.980 274.405 ;
        RECT 228.850 274.235 236.690 274.405 ;
        RECT 237.140 274.235 244.980 274.405 ;
        RECT 254.850 274.235 262.690 274.405 ;
        RECT 263.140 274.235 270.980 274.405 ;
        RECT 280.850 274.235 288.690 274.405 ;
        RECT 289.140 274.235 296.980 274.405 ;
        RECT 46.850 273.695 54.690 273.865 ;
        RECT 55.140 273.695 62.980 273.865 ;
        RECT 72.850 273.695 80.690 273.865 ;
        RECT 81.140 273.695 88.980 273.865 ;
        RECT 98.850 273.695 106.690 273.865 ;
        RECT 107.140 273.695 114.980 273.865 ;
        RECT 124.850 273.695 132.690 273.865 ;
        RECT 133.140 273.695 140.980 273.865 ;
        RECT 150.850 273.695 158.690 273.865 ;
        RECT 159.140 273.695 166.980 273.865 ;
        RECT 176.850 273.695 184.690 273.865 ;
        RECT 185.140 273.695 192.980 273.865 ;
        RECT 202.850 273.695 210.690 273.865 ;
        RECT 211.140 273.695 218.980 273.865 ;
        RECT 228.850 273.695 236.690 273.865 ;
        RECT 237.140 273.695 244.980 273.865 ;
        RECT 254.850 273.695 262.690 273.865 ;
        RECT 263.140 273.695 270.980 273.865 ;
        RECT 280.850 273.695 288.690 273.865 ;
        RECT 289.140 273.695 296.980 273.865 ;
        RECT 46.850 266.055 54.690 266.225 ;
        RECT 55.140 266.055 62.980 266.225 ;
        RECT 72.850 266.055 80.690 266.225 ;
        RECT 81.140 266.055 88.980 266.225 ;
        RECT 98.850 266.055 106.690 266.225 ;
        RECT 107.140 266.055 114.980 266.225 ;
        RECT 124.850 266.055 132.690 266.225 ;
        RECT 133.140 266.055 140.980 266.225 ;
        RECT 150.850 266.055 158.690 266.225 ;
        RECT 159.140 266.055 166.980 266.225 ;
        RECT 176.850 266.055 184.690 266.225 ;
        RECT 185.140 266.055 192.980 266.225 ;
        RECT 202.850 266.055 210.690 266.225 ;
        RECT 211.140 266.055 218.980 266.225 ;
        RECT 228.850 266.055 236.690 266.225 ;
        RECT 237.140 266.055 244.980 266.225 ;
        RECT 254.850 266.055 262.690 266.225 ;
        RECT 263.140 266.055 270.980 266.225 ;
        RECT 280.850 266.055 288.690 266.225 ;
        RECT 289.140 266.055 296.980 266.225 ;
        RECT 46.850 265.515 54.690 265.685 ;
        RECT 55.140 265.515 62.980 265.685 ;
        RECT 72.850 265.515 80.690 265.685 ;
        RECT 81.140 265.515 88.980 265.685 ;
        RECT 98.850 265.515 106.690 265.685 ;
        RECT 107.140 265.515 114.980 265.685 ;
        RECT 124.850 265.515 132.690 265.685 ;
        RECT 133.140 265.515 140.980 265.685 ;
        RECT 150.850 265.515 158.690 265.685 ;
        RECT 159.140 265.515 166.980 265.685 ;
        RECT 176.850 265.515 184.690 265.685 ;
        RECT 185.140 265.515 192.980 265.685 ;
        RECT 202.850 265.515 210.690 265.685 ;
        RECT 211.140 265.515 218.980 265.685 ;
        RECT 228.850 265.515 236.690 265.685 ;
        RECT 237.140 265.515 244.980 265.685 ;
        RECT 254.850 265.515 262.690 265.685 ;
        RECT 263.140 265.515 270.980 265.685 ;
        RECT 280.850 265.515 288.690 265.685 ;
        RECT 289.140 265.515 296.980 265.685 ;
        RECT 46.850 257.875 54.690 258.045 ;
        RECT 55.140 257.875 62.980 258.045 ;
        RECT 72.850 257.875 80.690 258.045 ;
        RECT 81.140 257.875 88.980 258.045 ;
        RECT 98.850 257.875 106.690 258.045 ;
        RECT 107.140 257.875 114.980 258.045 ;
        RECT 124.850 257.875 132.690 258.045 ;
        RECT 133.140 257.875 140.980 258.045 ;
        RECT 150.850 257.875 158.690 258.045 ;
        RECT 159.140 257.875 166.980 258.045 ;
        RECT 176.850 257.875 184.690 258.045 ;
        RECT 185.140 257.875 192.980 258.045 ;
        RECT 202.850 257.875 210.690 258.045 ;
        RECT 211.140 257.875 218.980 258.045 ;
        RECT 228.850 257.875 236.690 258.045 ;
        RECT 237.140 257.875 244.980 258.045 ;
        RECT 254.850 257.875 262.690 258.045 ;
        RECT 263.140 257.875 270.980 258.045 ;
        RECT 280.850 257.875 288.690 258.045 ;
        RECT 289.140 257.875 296.980 258.045 ;
        RECT 46.850 257.335 54.690 257.505 ;
        RECT 55.140 257.335 62.980 257.505 ;
        RECT 72.850 257.335 80.690 257.505 ;
        RECT 81.140 257.335 88.980 257.505 ;
        RECT 98.850 257.335 106.690 257.505 ;
        RECT 107.140 257.335 114.980 257.505 ;
        RECT 124.850 257.335 132.690 257.505 ;
        RECT 133.140 257.335 140.980 257.505 ;
        RECT 150.850 257.335 158.690 257.505 ;
        RECT 159.140 257.335 166.980 257.505 ;
        RECT 176.850 257.335 184.690 257.505 ;
        RECT 185.140 257.335 192.980 257.505 ;
        RECT 202.850 257.335 210.690 257.505 ;
        RECT 211.140 257.335 218.980 257.505 ;
        RECT 228.850 257.335 236.690 257.505 ;
        RECT 237.140 257.335 244.980 257.505 ;
        RECT 254.850 257.335 262.690 257.505 ;
        RECT 263.140 257.335 270.980 257.505 ;
        RECT 280.850 257.335 288.690 257.505 ;
        RECT 289.140 257.335 296.980 257.505 ;
        RECT 46.850 249.695 54.690 249.865 ;
        RECT 55.140 249.695 62.980 249.865 ;
        RECT 72.850 249.695 80.690 249.865 ;
        RECT 81.140 249.695 88.980 249.865 ;
        RECT 98.850 249.695 106.690 249.865 ;
        RECT 107.140 249.695 114.980 249.865 ;
        RECT 124.850 249.695 132.690 249.865 ;
        RECT 133.140 249.695 140.980 249.865 ;
        RECT 150.850 249.695 158.690 249.865 ;
        RECT 159.140 249.695 166.980 249.865 ;
        RECT 176.850 249.695 184.690 249.865 ;
        RECT 185.140 249.695 192.980 249.865 ;
        RECT 202.850 249.695 210.690 249.865 ;
        RECT 211.140 249.695 218.980 249.865 ;
        RECT 228.850 249.695 236.690 249.865 ;
        RECT 237.140 249.695 244.980 249.865 ;
        RECT 254.850 249.695 262.690 249.865 ;
        RECT 263.140 249.695 270.980 249.865 ;
        RECT 280.850 249.695 288.690 249.865 ;
        RECT 289.140 249.695 296.980 249.865 ;
        RECT 46.850 249.155 54.690 249.325 ;
        RECT 55.140 249.155 62.980 249.325 ;
        RECT 72.850 249.155 80.690 249.325 ;
        RECT 81.140 249.155 88.980 249.325 ;
        RECT 98.850 249.155 106.690 249.325 ;
        RECT 107.140 249.155 114.980 249.325 ;
        RECT 124.850 249.155 132.690 249.325 ;
        RECT 133.140 249.155 140.980 249.325 ;
        RECT 150.850 249.155 158.690 249.325 ;
        RECT 159.140 249.155 166.980 249.325 ;
        RECT 176.850 249.155 184.690 249.325 ;
        RECT 185.140 249.155 192.980 249.325 ;
        RECT 202.850 249.155 210.690 249.325 ;
        RECT 211.140 249.155 218.980 249.325 ;
        RECT 228.850 249.155 236.690 249.325 ;
        RECT 237.140 249.155 244.980 249.325 ;
        RECT 254.850 249.155 262.690 249.325 ;
        RECT 263.140 249.155 270.980 249.325 ;
        RECT 280.850 249.155 288.690 249.325 ;
        RECT 289.140 249.155 296.980 249.325 ;
        RECT 46.850 241.515 54.690 241.685 ;
        RECT 55.140 241.515 62.980 241.685 ;
        RECT 72.850 241.515 80.690 241.685 ;
        RECT 81.140 241.515 88.980 241.685 ;
        RECT 98.850 241.515 106.690 241.685 ;
        RECT 107.140 241.515 114.980 241.685 ;
        RECT 124.850 241.515 132.690 241.685 ;
        RECT 133.140 241.515 140.980 241.685 ;
        RECT 150.850 241.515 158.690 241.685 ;
        RECT 159.140 241.515 166.980 241.685 ;
        RECT 176.850 241.515 184.690 241.685 ;
        RECT 185.140 241.515 192.980 241.685 ;
        RECT 202.850 241.515 210.690 241.685 ;
        RECT 211.140 241.515 218.980 241.685 ;
        RECT 228.850 241.515 236.690 241.685 ;
        RECT 237.140 241.515 244.980 241.685 ;
        RECT 254.850 241.515 262.690 241.685 ;
        RECT 263.140 241.515 270.980 241.685 ;
        RECT 280.850 241.515 288.690 241.685 ;
        RECT 289.140 241.515 296.980 241.685 ;
        RECT 46.850 240.975 54.690 241.145 ;
        RECT 55.140 240.975 62.980 241.145 ;
        RECT 72.850 240.975 80.690 241.145 ;
        RECT 81.140 240.975 88.980 241.145 ;
        RECT 98.850 240.975 106.690 241.145 ;
        RECT 107.140 240.975 114.980 241.145 ;
        RECT 124.850 240.975 132.690 241.145 ;
        RECT 133.140 240.975 140.980 241.145 ;
        RECT 150.850 240.975 158.690 241.145 ;
        RECT 159.140 240.975 166.980 241.145 ;
        RECT 176.850 240.975 184.690 241.145 ;
        RECT 185.140 240.975 192.980 241.145 ;
        RECT 202.850 240.975 210.690 241.145 ;
        RECT 211.140 240.975 218.980 241.145 ;
        RECT 228.850 240.975 236.690 241.145 ;
        RECT 237.140 240.975 244.980 241.145 ;
        RECT 254.850 240.975 262.690 241.145 ;
        RECT 263.140 240.975 270.980 241.145 ;
        RECT 280.850 240.975 288.690 241.145 ;
        RECT 289.140 240.975 296.980 241.145 ;
        RECT 46.850 233.335 54.690 233.505 ;
        RECT 55.140 233.335 62.980 233.505 ;
        RECT 72.850 233.335 80.690 233.505 ;
        RECT 81.140 233.335 88.980 233.505 ;
        RECT 98.850 233.335 106.690 233.505 ;
        RECT 107.140 233.335 114.980 233.505 ;
        RECT 124.850 233.335 132.690 233.505 ;
        RECT 133.140 233.335 140.980 233.505 ;
        RECT 150.850 233.335 158.690 233.505 ;
        RECT 159.140 233.335 166.980 233.505 ;
        RECT 176.850 233.335 184.690 233.505 ;
        RECT 185.140 233.335 192.980 233.505 ;
        RECT 202.850 233.335 210.690 233.505 ;
        RECT 211.140 233.335 218.980 233.505 ;
        RECT 228.850 233.335 236.690 233.505 ;
        RECT 237.140 233.335 244.980 233.505 ;
        RECT 254.850 233.335 262.690 233.505 ;
        RECT 263.140 233.335 270.980 233.505 ;
        RECT 280.850 233.335 288.690 233.505 ;
        RECT 289.140 233.335 296.980 233.505 ;
        RECT 46.850 232.795 54.690 232.965 ;
        RECT 55.140 232.795 62.980 232.965 ;
        RECT 72.850 232.795 80.690 232.965 ;
        RECT 81.140 232.795 88.980 232.965 ;
        RECT 98.850 232.795 106.690 232.965 ;
        RECT 107.140 232.795 114.980 232.965 ;
        RECT 124.850 232.795 132.690 232.965 ;
        RECT 133.140 232.795 140.980 232.965 ;
        RECT 150.850 232.795 158.690 232.965 ;
        RECT 159.140 232.795 166.980 232.965 ;
        RECT 176.850 232.795 184.690 232.965 ;
        RECT 185.140 232.795 192.980 232.965 ;
        RECT 202.850 232.795 210.690 232.965 ;
        RECT 211.140 232.795 218.980 232.965 ;
        RECT 228.850 232.795 236.690 232.965 ;
        RECT 237.140 232.795 244.980 232.965 ;
        RECT 254.850 232.795 262.690 232.965 ;
        RECT 263.140 232.795 270.980 232.965 ;
        RECT 280.850 232.795 288.690 232.965 ;
        RECT 289.140 232.795 296.980 232.965 ;
        RECT 46.850 225.155 54.690 225.325 ;
        RECT 55.140 225.155 62.980 225.325 ;
        RECT 72.850 225.155 80.690 225.325 ;
        RECT 81.140 225.155 88.980 225.325 ;
        RECT 98.850 225.155 106.690 225.325 ;
        RECT 107.140 225.155 114.980 225.325 ;
        RECT 124.850 225.155 132.690 225.325 ;
        RECT 133.140 225.155 140.980 225.325 ;
        RECT 150.850 225.155 158.690 225.325 ;
        RECT 159.140 225.155 166.980 225.325 ;
        RECT 176.850 225.155 184.690 225.325 ;
        RECT 185.140 225.155 192.980 225.325 ;
        RECT 202.850 225.155 210.690 225.325 ;
        RECT 211.140 225.155 218.980 225.325 ;
        RECT 228.850 225.155 236.690 225.325 ;
        RECT 237.140 225.155 244.980 225.325 ;
        RECT 254.850 225.155 262.690 225.325 ;
        RECT 263.140 225.155 270.980 225.325 ;
        RECT 280.850 225.155 288.690 225.325 ;
        RECT 289.140 225.155 296.980 225.325 ;
        RECT 46.850 224.615 54.690 224.785 ;
        RECT 55.140 224.615 62.980 224.785 ;
        RECT 72.850 224.615 80.690 224.785 ;
        RECT 81.140 224.615 88.980 224.785 ;
        RECT 98.850 224.615 106.690 224.785 ;
        RECT 107.140 224.615 114.980 224.785 ;
        RECT 124.850 224.615 132.690 224.785 ;
        RECT 133.140 224.615 140.980 224.785 ;
        RECT 150.850 224.615 158.690 224.785 ;
        RECT 159.140 224.615 166.980 224.785 ;
        RECT 176.850 224.615 184.690 224.785 ;
        RECT 185.140 224.615 192.980 224.785 ;
        RECT 202.850 224.615 210.690 224.785 ;
        RECT 211.140 224.615 218.980 224.785 ;
        RECT 228.850 224.615 236.690 224.785 ;
        RECT 237.140 224.615 244.980 224.785 ;
        RECT 254.850 224.615 262.690 224.785 ;
        RECT 263.140 224.615 270.980 224.785 ;
        RECT 280.850 224.615 288.690 224.785 ;
        RECT 289.140 224.615 296.980 224.785 ;
        RECT 46.850 216.975 54.690 217.145 ;
        RECT 55.140 216.975 62.980 217.145 ;
        RECT 72.850 216.975 80.690 217.145 ;
        RECT 81.140 216.975 88.980 217.145 ;
        RECT 98.850 216.975 106.690 217.145 ;
        RECT 107.140 216.975 114.980 217.145 ;
        RECT 124.850 216.975 132.690 217.145 ;
        RECT 133.140 216.975 140.980 217.145 ;
        RECT 150.850 216.975 158.690 217.145 ;
        RECT 159.140 216.975 166.980 217.145 ;
        RECT 176.850 216.975 184.690 217.145 ;
        RECT 185.140 216.975 192.980 217.145 ;
        RECT 202.850 216.975 210.690 217.145 ;
        RECT 211.140 216.975 218.980 217.145 ;
        RECT 228.850 216.975 236.690 217.145 ;
        RECT 237.140 216.975 244.980 217.145 ;
        RECT 254.850 216.975 262.690 217.145 ;
        RECT 263.140 216.975 270.980 217.145 ;
        RECT 280.850 216.975 288.690 217.145 ;
        RECT 289.140 216.975 296.980 217.145 ;
        RECT 46.850 216.435 54.690 216.605 ;
        RECT 55.140 216.435 62.980 216.605 ;
        RECT 72.850 216.435 80.690 216.605 ;
        RECT 81.140 216.435 88.980 216.605 ;
        RECT 98.850 216.435 106.690 216.605 ;
        RECT 107.140 216.435 114.980 216.605 ;
        RECT 124.850 216.435 132.690 216.605 ;
        RECT 133.140 216.435 140.980 216.605 ;
        RECT 150.850 216.435 158.690 216.605 ;
        RECT 159.140 216.435 166.980 216.605 ;
        RECT 176.850 216.435 184.690 216.605 ;
        RECT 185.140 216.435 192.980 216.605 ;
        RECT 202.850 216.435 210.690 216.605 ;
        RECT 211.140 216.435 218.980 216.605 ;
        RECT 228.850 216.435 236.690 216.605 ;
        RECT 237.140 216.435 244.980 216.605 ;
        RECT 254.850 216.435 262.690 216.605 ;
        RECT 263.140 216.435 270.980 216.605 ;
        RECT 280.850 216.435 288.690 216.605 ;
        RECT 289.140 216.435 296.980 216.605 ;
        RECT 46.850 208.795 54.690 208.965 ;
        RECT 55.140 208.795 62.980 208.965 ;
        RECT 72.850 208.795 80.690 208.965 ;
        RECT 81.140 208.795 88.980 208.965 ;
        RECT 98.850 208.795 106.690 208.965 ;
        RECT 107.140 208.795 114.980 208.965 ;
        RECT 124.850 208.795 132.690 208.965 ;
        RECT 133.140 208.795 140.980 208.965 ;
        RECT 150.850 208.795 158.690 208.965 ;
        RECT 159.140 208.795 166.980 208.965 ;
        RECT 176.850 208.795 184.690 208.965 ;
        RECT 185.140 208.795 192.980 208.965 ;
        RECT 202.850 208.795 210.690 208.965 ;
        RECT 211.140 208.795 218.980 208.965 ;
        RECT 228.850 208.795 236.690 208.965 ;
        RECT 237.140 208.795 244.980 208.965 ;
        RECT 254.850 208.795 262.690 208.965 ;
        RECT 263.140 208.795 270.980 208.965 ;
        RECT 280.850 208.795 288.690 208.965 ;
        RECT 289.140 208.795 296.980 208.965 ;
        RECT 46.850 208.255 54.690 208.425 ;
        RECT 55.140 208.255 62.980 208.425 ;
        RECT 72.850 208.255 80.690 208.425 ;
        RECT 81.140 208.255 88.980 208.425 ;
        RECT 98.850 208.255 106.690 208.425 ;
        RECT 107.140 208.255 114.980 208.425 ;
        RECT 124.850 208.255 132.690 208.425 ;
        RECT 133.140 208.255 140.980 208.425 ;
        RECT 150.850 208.255 158.690 208.425 ;
        RECT 159.140 208.255 166.980 208.425 ;
        RECT 176.850 208.255 184.690 208.425 ;
        RECT 185.140 208.255 192.980 208.425 ;
        RECT 202.850 208.255 210.690 208.425 ;
        RECT 211.140 208.255 218.980 208.425 ;
        RECT 228.850 208.255 236.690 208.425 ;
        RECT 237.140 208.255 244.980 208.425 ;
        RECT 254.850 208.255 262.690 208.425 ;
        RECT 263.140 208.255 270.980 208.425 ;
        RECT 280.850 208.255 288.690 208.425 ;
        RECT 289.140 208.255 296.980 208.425 ;
        RECT 46.850 200.615 54.690 200.785 ;
        RECT 55.140 200.615 62.980 200.785 ;
        RECT 72.850 200.615 80.690 200.785 ;
        RECT 81.140 200.615 88.980 200.785 ;
        RECT 98.850 200.615 106.690 200.785 ;
        RECT 107.140 200.615 114.980 200.785 ;
        RECT 124.850 200.615 132.690 200.785 ;
        RECT 133.140 200.615 140.980 200.785 ;
        RECT 150.850 200.615 158.690 200.785 ;
        RECT 159.140 200.615 166.980 200.785 ;
        RECT 176.850 200.615 184.690 200.785 ;
        RECT 185.140 200.615 192.980 200.785 ;
        RECT 202.850 200.615 210.690 200.785 ;
        RECT 211.140 200.615 218.980 200.785 ;
        RECT 228.850 200.615 236.690 200.785 ;
        RECT 237.140 200.615 244.980 200.785 ;
        RECT 254.850 200.615 262.690 200.785 ;
        RECT 263.140 200.615 270.980 200.785 ;
        RECT 280.850 200.615 288.690 200.785 ;
        RECT 289.140 200.615 296.980 200.785 ;
        RECT 46.850 200.075 54.690 200.245 ;
        RECT 55.140 200.075 62.980 200.245 ;
        RECT 72.850 200.075 80.690 200.245 ;
        RECT 81.140 200.075 88.980 200.245 ;
        RECT 98.850 200.075 106.690 200.245 ;
        RECT 107.140 200.075 114.980 200.245 ;
        RECT 124.850 200.075 132.690 200.245 ;
        RECT 133.140 200.075 140.980 200.245 ;
        RECT 150.850 200.075 158.690 200.245 ;
        RECT 159.140 200.075 166.980 200.245 ;
        RECT 176.850 200.075 184.690 200.245 ;
        RECT 185.140 200.075 192.980 200.245 ;
        RECT 202.850 200.075 210.690 200.245 ;
        RECT 211.140 200.075 218.980 200.245 ;
        RECT 228.850 200.075 236.690 200.245 ;
        RECT 237.140 200.075 244.980 200.245 ;
        RECT 254.850 200.075 262.690 200.245 ;
        RECT 263.140 200.075 270.980 200.245 ;
        RECT 280.850 200.075 288.690 200.245 ;
        RECT 289.140 200.075 296.980 200.245 ;
        RECT 46.850 192.435 54.690 192.605 ;
        RECT 55.140 192.435 62.980 192.605 ;
        RECT 72.850 192.435 80.690 192.605 ;
        RECT 81.140 192.435 88.980 192.605 ;
        RECT 98.850 192.435 106.690 192.605 ;
        RECT 107.140 192.435 114.980 192.605 ;
        RECT 124.850 192.435 132.690 192.605 ;
        RECT 133.140 192.435 140.980 192.605 ;
        RECT 150.850 192.435 158.690 192.605 ;
        RECT 159.140 192.435 166.980 192.605 ;
        RECT 176.850 192.435 184.690 192.605 ;
        RECT 185.140 192.435 192.980 192.605 ;
        RECT 202.850 192.435 210.690 192.605 ;
        RECT 211.140 192.435 218.980 192.605 ;
        RECT 228.850 192.435 236.690 192.605 ;
        RECT 237.140 192.435 244.980 192.605 ;
        RECT 254.850 192.435 262.690 192.605 ;
        RECT 263.140 192.435 270.980 192.605 ;
        RECT 280.850 192.435 288.690 192.605 ;
        RECT 289.140 192.435 296.980 192.605 ;
        RECT 46.850 191.895 54.690 192.065 ;
        RECT 55.140 191.895 62.980 192.065 ;
        RECT 72.850 191.895 80.690 192.065 ;
        RECT 81.140 191.895 88.980 192.065 ;
        RECT 98.850 191.895 106.690 192.065 ;
        RECT 107.140 191.895 114.980 192.065 ;
        RECT 124.850 191.895 132.690 192.065 ;
        RECT 133.140 191.895 140.980 192.065 ;
        RECT 150.850 191.895 158.690 192.065 ;
        RECT 159.140 191.895 166.980 192.065 ;
        RECT 176.850 191.895 184.690 192.065 ;
        RECT 185.140 191.895 192.980 192.065 ;
        RECT 202.850 191.895 210.690 192.065 ;
        RECT 211.140 191.895 218.980 192.065 ;
        RECT 228.850 191.895 236.690 192.065 ;
        RECT 237.140 191.895 244.980 192.065 ;
        RECT 254.850 191.895 262.690 192.065 ;
        RECT 263.140 191.895 270.980 192.065 ;
        RECT 280.850 191.895 288.690 192.065 ;
        RECT 289.140 191.895 296.980 192.065 ;
        RECT 46.850 184.255 54.690 184.425 ;
        RECT 55.140 184.255 62.980 184.425 ;
        RECT 72.850 184.255 80.690 184.425 ;
        RECT 81.140 184.255 88.980 184.425 ;
        RECT 98.850 184.255 106.690 184.425 ;
        RECT 107.140 184.255 114.980 184.425 ;
        RECT 124.850 184.255 132.690 184.425 ;
        RECT 133.140 184.255 140.980 184.425 ;
        RECT 150.850 184.255 158.690 184.425 ;
        RECT 159.140 184.255 166.980 184.425 ;
        RECT 176.850 184.255 184.690 184.425 ;
        RECT 185.140 184.255 192.980 184.425 ;
        RECT 202.850 184.255 210.690 184.425 ;
        RECT 211.140 184.255 218.980 184.425 ;
        RECT 228.850 184.255 236.690 184.425 ;
        RECT 237.140 184.255 244.980 184.425 ;
        RECT 254.850 184.255 262.690 184.425 ;
        RECT 263.140 184.255 270.980 184.425 ;
        RECT 280.850 184.255 288.690 184.425 ;
        RECT 289.140 184.255 296.980 184.425 ;
        RECT 46.850 183.715 54.690 183.885 ;
        RECT 55.140 183.715 62.980 183.885 ;
        RECT 72.850 183.715 80.690 183.885 ;
        RECT 81.140 183.715 88.980 183.885 ;
        RECT 98.850 183.715 106.690 183.885 ;
        RECT 107.140 183.715 114.980 183.885 ;
        RECT 124.850 183.715 132.690 183.885 ;
        RECT 133.140 183.715 140.980 183.885 ;
        RECT 150.850 183.715 158.690 183.885 ;
        RECT 159.140 183.715 166.980 183.885 ;
        RECT 176.850 183.715 184.690 183.885 ;
        RECT 185.140 183.715 192.980 183.885 ;
        RECT 202.850 183.715 210.690 183.885 ;
        RECT 211.140 183.715 218.980 183.885 ;
        RECT 228.850 183.715 236.690 183.885 ;
        RECT 237.140 183.715 244.980 183.885 ;
        RECT 254.850 183.715 262.690 183.885 ;
        RECT 263.140 183.715 270.980 183.885 ;
        RECT 280.850 183.715 288.690 183.885 ;
        RECT 289.140 183.715 296.980 183.885 ;
        RECT 46.850 176.075 54.690 176.245 ;
        RECT 55.140 176.075 62.980 176.245 ;
        RECT 72.850 176.075 80.690 176.245 ;
        RECT 81.140 176.075 88.980 176.245 ;
        RECT 98.850 176.075 106.690 176.245 ;
        RECT 107.140 176.075 114.980 176.245 ;
        RECT 124.850 176.075 132.690 176.245 ;
        RECT 133.140 176.075 140.980 176.245 ;
        RECT 150.850 176.075 158.690 176.245 ;
        RECT 159.140 176.075 166.980 176.245 ;
        RECT 176.850 176.075 184.690 176.245 ;
        RECT 185.140 176.075 192.980 176.245 ;
        RECT 202.850 176.075 210.690 176.245 ;
        RECT 211.140 176.075 218.980 176.245 ;
        RECT 228.850 176.075 236.690 176.245 ;
        RECT 237.140 176.075 244.980 176.245 ;
        RECT 254.850 176.075 262.690 176.245 ;
        RECT 263.140 176.075 270.980 176.245 ;
        RECT 280.850 176.075 288.690 176.245 ;
        RECT 289.140 176.075 296.980 176.245 ;
        RECT 46.850 175.535 54.690 175.705 ;
        RECT 55.140 175.535 62.980 175.705 ;
        RECT 72.850 175.535 80.690 175.705 ;
        RECT 81.140 175.535 88.980 175.705 ;
        RECT 98.850 175.535 106.690 175.705 ;
        RECT 107.140 175.535 114.980 175.705 ;
        RECT 124.850 175.535 132.690 175.705 ;
        RECT 133.140 175.535 140.980 175.705 ;
        RECT 150.850 175.535 158.690 175.705 ;
        RECT 159.140 175.535 166.980 175.705 ;
        RECT 176.850 175.535 184.690 175.705 ;
        RECT 185.140 175.535 192.980 175.705 ;
        RECT 202.850 175.535 210.690 175.705 ;
        RECT 211.140 175.535 218.980 175.705 ;
        RECT 228.850 175.535 236.690 175.705 ;
        RECT 237.140 175.535 244.980 175.705 ;
        RECT 254.850 175.535 262.690 175.705 ;
        RECT 263.140 175.535 270.980 175.705 ;
        RECT 280.850 175.535 288.690 175.705 ;
        RECT 289.140 175.535 296.980 175.705 ;
        RECT 46.850 167.895 54.690 168.065 ;
        RECT 55.140 167.895 62.980 168.065 ;
        RECT 72.850 167.895 80.690 168.065 ;
        RECT 81.140 167.895 88.980 168.065 ;
        RECT 98.850 167.895 106.690 168.065 ;
        RECT 107.140 167.895 114.980 168.065 ;
        RECT 124.850 167.895 132.690 168.065 ;
        RECT 133.140 167.895 140.980 168.065 ;
        RECT 150.850 167.895 158.690 168.065 ;
        RECT 159.140 167.895 166.980 168.065 ;
        RECT 176.850 167.895 184.690 168.065 ;
        RECT 185.140 167.895 192.980 168.065 ;
        RECT 202.850 167.895 210.690 168.065 ;
        RECT 211.140 167.895 218.980 168.065 ;
        RECT 228.850 167.895 236.690 168.065 ;
        RECT 237.140 167.895 244.980 168.065 ;
        RECT 254.850 167.895 262.690 168.065 ;
        RECT 263.140 167.895 270.980 168.065 ;
        RECT 280.850 167.895 288.690 168.065 ;
        RECT 289.140 167.895 296.980 168.065 ;
        RECT 168.430 160.230 168.600 160.400 ;
        RECT 174.440 160.440 174.810 160.800 ;
        RECT 173.090 155.590 173.460 155.920 ;
        RECT 386.380 148.990 386.740 151.150 ;
        RECT 387.990 149.000 388.350 151.160 ;
        RECT 129.340 137.285 129.510 137.455 ;
        RECT 151.240 136.845 151.410 137.015 ;
        RECT 172.030 136.615 172.200 136.785 ;
        RECT 120.870 136.395 124.790 136.565 ;
        RECT 129.560 135.820 129.730 136.600 ;
        RECT 142.770 135.955 146.690 136.125 ;
        RECT 151.460 135.380 151.630 136.160 ;
        RECT 163.560 135.725 167.480 135.895 ;
        RECT 172.250 135.150 172.420 135.930 ;
        RECT 121.890 132.830 122.060 133.000 ;
        RECT 129.260 132.780 129.430 132.950 ;
        RECT 129.480 132.295 129.650 132.465 ;
        RECT 143.790 132.390 143.960 132.560 ;
        RECT 151.160 132.340 151.330 132.510 ;
        RECT 164.580 132.160 164.750 132.330 ;
        RECT 171.950 132.110 172.120 132.280 ;
        RECT 129.260 131.810 129.430 131.980 ;
        RECT 151.380 131.855 151.550 132.025 ;
        RECT 172.170 131.625 172.340 131.795 ;
        RECT 151.160 131.370 151.330 131.540 ;
        RECT 171.950 131.140 172.120 131.310 ;
        RECT 311.590 131.750 311.810 131.960 ;
        RECT 318.385 131.910 318.555 132.080 ;
        RECT 320.380 131.140 320.580 132.340 ;
        RECT 323.420 131.950 323.630 132.160 ;
        RECT 325.305 131.810 325.475 131.980 ;
        RECT 332.150 131.100 332.330 131.290 ;
        RECT 334.070 131.160 334.280 132.380 ;
        RECT 121.890 125.280 122.060 125.450 ;
        RECT 321.550 125.710 321.870 126.110 ;
        RECT 323.415 125.710 323.585 125.880 ;
        RECT 143.790 124.840 143.960 125.010 ;
        RECT 164.580 124.610 164.750 124.780 ;
        RECT 330.220 124.970 330.440 126.500 ;
        RECT 332.180 125.090 332.380 126.260 ;
        RECT 386.390 123.200 386.750 125.360 ;
        RECT 114.950 116.610 116.935 116.800 ;
        RECT 117.605 116.610 119.590 116.800 ;
        RECT 121.100 116.590 123.085 116.780 ;
        RECT 386.260 116.680 386.620 118.840 ;
        RECT 387.860 116.680 388.220 118.840 ;
        RECT 118.280 114.870 120.265 115.060 ;
        RECT 44.530 71.730 44.900 72.180 ;
        RECT 81.450 72.055 81.620 72.225 ;
        RECT 47.210 71.340 47.620 71.750 ;
        RECT 72.980 71.165 76.900 71.335 ;
        RECT 45.790 70.290 47.350 70.460 ;
        RECT 81.670 70.590 81.840 71.370 ;
        RECT 43.740 69.770 44.360 69.940 ;
        RECT 27.245 69.280 27.415 69.450 ;
        RECT 29.565 69.280 29.735 69.450 ;
        RECT 45.980 69.270 47.550 69.440 ;
        RECT 47.110 68.260 47.520 68.670 ;
        RECT 27.275 66.750 27.445 66.920 ;
        RECT 29.595 66.750 29.765 66.920 ;
        RECT 45.830 67.230 47.390 67.400 ;
        RECT 74.000 67.600 74.170 67.770 ;
        RECT 81.370 67.550 81.540 67.720 ;
        RECT 81.590 67.065 81.760 67.235 ;
        RECT 43.780 66.710 44.400 66.880 ;
        RECT 81.370 66.580 81.540 66.750 ;
        RECT 46.020 66.210 47.590 66.380 ;
        RECT 47.140 65.370 47.550 65.780 ;
        RECT 27.265 64.160 27.435 64.330 ;
        RECT 29.585 64.160 29.755 64.330 ;
        RECT 45.810 64.340 47.370 64.510 ;
        RECT 43.760 63.820 44.380 63.990 ;
        RECT 46.000 63.320 47.570 63.490 ;
        RECT 47.170 62.490 47.580 62.900 ;
        RECT 27.265 61.610 27.435 61.780 ;
        RECT 29.585 61.610 29.755 61.780 ;
        RECT 21.210 60.990 21.380 61.210 ;
        RECT 25.000 60.520 25.170 60.740 ;
        RECT 45.850 61.470 47.410 61.640 ;
        RECT 43.800 60.950 44.420 61.120 ;
        RECT 21.210 60.030 21.380 60.250 ;
        RECT 25.000 59.560 25.170 59.780 ;
        RECT 46.040 60.450 47.610 60.620 ;
        RECT 74.000 60.050 74.170 60.220 ;
        RECT 47.150 59.620 47.560 60.030 ;
        RECT 21.210 59.080 21.380 59.300 ;
        RECT 27.265 59.060 27.435 59.230 ;
        RECT 29.585 59.060 29.755 59.230 ;
        RECT 25.000 58.570 25.170 58.790 ;
        RECT 25.000 57.630 25.170 57.850 ;
        RECT 45.850 58.580 47.410 58.750 ;
        RECT 43.800 58.060 44.420 58.230 ;
        RECT 46.040 57.560 47.610 57.730 ;
        RECT 27.265 56.510 27.435 56.680 ;
        RECT 29.585 56.510 29.755 56.680 ;
        RECT 47.160 56.710 47.570 57.120 ;
        RECT 45.850 55.690 47.410 55.860 ;
        RECT 43.800 55.170 44.420 55.340 ;
        RECT 27.265 53.960 27.435 54.130 ;
        RECT 29.585 53.960 29.755 54.130 ;
        RECT 46.040 54.670 47.610 54.840 ;
        RECT 47.260 53.800 47.670 54.210 ;
        RECT 45.870 52.780 47.430 52.950 ;
        RECT 43.820 52.260 44.440 52.430 ;
        RECT 27.265 51.410 27.435 51.580 ;
        RECT 29.585 51.410 29.755 51.580 ;
        RECT 46.060 51.760 47.630 51.930 ;
        RECT 47.240 50.920 47.650 51.330 ;
        RECT 45.850 49.900 47.410 50.070 ;
        RECT 43.800 49.380 44.420 49.550 ;
        RECT 27.265 48.860 27.435 49.030 ;
        RECT 29.585 48.860 29.755 49.030 ;
        RECT 46.040 48.880 47.610 49.050 ;
        RECT 43.440 48.420 43.750 48.740 ;
        RECT 45.830 47.050 47.390 47.220 ;
        RECT 43.780 46.530 44.400 46.700 ;
        RECT 81.840 46.305 82.010 46.475 ;
        RECT 46.020 46.030 47.590 46.200 ;
        RECT 73.370 45.415 77.290 45.585 ;
        RECT 82.060 44.840 82.230 45.620 ;
        RECT 74.390 41.850 74.560 42.020 ;
        RECT 81.760 41.800 81.930 41.970 ;
        RECT 81.980 41.315 82.150 41.485 ;
        RECT 81.760 40.830 81.930 41.000 ;
        RECT 74.390 34.300 74.560 34.470 ;
        RECT 116.160 110.480 116.330 110.930 ;
        RECT 116.960 109.735 117.880 109.905 ;
        RECT 119.250 109.735 120.170 109.905 ;
        RECT 121.540 109.735 122.460 109.905 ;
        RECT 116.190 108.780 116.360 109.220 ;
        RECT 118.480 108.780 118.650 109.220 ;
        RECT 120.770 108.780 120.940 109.220 ;
        RECT 123.060 108.780 123.230 109.220 ;
        RECT 116.960 108.095 117.880 108.265 ;
        RECT 119.250 108.095 120.170 108.265 ;
        RECT 121.540 108.095 122.460 108.265 ;
        RECT 115.580 104.685 117.500 104.855 ;
        RECT 131.420 105.465 133.340 105.635 ;
        RECT 115.580 103.045 117.500 103.215 ;
        RECT 131.420 103.825 133.340 103.995 ;
        RECT 142.340 105.055 144.260 105.225 ;
        RECT 142.340 103.415 144.260 103.585 ;
        RECT 122.920 100.510 123.230 100.850 ;
        RECT 130.125 100.580 130.600 100.975 ;
        RECT 135.540 100.440 135.950 100.810 ;
        RECT 143.490 100.580 143.965 100.975 ;
        RECT 145.700 100.580 146.140 100.890 ;
        RECT 149.670 100.650 150.510 101.540 ;
        RECT 112.560 99.815 112.730 99.985 ;
        RECT 113.850 99.815 114.020 99.985 ;
        RECT 115.140 99.815 115.310 99.985 ;
        RECT 116.430 99.815 116.600 99.985 ;
        RECT 117.720 99.815 117.890 99.985 ;
        RECT 119.010 99.815 119.180 99.985 ;
        RECT 120.300 99.815 120.470 99.985 ;
        RECT 121.590 99.815 121.760 99.985 ;
        RECT 112.560 98.265 112.730 98.435 ;
        RECT 112.560 97.725 112.730 97.895 ;
        RECT 112.560 96.175 112.730 96.345 ;
        RECT 112.560 95.635 112.730 95.805 ;
        RECT 112.560 94.085 112.730 94.255 ;
        RECT 112.560 93.545 112.730 93.715 ;
        RECT 112.560 91.995 112.730 92.165 ;
        RECT 112.560 91.455 112.730 91.625 ;
        RECT 112.560 89.905 112.730 90.075 ;
        RECT 112.560 89.365 112.730 89.535 ;
        RECT 112.560 87.815 112.730 87.985 ;
        RECT 112.560 87.275 112.730 87.445 ;
        RECT 112.560 85.725 112.730 85.895 ;
        RECT 113.850 98.265 114.020 98.435 ;
        RECT 113.850 97.725 114.020 97.895 ;
        RECT 113.850 96.175 114.020 96.345 ;
        RECT 113.850 95.635 114.020 95.805 ;
        RECT 113.850 94.085 114.020 94.255 ;
        RECT 113.850 93.545 114.020 93.715 ;
        RECT 113.850 91.995 114.020 92.165 ;
        RECT 113.850 91.455 114.020 91.625 ;
        RECT 113.850 89.905 114.020 90.075 ;
        RECT 113.850 89.365 114.020 89.535 ;
        RECT 113.850 87.815 114.020 87.985 ;
        RECT 113.850 87.275 114.020 87.445 ;
        RECT 113.850 85.725 114.020 85.895 ;
        RECT 115.140 98.265 115.310 98.435 ;
        RECT 115.140 97.725 115.310 97.895 ;
        RECT 115.140 96.175 115.310 96.345 ;
        RECT 115.140 95.635 115.310 95.805 ;
        RECT 115.140 94.085 115.310 94.255 ;
        RECT 115.140 93.545 115.310 93.715 ;
        RECT 115.140 91.995 115.310 92.165 ;
        RECT 115.140 91.455 115.310 91.625 ;
        RECT 115.140 89.905 115.310 90.075 ;
        RECT 115.140 89.365 115.310 89.535 ;
        RECT 115.140 87.815 115.310 87.985 ;
        RECT 115.140 87.275 115.310 87.445 ;
        RECT 115.140 85.725 115.310 85.895 ;
        RECT 116.430 98.265 116.600 98.435 ;
        RECT 116.430 97.725 116.600 97.895 ;
        RECT 116.430 96.175 116.600 96.345 ;
        RECT 116.430 95.635 116.600 95.805 ;
        RECT 116.430 94.085 116.600 94.255 ;
        RECT 116.430 93.545 116.600 93.715 ;
        RECT 116.430 91.995 116.600 92.165 ;
        RECT 116.430 91.455 116.600 91.625 ;
        RECT 116.430 89.905 116.600 90.075 ;
        RECT 116.430 89.365 116.600 89.535 ;
        RECT 116.430 87.815 116.600 87.985 ;
        RECT 116.430 87.275 116.600 87.445 ;
        RECT 116.430 85.725 116.600 85.895 ;
        RECT 117.720 98.265 117.890 98.435 ;
        RECT 117.720 97.725 117.890 97.895 ;
        RECT 117.720 96.175 117.890 96.345 ;
        RECT 117.720 95.635 117.890 95.805 ;
        RECT 117.720 94.085 117.890 94.255 ;
        RECT 117.720 93.545 117.890 93.715 ;
        RECT 117.720 91.995 117.890 92.165 ;
        RECT 117.720 91.455 117.890 91.625 ;
        RECT 117.720 89.905 117.890 90.075 ;
        RECT 117.720 89.365 117.890 89.535 ;
        RECT 117.720 87.815 117.890 87.985 ;
        RECT 117.720 87.275 117.890 87.445 ;
        RECT 117.720 85.725 117.890 85.895 ;
        RECT 119.010 98.265 119.180 98.435 ;
        RECT 119.010 97.725 119.180 97.895 ;
        RECT 119.010 96.175 119.180 96.345 ;
        RECT 119.010 95.635 119.180 95.805 ;
        RECT 119.010 94.085 119.180 94.255 ;
        RECT 119.010 93.545 119.180 93.715 ;
        RECT 119.010 91.995 119.180 92.165 ;
        RECT 119.010 91.455 119.180 91.625 ;
        RECT 119.010 89.905 119.180 90.075 ;
        RECT 119.010 89.365 119.180 89.535 ;
        RECT 119.010 87.815 119.180 87.985 ;
        RECT 119.010 87.275 119.180 87.445 ;
        RECT 119.010 85.725 119.180 85.895 ;
        RECT 120.300 98.265 120.470 98.435 ;
        RECT 120.300 97.725 120.470 97.895 ;
        RECT 120.300 96.175 120.470 96.345 ;
        RECT 120.300 95.635 120.470 95.805 ;
        RECT 120.300 94.085 120.470 94.255 ;
        RECT 120.300 93.545 120.470 93.715 ;
        RECT 120.300 91.995 120.470 92.165 ;
        RECT 120.300 91.455 120.470 91.625 ;
        RECT 120.300 89.905 120.470 90.075 ;
        RECT 120.300 89.365 120.470 89.535 ;
        RECT 120.300 87.815 120.470 87.985 ;
        RECT 120.300 87.275 120.470 87.445 ;
        RECT 120.300 85.725 120.470 85.895 ;
        RECT 121.590 98.265 121.760 98.435 ;
        RECT 121.590 97.725 121.760 97.895 ;
        RECT 121.590 96.175 121.760 96.345 ;
        RECT 121.590 95.635 121.760 95.805 ;
        RECT 121.590 94.085 121.760 94.255 ;
        RECT 121.590 93.545 121.760 93.715 ;
        RECT 121.590 91.995 121.760 92.165 ;
        RECT 121.590 91.455 121.760 91.625 ;
        RECT 121.590 89.905 121.760 90.075 ;
        RECT 121.590 89.365 121.760 89.535 ;
        RECT 121.590 87.815 121.760 87.985 ;
        RECT 121.590 87.275 121.760 87.445 ;
        RECT 121.590 85.725 121.760 85.895 ;
        RECT 125.910 99.815 126.080 99.985 ;
        RECT 127.200 99.815 127.370 99.985 ;
        RECT 128.490 99.815 128.660 99.985 ;
        RECT 129.780 99.815 129.950 99.985 ;
        RECT 131.070 99.815 131.240 99.985 ;
        RECT 132.360 99.815 132.530 99.985 ;
        RECT 133.650 99.815 133.820 99.985 ;
        RECT 134.940 99.815 135.110 99.985 ;
        RECT 125.910 98.265 126.080 98.435 ;
        RECT 125.910 97.725 126.080 97.895 ;
        RECT 125.910 96.175 126.080 96.345 ;
        RECT 125.910 95.635 126.080 95.805 ;
        RECT 125.910 94.085 126.080 94.255 ;
        RECT 125.910 93.545 126.080 93.715 ;
        RECT 125.910 91.995 126.080 92.165 ;
        RECT 125.910 91.455 126.080 91.625 ;
        RECT 125.910 89.905 126.080 90.075 ;
        RECT 125.910 89.365 126.080 89.535 ;
        RECT 125.910 87.815 126.080 87.985 ;
        RECT 125.910 87.275 126.080 87.445 ;
        RECT 125.910 85.725 126.080 85.895 ;
        RECT 127.200 98.265 127.370 98.435 ;
        RECT 127.200 97.725 127.370 97.895 ;
        RECT 127.200 96.175 127.370 96.345 ;
        RECT 127.200 95.635 127.370 95.805 ;
        RECT 127.200 94.085 127.370 94.255 ;
        RECT 127.200 93.545 127.370 93.715 ;
        RECT 127.200 91.995 127.370 92.165 ;
        RECT 127.200 91.455 127.370 91.625 ;
        RECT 127.200 89.905 127.370 90.075 ;
        RECT 127.200 89.365 127.370 89.535 ;
        RECT 127.200 87.815 127.370 87.985 ;
        RECT 127.200 87.275 127.370 87.445 ;
        RECT 127.200 85.725 127.370 85.895 ;
        RECT 128.490 98.265 128.660 98.435 ;
        RECT 128.490 97.725 128.660 97.895 ;
        RECT 128.490 96.175 128.660 96.345 ;
        RECT 128.490 95.635 128.660 95.805 ;
        RECT 128.490 94.085 128.660 94.255 ;
        RECT 128.490 93.545 128.660 93.715 ;
        RECT 128.490 91.995 128.660 92.165 ;
        RECT 128.490 91.455 128.660 91.625 ;
        RECT 128.490 89.905 128.660 90.075 ;
        RECT 128.490 89.365 128.660 89.535 ;
        RECT 128.490 87.815 128.660 87.985 ;
        RECT 128.490 87.275 128.660 87.445 ;
        RECT 128.490 85.725 128.660 85.895 ;
        RECT 129.780 98.265 129.950 98.435 ;
        RECT 129.780 97.725 129.950 97.895 ;
        RECT 129.780 96.175 129.950 96.345 ;
        RECT 129.780 95.635 129.950 95.805 ;
        RECT 129.780 94.085 129.950 94.255 ;
        RECT 129.780 93.545 129.950 93.715 ;
        RECT 129.780 91.995 129.950 92.165 ;
        RECT 129.780 91.455 129.950 91.625 ;
        RECT 129.780 89.905 129.950 90.075 ;
        RECT 129.780 89.365 129.950 89.535 ;
        RECT 129.780 87.815 129.950 87.985 ;
        RECT 129.780 87.275 129.950 87.445 ;
        RECT 129.780 85.725 129.950 85.895 ;
        RECT 131.070 98.265 131.240 98.435 ;
        RECT 131.070 97.725 131.240 97.895 ;
        RECT 131.070 96.175 131.240 96.345 ;
        RECT 131.070 95.635 131.240 95.805 ;
        RECT 131.070 94.085 131.240 94.255 ;
        RECT 131.070 93.545 131.240 93.715 ;
        RECT 131.070 91.995 131.240 92.165 ;
        RECT 131.070 91.455 131.240 91.625 ;
        RECT 131.070 89.905 131.240 90.075 ;
        RECT 131.070 89.365 131.240 89.535 ;
        RECT 131.070 87.815 131.240 87.985 ;
        RECT 131.070 87.275 131.240 87.445 ;
        RECT 131.070 85.725 131.240 85.895 ;
        RECT 132.360 98.265 132.530 98.435 ;
        RECT 132.360 97.725 132.530 97.895 ;
        RECT 132.360 96.175 132.530 96.345 ;
        RECT 132.360 95.635 132.530 95.805 ;
        RECT 132.360 94.085 132.530 94.255 ;
        RECT 132.360 93.545 132.530 93.715 ;
        RECT 132.360 91.995 132.530 92.165 ;
        RECT 132.360 91.455 132.530 91.625 ;
        RECT 132.360 89.905 132.530 90.075 ;
        RECT 132.360 89.365 132.530 89.535 ;
        RECT 132.360 87.815 132.530 87.985 ;
        RECT 132.360 87.275 132.530 87.445 ;
        RECT 132.360 85.725 132.530 85.895 ;
        RECT 133.650 98.265 133.820 98.435 ;
        RECT 133.650 97.725 133.820 97.895 ;
        RECT 133.650 96.175 133.820 96.345 ;
        RECT 133.650 95.635 133.820 95.805 ;
        RECT 133.650 94.085 133.820 94.255 ;
        RECT 133.650 93.545 133.820 93.715 ;
        RECT 133.650 91.995 133.820 92.165 ;
        RECT 133.650 91.455 133.820 91.625 ;
        RECT 133.650 89.905 133.820 90.075 ;
        RECT 133.650 89.365 133.820 89.535 ;
        RECT 133.650 87.815 133.820 87.985 ;
        RECT 133.650 87.275 133.820 87.445 ;
        RECT 133.650 85.725 133.820 85.895 ;
        RECT 134.940 98.265 135.110 98.435 ;
        RECT 134.940 97.725 135.110 97.895 ;
        RECT 134.940 96.175 135.110 96.345 ;
        RECT 134.940 95.635 135.110 95.805 ;
        RECT 134.940 94.085 135.110 94.255 ;
        RECT 134.940 93.545 135.110 93.715 ;
        RECT 134.940 91.995 135.110 92.165 ;
        RECT 134.940 91.455 135.110 91.625 ;
        RECT 134.940 89.905 135.110 90.075 ;
        RECT 134.940 89.365 135.110 89.535 ;
        RECT 134.940 87.815 135.110 87.985 ;
        RECT 134.940 87.275 135.110 87.445 ;
        RECT 134.940 85.725 135.110 85.895 ;
        RECT 139.225 99.820 139.395 99.990 ;
        RECT 140.515 99.820 140.685 99.990 ;
        RECT 141.805 99.820 141.975 99.990 ;
        RECT 143.095 99.820 143.265 99.990 ;
        RECT 144.385 99.820 144.555 99.990 ;
        RECT 145.675 99.820 145.845 99.990 ;
        RECT 146.965 99.820 147.135 99.990 ;
        RECT 148.255 99.820 148.425 99.990 ;
        RECT 139.225 98.270 139.395 98.440 ;
        RECT 139.225 97.730 139.395 97.900 ;
        RECT 139.225 96.180 139.395 96.350 ;
        RECT 139.225 95.640 139.395 95.810 ;
        RECT 139.225 94.090 139.395 94.260 ;
        RECT 139.225 93.550 139.395 93.720 ;
        RECT 139.225 92.000 139.395 92.170 ;
        RECT 139.225 91.460 139.395 91.630 ;
        RECT 139.225 89.910 139.395 90.080 ;
        RECT 139.225 89.370 139.395 89.540 ;
        RECT 139.225 87.820 139.395 87.990 ;
        RECT 139.225 87.280 139.395 87.450 ;
        RECT 139.225 85.730 139.395 85.900 ;
        RECT 140.515 98.270 140.685 98.440 ;
        RECT 140.515 97.730 140.685 97.900 ;
        RECT 140.515 96.180 140.685 96.350 ;
        RECT 140.515 95.640 140.685 95.810 ;
        RECT 140.515 94.090 140.685 94.260 ;
        RECT 140.515 93.550 140.685 93.720 ;
        RECT 140.515 92.000 140.685 92.170 ;
        RECT 140.515 91.460 140.685 91.630 ;
        RECT 140.515 89.910 140.685 90.080 ;
        RECT 140.515 89.370 140.685 89.540 ;
        RECT 140.515 87.820 140.685 87.990 ;
        RECT 140.515 87.280 140.685 87.450 ;
        RECT 140.515 85.730 140.685 85.900 ;
        RECT 141.805 98.270 141.975 98.440 ;
        RECT 141.805 97.730 141.975 97.900 ;
        RECT 141.805 96.180 141.975 96.350 ;
        RECT 141.805 95.640 141.975 95.810 ;
        RECT 141.805 94.090 141.975 94.260 ;
        RECT 141.805 93.550 141.975 93.720 ;
        RECT 141.805 92.000 141.975 92.170 ;
        RECT 141.805 91.460 141.975 91.630 ;
        RECT 141.805 89.910 141.975 90.080 ;
        RECT 141.805 89.370 141.975 89.540 ;
        RECT 141.805 87.820 141.975 87.990 ;
        RECT 141.805 87.280 141.975 87.450 ;
        RECT 141.805 85.730 141.975 85.900 ;
        RECT 143.095 98.270 143.265 98.440 ;
        RECT 143.095 97.730 143.265 97.900 ;
        RECT 143.095 96.180 143.265 96.350 ;
        RECT 143.095 95.640 143.265 95.810 ;
        RECT 143.095 94.090 143.265 94.260 ;
        RECT 143.095 93.550 143.265 93.720 ;
        RECT 143.095 92.000 143.265 92.170 ;
        RECT 143.095 91.460 143.265 91.630 ;
        RECT 143.095 89.910 143.265 90.080 ;
        RECT 143.095 89.370 143.265 89.540 ;
        RECT 143.095 87.820 143.265 87.990 ;
        RECT 143.095 87.280 143.265 87.450 ;
        RECT 143.095 85.730 143.265 85.900 ;
        RECT 144.385 98.270 144.555 98.440 ;
        RECT 144.385 97.730 144.555 97.900 ;
        RECT 144.385 96.180 144.555 96.350 ;
        RECT 144.385 95.640 144.555 95.810 ;
        RECT 144.385 94.090 144.555 94.260 ;
        RECT 144.385 93.550 144.555 93.720 ;
        RECT 144.385 92.000 144.555 92.170 ;
        RECT 144.385 91.460 144.555 91.630 ;
        RECT 144.385 89.910 144.555 90.080 ;
        RECT 144.385 89.370 144.555 89.540 ;
        RECT 144.385 87.820 144.555 87.990 ;
        RECT 144.385 87.280 144.555 87.450 ;
        RECT 144.385 85.730 144.555 85.900 ;
        RECT 145.675 98.270 145.845 98.440 ;
        RECT 145.675 97.730 145.845 97.900 ;
        RECT 145.675 96.180 145.845 96.350 ;
        RECT 145.675 95.640 145.845 95.810 ;
        RECT 145.675 94.090 145.845 94.260 ;
        RECT 145.675 93.550 145.845 93.720 ;
        RECT 145.675 92.000 145.845 92.170 ;
        RECT 145.675 91.460 145.845 91.630 ;
        RECT 145.675 89.910 145.845 90.080 ;
        RECT 145.675 89.370 145.845 89.540 ;
        RECT 145.675 87.820 145.845 87.990 ;
        RECT 145.675 87.280 145.845 87.450 ;
        RECT 145.675 85.730 145.845 85.900 ;
        RECT 146.965 98.270 147.135 98.440 ;
        RECT 146.965 97.730 147.135 97.900 ;
        RECT 146.965 96.180 147.135 96.350 ;
        RECT 146.965 95.640 147.135 95.810 ;
        RECT 146.965 94.090 147.135 94.260 ;
        RECT 146.965 93.550 147.135 93.720 ;
        RECT 146.965 92.000 147.135 92.170 ;
        RECT 146.965 91.460 147.135 91.630 ;
        RECT 146.965 89.910 147.135 90.080 ;
        RECT 146.965 89.370 147.135 89.540 ;
        RECT 146.965 87.820 147.135 87.990 ;
        RECT 146.965 87.280 147.135 87.450 ;
        RECT 146.965 85.730 147.135 85.900 ;
        RECT 148.255 98.270 148.425 98.440 ;
        RECT 148.255 97.730 148.425 97.900 ;
        RECT 148.255 96.180 148.425 96.350 ;
        RECT 148.255 95.640 148.425 95.810 ;
        RECT 148.255 94.090 148.425 94.260 ;
        RECT 148.255 93.550 148.425 93.720 ;
        RECT 148.255 92.000 148.425 92.170 ;
        RECT 148.255 91.460 148.425 91.630 ;
        RECT 148.255 89.910 148.425 90.080 ;
        RECT 148.255 89.370 148.425 89.540 ;
        RECT 148.255 87.820 148.425 87.990 ;
        RECT 148.255 87.280 148.425 87.450 ;
        RECT 148.255 85.730 148.425 85.900 ;
        RECT 116.470 83.830 116.890 84.000 ;
        RECT 131.130 83.870 131.550 84.040 ;
        RECT 131.860 83.350 132.110 83.590 ;
        RECT 143.690 83.870 144.110 84.040 ;
        RECT 116.470 82.860 116.890 83.030 ;
        RECT 131.130 82.900 131.550 83.070 ;
        RECT 143.690 82.900 144.110 83.070 ;
        RECT 115.950 76.715 117.870 76.885 ;
        RECT 129.660 76.835 131.580 77.005 ;
        RECT 134.440 75.840 134.970 76.220 ;
        RECT 115.950 75.075 117.870 75.245 ;
        RECT 129.660 75.195 131.580 75.365 ;
        RECT 119.740 74.760 120.090 75.110 ;
        RECT 142.840 76.875 144.760 77.045 ;
        RECT 145.600 75.760 146.200 76.460 ;
        RECT 142.840 75.235 144.760 75.405 ;
        RECT 110.630 71.950 111.420 72.770 ;
        RECT 124.160 71.850 124.750 72.520 ;
        RECT 137.190 71.850 137.750 72.470 ;
        RECT 112.560 71.230 112.730 71.400 ;
        RECT 113.850 71.230 114.020 71.400 ;
        RECT 115.140 71.230 115.310 71.400 ;
        RECT 116.430 71.230 116.600 71.400 ;
        RECT 117.720 71.230 117.890 71.400 ;
        RECT 119.010 71.230 119.180 71.400 ;
        RECT 120.300 71.230 120.470 71.400 ;
        RECT 121.590 71.230 121.760 71.400 ;
        RECT 112.560 69.680 112.730 69.850 ;
        RECT 112.560 69.140 112.730 69.310 ;
        RECT 112.560 67.590 112.730 67.760 ;
        RECT 112.560 67.050 112.730 67.220 ;
        RECT 112.560 65.500 112.730 65.670 ;
        RECT 112.560 64.960 112.730 65.130 ;
        RECT 112.560 63.410 112.730 63.580 ;
        RECT 112.560 62.870 112.730 63.040 ;
        RECT 112.560 61.320 112.730 61.490 ;
        RECT 112.560 60.780 112.730 60.950 ;
        RECT 112.560 59.230 112.730 59.400 ;
        RECT 112.560 58.690 112.730 58.860 ;
        RECT 112.560 57.140 112.730 57.310 ;
        RECT 113.850 69.680 114.020 69.850 ;
        RECT 113.850 69.140 114.020 69.310 ;
        RECT 113.850 67.590 114.020 67.760 ;
        RECT 113.850 67.050 114.020 67.220 ;
        RECT 113.850 65.500 114.020 65.670 ;
        RECT 113.850 64.960 114.020 65.130 ;
        RECT 113.850 63.410 114.020 63.580 ;
        RECT 113.850 62.870 114.020 63.040 ;
        RECT 113.850 61.320 114.020 61.490 ;
        RECT 113.850 60.780 114.020 60.950 ;
        RECT 113.850 59.230 114.020 59.400 ;
        RECT 113.850 58.690 114.020 58.860 ;
        RECT 113.850 57.140 114.020 57.310 ;
        RECT 115.140 69.680 115.310 69.850 ;
        RECT 115.140 69.140 115.310 69.310 ;
        RECT 115.140 67.590 115.310 67.760 ;
        RECT 115.140 67.050 115.310 67.220 ;
        RECT 115.140 65.500 115.310 65.670 ;
        RECT 115.140 64.960 115.310 65.130 ;
        RECT 115.140 63.410 115.310 63.580 ;
        RECT 115.140 62.870 115.310 63.040 ;
        RECT 115.140 61.320 115.310 61.490 ;
        RECT 115.140 60.780 115.310 60.950 ;
        RECT 115.140 59.230 115.310 59.400 ;
        RECT 115.140 58.690 115.310 58.860 ;
        RECT 115.140 57.140 115.310 57.310 ;
        RECT 116.430 69.680 116.600 69.850 ;
        RECT 116.430 69.140 116.600 69.310 ;
        RECT 116.430 67.590 116.600 67.760 ;
        RECT 116.430 67.050 116.600 67.220 ;
        RECT 116.430 65.500 116.600 65.670 ;
        RECT 116.430 64.960 116.600 65.130 ;
        RECT 116.430 63.410 116.600 63.580 ;
        RECT 116.430 62.870 116.600 63.040 ;
        RECT 116.430 61.320 116.600 61.490 ;
        RECT 116.430 60.780 116.600 60.950 ;
        RECT 116.430 59.230 116.600 59.400 ;
        RECT 116.430 58.690 116.600 58.860 ;
        RECT 116.430 57.140 116.600 57.310 ;
        RECT 117.720 69.680 117.890 69.850 ;
        RECT 117.720 69.140 117.890 69.310 ;
        RECT 117.720 67.590 117.890 67.760 ;
        RECT 117.720 67.050 117.890 67.220 ;
        RECT 117.720 65.500 117.890 65.670 ;
        RECT 117.720 64.960 117.890 65.130 ;
        RECT 117.720 63.410 117.890 63.580 ;
        RECT 117.720 62.870 117.890 63.040 ;
        RECT 117.720 61.320 117.890 61.490 ;
        RECT 117.720 60.780 117.890 60.950 ;
        RECT 117.720 59.230 117.890 59.400 ;
        RECT 117.720 58.690 117.890 58.860 ;
        RECT 117.720 57.140 117.890 57.310 ;
        RECT 119.010 69.680 119.180 69.850 ;
        RECT 119.010 69.140 119.180 69.310 ;
        RECT 119.010 67.590 119.180 67.760 ;
        RECT 119.010 67.050 119.180 67.220 ;
        RECT 119.010 65.500 119.180 65.670 ;
        RECT 119.010 64.960 119.180 65.130 ;
        RECT 119.010 63.410 119.180 63.580 ;
        RECT 119.010 62.870 119.180 63.040 ;
        RECT 119.010 61.320 119.180 61.490 ;
        RECT 119.010 60.780 119.180 60.950 ;
        RECT 119.010 59.230 119.180 59.400 ;
        RECT 119.010 58.690 119.180 58.860 ;
        RECT 119.010 57.140 119.180 57.310 ;
        RECT 120.300 69.680 120.470 69.850 ;
        RECT 120.300 69.140 120.470 69.310 ;
        RECT 120.300 67.590 120.470 67.760 ;
        RECT 120.300 67.050 120.470 67.220 ;
        RECT 120.300 65.500 120.470 65.670 ;
        RECT 120.300 64.960 120.470 65.130 ;
        RECT 120.300 63.410 120.470 63.580 ;
        RECT 120.300 62.870 120.470 63.040 ;
        RECT 120.300 61.320 120.470 61.490 ;
        RECT 120.300 60.780 120.470 60.950 ;
        RECT 120.300 59.230 120.470 59.400 ;
        RECT 120.300 58.690 120.470 58.860 ;
        RECT 120.300 57.140 120.470 57.310 ;
        RECT 125.910 71.230 126.080 71.400 ;
        RECT 127.200 71.230 127.370 71.400 ;
        RECT 128.490 71.230 128.660 71.400 ;
        RECT 129.780 71.230 129.950 71.400 ;
        RECT 131.070 71.230 131.240 71.400 ;
        RECT 132.360 71.230 132.530 71.400 ;
        RECT 133.650 71.230 133.820 71.400 ;
        RECT 134.940 71.230 135.110 71.400 ;
        RECT 121.590 69.680 121.760 69.850 ;
        RECT 121.590 69.140 121.760 69.310 ;
        RECT 121.590 67.590 121.760 67.760 ;
        RECT 121.590 67.050 121.760 67.220 ;
        RECT 121.590 65.500 121.760 65.670 ;
        RECT 121.590 64.960 121.760 65.130 ;
        RECT 121.590 63.410 121.760 63.580 ;
        RECT 121.590 62.870 121.760 63.040 ;
        RECT 121.590 61.320 121.760 61.490 ;
        RECT 121.590 60.780 121.760 60.950 ;
        RECT 121.590 59.230 121.760 59.400 ;
        RECT 121.590 58.690 121.760 58.860 ;
        RECT 125.910 69.680 126.080 69.850 ;
        RECT 125.910 69.140 126.080 69.310 ;
        RECT 125.910 67.590 126.080 67.760 ;
        RECT 125.910 67.050 126.080 67.220 ;
        RECT 125.910 65.500 126.080 65.670 ;
        RECT 125.910 64.960 126.080 65.130 ;
        RECT 125.910 63.410 126.080 63.580 ;
        RECT 125.910 62.870 126.080 63.040 ;
        RECT 125.910 61.320 126.080 61.490 ;
        RECT 125.910 60.780 126.080 60.950 ;
        RECT 125.910 59.230 126.080 59.400 ;
        RECT 125.910 58.690 126.080 58.860 ;
        RECT 121.590 57.140 121.760 57.310 ;
        RECT 125.910 57.140 126.080 57.310 ;
        RECT 127.200 69.680 127.370 69.850 ;
        RECT 127.200 69.140 127.370 69.310 ;
        RECT 127.200 67.590 127.370 67.760 ;
        RECT 127.200 67.050 127.370 67.220 ;
        RECT 127.200 65.500 127.370 65.670 ;
        RECT 127.200 64.960 127.370 65.130 ;
        RECT 127.200 63.410 127.370 63.580 ;
        RECT 127.200 62.870 127.370 63.040 ;
        RECT 127.200 61.320 127.370 61.490 ;
        RECT 127.200 60.780 127.370 60.950 ;
        RECT 127.200 59.230 127.370 59.400 ;
        RECT 127.200 58.690 127.370 58.860 ;
        RECT 127.200 57.140 127.370 57.310 ;
        RECT 128.490 69.680 128.660 69.850 ;
        RECT 128.490 69.140 128.660 69.310 ;
        RECT 128.490 67.590 128.660 67.760 ;
        RECT 128.490 67.050 128.660 67.220 ;
        RECT 128.490 65.500 128.660 65.670 ;
        RECT 128.490 64.960 128.660 65.130 ;
        RECT 128.490 63.410 128.660 63.580 ;
        RECT 128.490 62.870 128.660 63.040 ;
        RECT 128.490 61.320 128.660 61.490 ;
        RECT 128.490 60.780 128.660 60.950 ;
        RECT 128.490 59.230 128.660 59.400 ;
        RECT 128.490 58.690 128.660 58.860 ;
        RECT 128.490 57.140 128.660 57.310 ;
        RECT 129.780 69.680 129.950 69.850 ;
        RECT 129.780 69.140 129.950 69.310 ;
        RECT 129.780 67.590 129.950 67.760 ;
        RECT 129.780 67.050 129.950 67.220 ;
        RECT 129.780 65.500 129.950 65.670 ;
        RECT 129.780 64.960 129.950 65.130 ;
        RECT 129.780 63.410 129.950 63.580 ;
        RECT 129.780 62.870 129.950 63.040 ;
        RECT 129.780 61.320 129.950 61.490 ;
        RECT 129.780 60.780 129.950 60.950 ;
        RECT 129.780 59.230 129.950 59.400 ;
        RECT 129.780 58.690 129.950 58.860 ;
        RECT 129.780 57.140 129.950 57.310 ;
        RECT 131.070 69.680 131.240 69.850 ;
        RECT 131.070 69.140 131.240 69.310 ;
        RECT 131.070 67.590 131.240 67.760 ;
        RECT 131.070 67.050 131.240 67.220 ;
        RECT 131.070 65.500 131.240 65.670 ;
        RECT 131.070 64.960 131.240 65.130 ;
        RECT 131.070 63.410 131.240 63.580 ;
        RECT 131.070 62.870 131.240 63.040 ;
        RECT 131.070 61.320 131.240 61.490 ;
        RECT 131.070 60.780 131.240 60.950 ;
        RECT 131.070 59.230 131.240 59.400 ;
        RECT 131.070 58.690 131.240 58.860 ;
        RECT 131.070 57.140 131.240 57.310 ;
        RECT 132.360 69.680 132.530 69.850 ;
        RECT 132.360 69.140 132.530 69.310 ;
        RECT 132.360 67.590 132.530 67.760 ;
        RECT 132.360 67.050 132.530 67.220 ;
        RECT 132.360 65.500 132.530 65.670 ;
        RECT 132.360 64.960 132.530 65.130 ;
        RECT 132.360 63.410 132.530 63.580 ;
        RECT 132.360 62.870 132.530 63.040 ;
        RECT 132.360 61.320 132.530 61.490 ;
        RECT 132.360 60.780 132.530 60.950 ;
        RECT 132.360 59.230 132.530 59.400 ;
        RECT 132.360 58.690 132.530 58.860 ;
        RECT 132.360 57.140 132.530 57.310 ;
        RECT 133.650 69.680 133.820 69.850 ;
        RECT 133.650 69.140 133.820 69.310 ;
        RECT 133.650 67.590 133.820 67.760 ;
        RECT 133.650 67.050 133.820 67.220 ;
        RECT 133.650 65.500 133.820 65.670 ;
        RECT 133.650 64.960 133.820 65.130 ;
        RECT 133.650 63.410 133.820 63.580 ;
        RECT 133.650 62.870 133.820 63.040 ;
        RECT 133.650 61.320 133.820 61.490 ;
        RECT 133.650 60.780 133.820 60.950 ;
        RECT 133.650 59.230 133.820 59.400 ;
        RECT 133.650 58.690 133.820 58.860 ;
        RECT 133.650 57.140 133.820 57.310 ;
        RECT 139.225 71.235 139.395 71.405 ;
        RECT 140.515 71.235 140.685 71.405 ;
        RECT 141.805 71.235 141.975 71.405 ;
        RECT 143.095 71.235 143.265 71.405 ;
        RECT 144.385 71.235 144.555 71.405 ;
        RECT 145.675 71.235 145.845 71.405 ;
        RECT 146.965 71.235 147.135 71.405 ;
        RECT 148.255 71.235 148.425 71.405 ;
        RECT 134.940 69.680 135.110 69.850 ;
        RECT 134.940 69.140 135.110 69.310 ;
        RECT 134.940 67.590 135.110 67.760 ;
        RECT 134.940 67.050 135.110 67.220 ;
        RECT 134.940 65.500 135.110 65.670 ;
        RECT 134.940 64.960 135.110 65.130 ;
        RECT 134.940 63.410 135.110 63.580 ;
        RECT 134.940 62.870 135.110 63.040 ;
        RECT 134.940 61.320 135.110 61.490 ;
        RECT 134.940 60.780 135.110 60.950 ;
        RECT 134.940 59.230 135.110 59.400 ;
        RECT 134.940 58.690 135.110 58.860 ;
        RECT 139.225 69.685 139.395 69.855 ;
        RECT 139.225 69.145 139.395 69.315 ;
        RECT 139.225 67.595 139.395 67.765 ;
        RECT 139.225 67.055 139.395 67.225 ;
        RECT 139.225 65.505 139.395 65.675 ;
        RECT 139.225 64.965 139.395 65.135 ;
        RECT 139.225 63.415 139.395 63.585 ;
        RECT 139.225 62.875 139.395 63.045 ;
        RECT 139.225 61.325 139.395 61.495 ;
        RECT 139.225 60.785 139.395 60.955 ;
        RECT 139.225 59.235 139.395 59.405 ;
        RECT 139.225 58.695 139.395 58.865 ;
        RECT 134.940 57.140 135.110 57.310 ;
        RECT 139.225 57.145 139.395 57.315 ;
        RECT 140.515 69.685 140.685 69.855 ;
        RECT 140.515 69.145 140.685 69.315 ;
        RECT 140.515 67.595 140.685 67.765 ;
        RECT 140.515 67.055 140.685 67.225 ;
        RECT 140.515 65.505 140.685 65.675 ;
        RECT 140.515 64.965 140.685 65.135 ;
        RECT 140.515 63.415 140.685 63.585 ;
        RECT 140.515 62.875 140.685 63.045 ;
        RECT 140.515 61.325 140.685 61.495 ;
        RECT 140.515 60.785 140.685 60.955 ;
        RECT 140.515 59.235 140.685 59.405 ;
        RECT 140.515 58.695 140.685 58.865 ;
        RECT 140.515 57.145 140.685 57.315 ;
        RECT 141.805 69.685 141.975 69.855 ;
        RECT 141.805 69.145 141.975 69.315 ;
        RECT 141.805 67.595 141.975 67.765 ;
        RECT 141.805 67.055 141.975 67.225 ;
        RECT 141.805 65.505 141.975 65.675 ;
        RECT 141.805 64.965 141.975 65.135 ;
        RECT 141.805 63.415 141.975 63.585 ;
        RECT 141.805 62.875 141.975 63.045 ;
        RECT 141.805 61.325 141.975 61.495 ;
        RECT 141.805 60.785 141.975 60.955 ;
        RECT 141.805 59.235 141.975 59.405 ;
        RECT 141.805 58.695 141.975 58.865 ;
        RECT 141.805 57.145 141.975 57.315 ;
        RECT 143.095 69.685 143.265 69.855 ;
        RECT 143.095 69.145 143.265 69.315 ;
        RECT 143.095 67.595 143.265 67.765 ;
        RECT 143.095 67.055 143.265 67.225 ;
        RECT 143.095 65.505 143.265 65.675 ;
        RECT 143.095 64.965 143.265 65.135 ;
        RECT 143.095 63.415 143.265 63.585 ;
        RECT 143.095 62.875 143.265 63.045 ;
        RECT 143.095 61.325 143.265 61.495 ;
        RECT 143.095 60.785 143.265 60.955 ;
        RECT 143.095 59.235 143.265 59.405 ;
        RECT 143.095 58.695 143.265 58.865 ;
        RECT 143.095 57.145 143.265 57.315 ;
        RECT 144.385 69.685 144.555 69.855 ;
        RECT 144.385 69.145 144.555 69.315 ;
        RECT 144.385 67.595 144.555 67.765 ;
        RECT 144.385 67.055 144.555 67.225 ;
        RECT 144.385 65.505 144.555 65.675 ;
        RECT 144.385 64.965 144.555 65.135 ;
        RECT 144.385 63.415 144.555 63.585 ;
        RECT 144.385 62.875 144.555 63.045 ;
        RECT 144.385 61.325 144.555 61.495 ;
        RECT 144.385 60.785 144.555 60.955 ;
        RECT 144.385 59.235 144.555 59.405 ;
        RECT 144.385 58.695 144.555 58.865 ;
        RECT 144.385 57.145 144.555 57.315 ;
        RECT 145.675 69.685 145.845 69.855 ;
        RECT 145.675 69.145 145.845 69.315 ;
        RECT 145.675 67.595 145.845 67.765 ;
        RECT 145.675 67.055 145.845 67.225 ;
        RECT 145.675 65.505 145.845 65.675 ;
        RECT 145.675 64.965 145.845 65.135 ;
        RECT 145.675 63.415 145.845 63.585 ;
        RECT 145.675 62.875 145.845 63.045 ;
        RECT 145.675 61.325 145.845 61.495 ;
        RECT 145.675 60.785 145.845 60.955 ;
        RECT 145.675 59.235 145.845 59.405 ;
        RECT 145.675 58.695 145.845 58.865 ;
        RECT 145.675 57.145 145.845 57.315 ;
        RECT 146.965 69.685 147.135 69.855 ;
        RECT 146.965 69.145 147.135 69.315 ;
        RECT 146.965 67.595 147.135 67.765 ;
        RECT 146.965 67.055 147.135 67.225 ;
        RECT 146.965 65.505 147.135 65.675 ;
        RECT 146.965 64.965 147.135 65.135 ;
        RECT 146.965 63.415 147.135 63.585 ;
        RECT 146.965 62.875 147.135 63.045 ;
        RECT 146.965 61.325 147.135 61.495 ;
        RECT 146.965 60.785 147.135 60.955 ;
        RECT 146.965 59.235 147.135 59.405 ;
        RECT 146.965 58.695 147.135 58.865 ;
        RECT 146.965 57.145 147.135 57.315 ;
        RECT 148.255 69.685 148.425 69.855 ;
        RECT 148.255 69.145 148.425 69.315 ;
        RECT 148.255 67.595 148.425 67.765 ;
        RECT 148.255 67.055 148.425 67.225 ;
        RECT 148.255 65.505 148.425 65.675 ;
        RECT 148.255 64.965 148.425 65.135 ;
        RECT 148.255 63.415 148.425 63.585 ;
        RECT 148.255 62.875 148.425 63.045 ;
        RECT 148.255 61.325 148.425 61.495 ;
        RECT 148.255 60.785 148.425 60.955 ;
        RECT 148.255 59.235 148.425 59.405 ;
        RECT 148.255 58.695 148.425 58.865 ;
        RECT 148.255 57.145 148.425 57.315 ;
        RECT 116.380 55.290 116.800 55.460 ;
        RECT 116.380 54.320 116.800 54.490 ;
        RECT 130.660 55.000 131.080 55.170 ;
        RECT 142.770 54.980 143.190 55.150 ;
        RECT 130.660 54.030 131.080 54.200 ;
        RECT 142.770 54.010 143.190 54.180 ;
        RECT 116.230 47.245 118.150 47.415 ;
        RECT 129.930 47.485 131.850 47.655 ;
        RECT 119.090 46.050 119.580 46.820 ;
        RECT 132.890 46.490 133.190 47.010 ;
        RECT 116.230 45.605 118.150 45.775 ;
        RECT 129.930 45.845 131.850 46.015 ;
        RECT 142.610 47.255 144.530 47.425 ;
        RECT 145.550 46.250 145.860 46.800 ;
        RECT 142.610 45.615 144.530 45.785 ;
        RECT 130.125 42.475 130.600 42.870 ;
        RECT 143.490 42.475 143.965 42.870 ;
        RECT 149.060 42.650 150.310 44.100 ;
        RECT 112.560 41.710 112.730 41.880 ;
        RECT 113.850 41.710 114.020 41.880 ;
        RECT 115.140 41.710 115.310 41.880 ;
        RECT 116.430 41.710 116.600 41.880 ;
        RECT 117.720 41.710 117.890 41.880 ;
        RECT 119.010 41.710 119.180 41.880 ;
        RECT 120.300 41.710 120.470 41.880 ;
        RECT 121.590 41.710 121.760 41.880 ;
        RECT 112.560 40.160 112.730 40.330 ;
        RECT 112.560 39.620 112.730 39.790 ;
        RECT 112.560 38.070 112.730 38.240 ;
        RECT 112.560 37.530 112.730 37.700 ;
        RECT 112.560 35.980 112.730 36.150 ;
        RECT 112.560 35.440 112.730 35.610 ;
        RECT 112.560 33.890 112.730 34.060 ;
        RECT 112.560 33.350 112.730 33.520 ;
        RECT 112.560 31.800 112.730 31.970 ;
        RECT 112.560 31.260 112.730 31.430 ;
        RECT 112.560 29.710 112.730 29.880 ;
        RECT 112.560 29.170 112.730 29.340 ;
        RECT 112.560 27.620 112.730 27.790 ;
        RECT 113.850 40.160 114.020 40.330 ;
        RECT 113.850 39.620 114.020 39.790 ;
        RECT 113.850 38.070 114.020 38.240 ;
        RECT 113.850 37.530 114.020 37.700 ;
        RECT 113.850 35.980 114.020 36.150 ;
        RECT 113.850 35.440 114.020 35.610 ;
        RECT 113.850 33.890 114.020 34.060 ;
        RECT 113.850 33.350 114.020 33.520 ;
        RECT 113.850 31.800 114.020 31.970 ;
        RECT 113.850 31.260 114.020 31.430 ;
        RECT 113.850 29.710 114.020 29.880 ;
        RECT 113.850 29.170 114.020 29.340 ;
        RECT 113.850 27.620 114.020 27.790 ;
        RECT 115.140 40.160 115.310 40.330 ;
        RECT 115.140 39.620 115.310 39.790 ;
        RECT 115.140 38.070 115.310 38.240 ;
        RECT 115.140 37.530 115.310 37.700 ;
        RECT 115.140 35.980 115.310 36.150 ;
        RECT 115.140 35.440 115.310 35.610 ;
        RECT 115.140 33.890 115.310 34.060 ;
        RECT 115.140 33.350 115.310 33.520 ;
        RECT 115.140 31.800 115.310 31.970 ;
        RECT 115.140 31.260 115.310 31.430 ;
        RECT 115.140 29.710 115.310 29.880 ;
        RECT 115.140 29.170 115.310 29.340 ;
        RECT 115.140 27.620 115.310 27.790 ;
        RECT 116.430 40.160 116.600 40.330 ;
        RECT 116.430 39.620 116.600 39.790 ;
        RECT 116.430 38.070 116.600 38.240 ;
        RECT 116.430 37.530 116.600 37.700 ;
        RECT 116.430 35.980 116.600 36.150 ;
        RECT 116.430 35.440 116.600 35.610 ;
        RECT 116.430 33.890 116.600 34.060 ;
        RECT 116.430 33.350 116.600 33.520 ;
        RECT 116.430 31.800 116.600 31.970 ;
        RECT 116.430 31.260 116.600 31.430 ;
        RECT 116.430 29.710 116.600 29.880 ;
        RECT 116.430 29.170 116.600 29.340 ;
        RECT 116.430 27.620 116.600 27.790 ;
        RECT 117.720 40.160 117.890 40.330 ;
        RECT 117.720 39.620 117.890 39.790 ;
        RECT 117.720 38.070 117.890 38.240 ;
        RECT 117.720 37.530 117.890 37.700 ;
        RECT 117.720 35.980 117.890 36.150 ;
        RECT 117.720 35.440 117.890 35.610 ;
        RECT 117.720 33.890 117.890 34.060 ;
        RECT 117.720 33.350 117.890 33.520 ;
        RECT 117.720 31.800 117.890 31.970 ;
        RECT 117.720 31.260 117.890 31.430 ;
        RECT 117.720 29.710 117.890 29.880 ;
        RECT 117.720 29.170 117.890 29.340 ;
        RECT 117.720 27.620 117.890 27.790 ;
        RECT 119.010 40.160 119.180 40.330 ;
        RECT 119.010 39.620 119.180 39.790 ;
        RECT 119.010 38.070 119.180 38.240 ;
        RECT 119.010 37.530 119.180 37.700 ;
        RECT 119.010 35.980 119.180 36.150 ;
        RECT 119.010 35.440 119.180 35.610 ;
        RECT 119.010 33.890 119.180 34.060 ;
        RECT 119.010 33.350 119.180 33.520 ;
        RECT 119.010 31.800 119.180 31.970 ;
        RECT 119.010 31.260 119.180 31.430 ;
        RECT 119.010 29.710 119.180 29.880 ;
        RECT 119.010 29.170 119.180 29.340 ;
        RECT 119.010 27.620 119.180 27.790 ;
        RECT 120.300 40.160 120.470 40.330 ;
        RECT 120.300 39.620 120.470 39.790 ;
        RECT 120.300 38.070 120.470 38.240 ;
        RECT 120.300 37.530 120.470 37.700 ;
        RECT 120.300 35.980 120.470 36.150 ;
        RECT 120.300 35.440 120.470 35.610 ;
        RECT 120.300 33.890 120.470 34.060 ;
        RECT 120.300 33.350 120.470 33.520 ;
        RECT 120.300 31.800 120.470 31.970 ;
        RECT 120.300 31.260 120.470 31.430 ;
        RECT 120.300 29.710 120.470 29.880 ;
        RECT 120.300 29.170 120.470 29.340 ;
        RECT 120.300 27.620 120.470 27.790 ;
        RECT 121.590 40.160 121.760 40.330 ;
        RECT 121.590 39.620 121.760 39.790 ;
        RECT 121.590 38.070 121.760 38.240 ;
        RECT 121.590 37.530 121.760 37.700 ;
        RECT 121.590 35.980 121.760 36.150 ;
        RECT 121.590 35.440 121.760 35.610 ;
        RECT 121.590 33.890 121.760 34.060 ;
        RECT 121.590 33.350 121.760 33.520 ;
        RECT 121.590 31.800 121.760 31.970 ;
        RECT 121.590 31.260 121.760 31.430 ;
        RECT 121.590 29.710 121.760 29.880 ;
        RECT 121.590 29.170 121.760 29.340 ;
        RECT 121.590 27.620 121.760 27.790 ;
        RECT 125.910 41.710 126.080 41.880 ;
        RECT 127.200 41.710 127.370 41.880 ;
        RECT 128.490 41.710 128.660 41.880 ;
        RECT 129.780 41.710 129.950 41.880 ;
        RECT 131.070 41.710 131.240 41.880 ;
        RECT 132.360 41.710 132.530 41.880 ;
        RECT 133.650 41.710 133.820 41.880 ;
        RECT 134.940 41.710 135.110 41.880 ;
        RECT 125.910 40.160 126.080 40.330 ;
        RECT 125.910 39.620 126.080 39.790 ;
        RECT 125.910 38.070 126.080 38.240 ;
        RECT 125.910 37.530 126.080 37.700 ;
        RECT 125.910 35.980 126.080 36.150 ;
        RECT 125.910 35.440 126.080 35.610 ;
        RECT 125.910 33.890 126.080 34.060 ;
        RECT 125.910 33.350 126.080 33.520 ;
        RECT 125.910 31.800 126.080 31.970 ;
        RECT 125.910 31.260 126.080 31.430 ;
        RECT 125.910 29.710 126.080 29.880 ;
        RECT 125.910 29.170 126.080 29.340 ;
        RECT 125.910 27.620 126.080 27.790 ;
        RECT 127.200 40.160 127.370 40.330 ;
        RECT 127.200 39.620 127.370 39.790 ;
        RECT 127.200 38.070 127.370 38.240 ;
        RECT 127.200 37.530 127.370 37.700 ;
        RECT 127.200 35.980 127.370 36.150 ;
        RECT 127.200 35.440 127.370 35.610 ;
        RECT 127.200 33.890 127.370 34.060 ;
        RECT 127.200 33.350 127.370 33.520 ;
        RECT 127.200 31.800 127.370 31.970 ;
        RECT 127.200 31.260 127.370 31.430 ;
        RECT 127.200 29.710 127.370 29.880 ;
        RECT 127.200 29.170 127.370 29.340 ;
        RECT 127.200 27.620 127.370 27.790 ;
        RECT 128.490 40.160 128.660 40.330 ;
        RECT 128.490 39.620 128.660 39.790 ;
        RECT 128.490 38.070 128.660 38.240 ;
        RECT 128.490 37.530 128.660 37.700 ;
        RECT 128.490 35.980 128.660 36.150 ;
        RECT 128.490 35.440 128.660 35.610 ;
        RECT 128.490 33.890 128.660 34.060 ;
        RECT 128.490 33.350 128.660 33.520 ;
        RECT 128.490 31.800 128.660 31.970 ;
        RECT 128.490 31.260 128.660 31.430 ;
        RECT 128.490 29.710 128.660 29.880 ;
        RECT 128.490 29.170 128.660 29.340 ;
        RECT 128.490 27.620 128.660 27.790 ;
        RECT 129.780 40.160 129.950 40.330 ;
        RECT 129.780 39.620 129.950 39.790 ;
        RECT 129.780 38.070 129.950 38.240 ;
        RECT 129.780 37.530 129.950 37.700 ;
        RECT 129.780 35.980 129.950 36.150 ;
        RECT 129.780 35.440 129.950 35.610 ;
        RECT 129.780 33.890 129.950 34.060 ;
        RECT 129.780 33.350 129.950 33.520 ;
        RECT 129.780 31.800 129.950 31.970 ;
        RECT 129.780 31.260 129.950 31.430 ;
        RECT 129.780 29.710 129.950 29.880 ;
        RECT 129.780 29.170 129.950 29.340 ;
        RECT 129.780 27.620 129.950 27.790 ;
        RECT 131.070 40.160 131.240 40.330 ;
        RECT 131.070 39.620 131.240 39.790 ;
        RECT 131.070 38.070 131.240 38.240 ;
        RECT 131.070 37.530 131.240 37.700 ;
        RECT 131.070 35.980 131.240 36.150 ;
        RECT 131.070 35.440 131.240 35.610 ;
        RECT 131.070 33.890 131.240 34.060 ;
        RECT 131.070 33.350 131.240 33.520 ;
        RECT 131.070 31.800 131.240 31.970 ;
        RECT 131.070 31.260 131.240 31.430 ;
        RECT 131.070 29.710 131.240 29.880 ;
        RECT 131.070 29.170 131.240 29.340 ;
        RECT 131.070 27.620 131.240 27.790 ;
        RECT 132.360 40.160 132.530 40.330 ;
        RECT 132.360 39.620 132.530 39.790 ;
        RECT 132.360 38.070 132.530 38.240 ;
        RECT 132.360 37.530 132.530 37.700 ;
        RECT 132.360 35.980 132.530 36.150 ;
        RECT 132.360 35.440 132.530 35.610 ;
        RECT 132.360 33.890 132.530 34.060 ;
        RECT 132.360 33.350 132.530 33.520 ;
        RECT 132.360 31.800 132.530 31.970 ;
        RECT 132.360 31.260 132.530 31.430 ;
        RECT 132.360 29.710 132.530 29.880 ;
        RECT 132.360 29.170 132.530 29.340 ;
        RECT 132.360 27.620 132.530 27.790 ;
        RECT 133.650 40.160 133.820 40.330 ;
        RECT 133.650 39.620 133.820 39.790 ;
        RECT 133.650 38.070 133.820 38.240 ;
        RECT 133.650 37.530 133.820 37.700 ;
        RECT 133.650 35.980 133.820 36.150 ;
        RECT 133.650 35.440 133.820 35.610 ;
        RECT 133.650 33.890 133.820 34.060 ;
        RECT 133.650 33.350 133.820 33.520 ;
        RECT 133.650 31.800 133.820 31.970 ;
        RECT 133.650 31.260 133.820 31.430 ;
        RECT 133.650 29.710 133.820 29.880 ;
        RECT 133.650 29.170 133.820 29.340 ;
        RECT 133.650 27.620 133.820 27.790 ;
        RECT 134.940 40.160 135.110 40.330 ;
        RECT 134.940 39.620 135.110 39.790 ;
        RECT 134.940 38.070 135.110 38.240 ;
        RECT 134.940 37.530 135.110 37.700 ;
        RECT 134.940 35.980 135.110 36.150 ;
        RECT 134.940 35.440 135.110 35.610 ;
        RECT 134.940 33.890 135.110 34.060 ;
        RECT 134.940 33.350 135.110 33.520 ;
        RECT 134.940 31.800 135.110 31.970 ;
        RECT 134.940 31.260 135.110 31.430 ;
        RECT 134.940 29.710 135.110 29.880 ;
        RECT 134.940 29.170 135.110 29.340 ;
        RECT 139.225 41.715 139.395 41.885 ;
        RECT 140.515 41.715 140.685 41.885 ;
        RECT 141.805 41.715 141.975 41.885 ;
        RECT 143.095 41.715 143.265 41.885 ;
        RECT 144.385 41.715 144.555 41.885 ;
        RECT 145.675 41.715 145.845 41.885 ;
        RECT 146.965 41.715 147.135 41.885 ;
        RECT 148.255 41.715 148.425 41.885 ;
        RECT 139.225 40.165 139.395 40.335 ;
        RECT 139.225 39.625 139.395 39.795 ;
        RECT 139.225 38.075 139.395 38.245 ;
        RECT 139.225 37.535 139.395 37.705 ;
        RECT 139.225 35.985 139.395 36.155 ;
        RECT 139.225 35.445 139.395 35.615 ;
        RECT 139.225 33.895 139.395 34.065 ;
        RECT 139.225 33.355 139.395 33.525 ;
        RECT 139.225 31.805 139.395 31.975 ;
        RECT 139.225 31.265 139.395 31.435 ;
        RECT 139.225 29.715 139.395 29.885 ;
        RECT 139.225 29.175 139.395 29.345 ;
        RECT 134.940 27.620 135.110 27.790 ;
        RECT 139.225 27.625 139.395 27.795 ;
        RECT 140.515 40.165 140.685 40.335 ;
        RECT 140.515 39.625 140.685 39.795 ;
        RECT 140.515 38.075 140.685 38.245 ;
        RECT 140.515 37.535 140.685 37.705 ;
        RECT 140.515 35.985 140.685 36.155 ;
        RECT 140.515 35.445 140.685 35.615 ;
        RECT 140.515 33.895 140.685 34.065 ;
        RECT 140.515 33.355 140.685 33.525 ;
        RECT 140.515 31.805 140.685 31.975 ;
        RECT 140.515 31.265 140.685 31.435 ;
        RECT 140.515 29.715 140.685 29.885 ;
        RECT 140.515 29.175 140.685 29.345 ;
        RECT 140.515 27.625 140.685 27.795 ;
        RECT 141.805 40.165 141.975 40.335 ;
        RECT 141.805 39.625 141.975 39.795 ;
        RECT 141.805 38.075 141.975 38.245 ;
        RECT 141.805 37.535 141.975 37.705 ;
        RECT 141.805 35.985 141.975 36.155 ;
        RECT 141.805 35.445 141.975 35.615 ;
        RECT 141.805 33.895 141.975 34.065 ;
        RECT 141.805 33.355 141.975 33.525 ;
        RECT 141.805 31.805 141.975 31.975 ;
        RECT 141.805 31.265 141.975 31.435 ;
        RECT 141.805 29.715 141.975 29.885 ;
        RECT 141.805 29.175 141.975 29.345 ;
        RECT 141.805 27.625 141.975 27.795 ;
        RECT 143.095 40.165 143.265 40.335 ;
        RECT 143.095 39.625 143.265 39.795 ;
        RECT 143.095 38.075 143.265 38.245 ;
        RECT 143.095 37.535 143.265 37.705 ;
        RECT 143.095 35.985 143.265 36.155 ;
        RECT 143.095 35.445 143.265 35.615 ;
        RECT 143.095 33.895 143.265 34.065 ;
        RECT 143.095 33.355 143.265 33.525 ;
        RECT 143.095 31.805 143.265 31.975 ;
        RECT 143.095 31.265 143.265 31.435 ;
        RECT 143.095 29.715 143.265 29.885 ;
        RECT 143.095 29.175 143.265 29.345 ;
        RECT 143.095 27.625 143.265 27.795 ;
        RECT 144.385 40.165 144.555 40.335 ;
        RECT 144.385 39.625 144.555 39.795 ;
        RECT 144.385 38.075 144.555 38.245 ;
        RECT 144.385 37.535 144.555 37.705 ;
        RECT 144.385 35.985 144.555 36.155 ;
        RECT 144.385 35.445 144.555 35.615 ;
        RECT 144.385 33.895 144.555 34.065 ;
        RECT 144.385 33.355 144.555 33.525 ;
        RECT 144.385 31.805 144.555 31.975 ;
        RECT 144.385 31.265 144.555 31.435 ;
        RECT 144.385 29.715 144.555 29.885 ;
        RECT 144.385 29.175 144.555 29.345 ;
        RECT 144.385 27.625 144.555 27.795 ;
        RECT 145.675 40.165 145.845 40.335 ;
        RECT 145.675 39.625 145.845 39.795 ;
        RECT 145.675 38.075 145.845 38.245 ;
        RECT 145.675 37.535 145.845 37.705 ;
        RECT 145.675 35.985 145.845 36.155 ;
        RECT 145.675 35.445 145.845 35.615 ;
        RECT 145.675 33.895 145.845 34.065 ;
        RECT 145.675 33.355 145.845 33.525 ;
        RECT 145.675 31.805 145.845 31.975 ;
        RECT 145.675 31.265 145.845 31.435 ;
        RECT 145.675 29.715 145.845 29.885 ;
        RECT 145.675 29.175 145.845 29.345 ;
        RECT 145.675 27.625 145.845 27.795 ;
        RECT 146.965 40.165 147.135 40.335 ;
        RECT 146.965 39.625 147.135 39.795 ;
        RECT 146.965 38.075 147.135 38.245 ;
        RECT 146.965 37.535 147.135 37.705 ;
        RECT 146.965 35.985 147.135 36.155 ;
        RECT 146.965 35.445 147.135 35.615 ;
        RECT 146.965 33.895 147.135 34.065 ;
        RECT 146.965 33.355 147.135 33.525 ;
        RECT 146.965 31.805 147.135 31.975 ;
        RECT 146.965 31.265 147.135 31.435 ;
        RECT 146.965 29.715 147.135 29.885 ;
        RECT 146.965 29.175 147.135 29.345 ;
        RECT 146.965 27.625 147.135 27.795 ;
        RECT 148.255 40.165 148.425 40.335 ;
        RECT 148.255 39.625 148.425 39.795 ;
        RECT 148.255 38.075 148.425 38.245 ;
        RECT 148.255 37.535 148.425 37.705 ;
        RECT 148.255 35.985 148.425 36.155 ;
        RECT 148.255 35.445 148.425 35.615 ;
        RECT 148.255 33.895 148.425 34.065 ;
        RECT 148.255 33.355 148.425 33.525 ;
        RECT 148.255 31.805 148.425 31.975 ;
        RECT 148.255 31.265 148.425 31.435 ;
        RECT 148.255 29.715 148.425 29.885 ;
        RECT 148.255 29.175 148.425 29.345 ;
        RECT 148.255 27.625 148.425 27.795 ;
        RECT 116.360 25.770 116.780 25.940 ;
        RECT 118.350 25.070 118.900 25.530 ;
        RECT 116.360 24.800 116.780 24.970 ;
        RECT 129.470 25.550 129.890 25.720 ;
        RECT 131.380 24.860 131.930 25.320 ;
        RECT 143.470 25.680 143.890 25.850 ;
        RECT 145.280 24.990 145.830 25.450 ;
        RECT 129.470 24.580 129.890 24.750 ;
        RECT 143.470 24.710 143.890 24.880 ;
        RECT 234.370 107.550 236.355 107.740 ;
        RECT 255.775 107.550 257.760 107.740 ;
        RECT 281.755 107.560 283.740 107.750 ;
        RECT 234.370 105.960 236.355 106.150 ;
        RECT 255.775 105.960 257.760 106.150 ;
        RECT 281.755 105.970 283.740 106.160 ;
        RECT 255.775 104.370 257.760 104.560 ;
        RECT 260.350 104.380 262.335 104.570 ;
        RECT 281.755 104.380 283.740 104.570 ;
        RECT 255.775 102.780 257.760 102.970 ;
        RECT 260.350 102.790 262.335 102.980 ;
        RECT 281.755 102.790 283.740 102.980 ;
        RECT 255.775 101.190 257.760 101.380 ;
        RECT 260.350 101.200 262.335 101.390 ;
        RECT 281.755 101.200 283.740 101.390 ;
        RECT 234.370 99.600 236.355 99.790 ;
        RECT 255.775 99.600 257.760 99.790 ;
        RECT 281.755 99.610 283.740 99.800 ;
        RECT 234.370 98.010 236.355 98.200 ;
        RECT 260.350 98.020 262.335 98.210 ;
        RECT 234.370 96.420 236.355 96.610 ;
        RECT 260.350 96.430 262.335 96.620 ;
        RECT 255.775 94.830 257.760 95.020 ;
        RECT 260.350 94.840 262.335 95.030 ;
        RECT 214.570 77.770 214.770 77.960 ;
        RECT 215.960 77.770 216.130 77.940 ;
        RECT 245.590 88.650 245.850 89.150 ;
        RECT 246.490 88.710 246.750 89.130 ;
        RECT 250.110 88.750 250.500 89.240 ;
        RECT 259.000 88.720 259.440 89.380 ;
        RECT 243.200 84.440 243.530 84.700 ;
        RECT 244.960 84.440 245.290 84.700 ;
        RECT 240.500 77.860 240.700 78.050 ;
        RECT 241.890 77.860 242.060 78.030 ;
        RECT 224.220 69.980 226.140 70.150 ;
        RECT 229.080 69.980 231.000 70.150 ;
        RECT 271.330 87.650 271.740 88.080 ;
        RECT 278.530 87.720 278.830 87.990 ;
        RECT 250.740 85.635 251.160 85.805 ;
        RECT 250.220 81.680 250.390 84.120 ;
        RECT 251.510 81.680 251.680 84.120 ;
        RECT 255.195 81.610 255.365 84.050 ;
        RECT 258.485 81.620 258.655 84.060 ;
        RECT 259.710 85.505 260.130 85.675 ;
        RECT 259.190 81.550 259.360 83.990 ;
        RECT 260.480 81.550 260.650 83.990 ;
        RECT 262.260 83.200 262.810 83.580 ;
        RECT 263.430 79.650 263.810 80.000 ;
        RECT 260.260 76.580 260.860 76.860 ;
        RECT 249.965 75.440 250.465 75.945 ;
        RECT 261.130 75.700 261.750 75.960 ;
        RECT 250.130 69.760 250.340 69.960 ;
        RECT 266.380 77.920 266.580 78.110 ;
        RECT 267.770 77.920 267.940 78.090 ;
        RECT 265.830 72.390 266.150 72.830 ;
        RECT 253.680 66.720 254.670 66.920 ;
        RECT 256.735 66.720 257.755 66.910 ;
        RECT 282.190 84.910 283.110 85.100 ;
        RECT 295.240 82.970 295.710 83.340 ;
        RECT 483.010 77.930 486.720 81.080 ;
        RECT 538.290 78.560 542.000 81.710 ;
        RECT 294.660 76.880 294.860 77.070 ;
        RECT 296.050 76.880 296.220 77.050 ;
        RECT 277.300 72.210 277.720 72.380 ;
        RECT 278.590 72.210 279.010 72.380 ;
        RECT 279.880 72.210 280.300 72.380 ;
        RECT 282.300 72.210 282.720 72.380 ;
        RECT 283.590 72.210 284.010 72.380 ;
        RECT 284.880 72.210 285.300 72.380 ;
        RECT 277.300 67.430 277.720 67.600 ;
        RECT 277.300 62.650 277.720 62.820 ;
        RECT 278.590 67.430 279.010 67.600 ;
        RECT 278.590 62.650 279.010 62.820 ;
        RECT 279.880 67.430 280.300 67.600 ;
        RECT 279.880 62.650 280.300 62.820 ;
        RECT 282.300 67.430 282.720 67.600 ;
        RECT 282.300 62.650 282.720 62.820 ;
        RECT 283.590 67.430 284.010 67.600 ;
        RECT 283.590 62.650 284.010 62.820 ;
        RECT 284.880 67.430 285.300 67.600 ;
        RECT 284.880 62.650 285.300 62.820 ;
        RECT 502.400 57.080 506.260 59.230 ;
        RECT 566.630 57.610 570.650 58.420 ;
        RECT 197.640 55.905 197.810 56.075 ;
        RECT 189.170 55.015 193.090 55.185 ;
        RECT 197.860 54.440 198.030 55.220 ;
        RECT 190.190 51.450 190.360 51.620 ;
        RECT 197.560 51.400 197.730 51.570 ;
        RECT 197.780 50.915 197.950 51.085 ;
        RECT 197.560 50.430 197.730 50.600 ;
        RECT 190.190 43.900 190.360 44.070 ;
        RECT 272.055 40.240 274.040 40.430 ;
        RECT 250.650 38.560 252.635 38.750 ;
        RECT 272.055 38.560 274.040 38.750 ;
        RECT 250.840 36.890 252.825 37.080 ;
        RECT 272.245 36.890 274.230 37.080 ;
        RECT 272.345 35.300 274.330 35.490 ;
        RECT 275.660 25.720 279.510 25.890 ;
        RECT 269.870 23.900 270.050 24.780 ;
        RECT 274.730 23.890 274.900 25.430 ;
        RECT 281.040 23.990 281.210 28.870 ;
        RECT 282.330 23.990 282.500 28.870 ;
        RECT 288.610 26.690 288.790 28.300 ;
        RECT 292.140 24.640 292.310 25.060 ;
        RECT 292.800 23.820 292.980 28.710 ;
        RECT 295.090 23.820 295.260 28.700 ;
        RECT 281.350 23.530 282.190 23.700 ;
        RECT 249.610 22.950 257.450 23.130 ;
        RECT 257.590 21.540 257.760 22.700 ;
        RECT 294.110 23.010 294.950 23.180 ;
        RECT 283.020 21.830 283.190 22.990 ;
        RECT 289.610 22.750 290.450 22.920 ;
        RECT 290.900 22.750 291.740 22.930 ;
        RECT 284.390 22.410 288.230 22.580 ;
        RECT 258.460 21.410 266.300 21.580 ;
        RECT 266.750 21.410 274.590 21.580 ;
        RECT 275.040 21.410 282.880 21.580 ;
        RECT 288.370 21.280 288.540 22.160 ;
        RECT 258.540 20.620 266.380 20.790 ;
        RECT 266.830 20.620 274.670 20.790 ;
        RECT 275.120 20.620 282.960 20.790 ;
        RECT 249.350 18.510 249.520 19.670 ;
        RECT 257.640 18.510 257.810 19.670 ;
        RECT 123.830 15.655 124.000 15.825 ;
        RECT 140.740 15.565 140.910 15.735 ;
        RECT 159.210 15.655 159.380 15.825 ;
        RECT 283.100 15.660 283.270 20.370 ;
        RECT 290.580 19.620 290.760 22.500 ;
        RECT 295.090 21.860 295.260 22.760 ;
        RECT 294.110 21.440 294.950 21.610 ;
        RECT 115.360 14.765 119.280 14.935 ;
        RECT 132.270 14.675 136.190 14.845 ;
        RECT 140.960 14.100 141.130 14.880 ;
        RECT 150.740 14.765 154.660 14.935 ;
        RECT 159.430 14.190 159.600 14.970 ;
        RECT 275.120 14.350 282.960 14.530 ;
        RECT 283.100 12.720 283.270 14.100 ;
        RECT 116.380 11.200 116.550 11.370 ;
        RECT 123.750 11.150 123.920 11.320 ;
        RECT 133.290 11.110 133.460 11.280 ;
        RECT 140.660 11.060 140.830 11.230 ;
        RECT 151.760 11.200 151.930 11.370 ;
        RECT 159.130 11.150 159.300 11.320 ;
        RECT 140.880 10.575 141.050 10.745 ;
        RECT 159.350 10.665 159.520 10.835 ;
        RECT 123.750 10.180 123.920 10.350 ;
        RECT 140.660 10.090 140.830 10.260 ;
        RECT 159.130 10.180 159.300 10.350 ;
        RECT 116.380 3.650 116.550 3.820 ;
        RECT 133.290 3.560 133.460 3.730 ;
        RECT 151.760 3.650 151.930 3.820 ;
      LAYER met1 ;
        RECT 46.790 330.925 54.750 331.155 ;
        RECT 55.080 330.925 63.040 331.155 ;
        RECT 72.790 330.925 80.750 331.155 ;
        RECT 81.080 330.925 89.040 331.155 ;
        RECT 98.790 330.925 106.750 331.155 ;
        RECT 107.080 330.925 115.040 331.155 ;
        RECT 124.790 330.925 132.750 331.155 ;
        RECT 133.080 330.925 141.040 331.155 ;
        RECT 150.790 330.925 158.750 331.155 ;
        RECT 159.080 330.925 167.040 331.155 ;
        RECT 176.790 330.925 184.750 331.155 ;
        RECT 185.080 330.925 193.040 331.155 ;
        RECT 202.790 330.925 210.750 331.155 ;
        RECT 211.080 330.925 219.040 331.155 ;
        RECT 228.790 330.925 236.750 331.155 ;
        RECT 237.080 330.925 245.040 331.155 ;
        RECT 254.790 330.925 262.750 331.155 ;
        RECT 263.080 330.925 271.040 331.155 ;
        RECT 280.790 330.925 288.750 331.155 ;
        RECT 289.080 330.925 297.040 331.155 ;
        RECT 46.890 323.515 54.680 323.530 ;
        RECT 55.190 323.515 62.980 323.570 ;
        RECT 72.890 323.515 80.680 323.530 ;
        RECT 81.190 323.515 88.980 323.570 ;
        RECT 98.890 323.515 106.680 323.530 ;
        RECT 107.190 323.515 114.980 323.570 ;
        RECT 124.890 323.515 132.680 323.530 ;
        RECT 133.190 323.515 140.980 323.570 ;
        RECT 150.890 323.515 158.680 323.530 ;
        RECT 159.190 323.515 166.980 323.570 ;
        RECT 176.890 323.515 184.680 323.530 ;
        RECT 185.190 323.515 192.980 323.570 ;
        RECT 202.890 323.515 210.680 323.530 ;
        RECT 211.190 323.515 218.980 323.570 ;
        RECT 228.890 323.515 236.680 323.530 ;
        RECT 237.190 323.515 244.980 323.570 ;
        RECT 254.890 323.515 262.680 323.530 ;
        RECT 263.190 323.515 270.980 323.570 ;
        RECT 280.890 323.515 288.680 323.530 ;
        RECT 289.190 323.515 296.980 323.570 ;
        RECT 46.790 323.285 54.750 323.515 ;
        RECT 55.080 323.285 63.040 323.515 ;
        RECT 72.790 323.285 80.750 323.515 ;
        RECT 81.080 323.285 89.040 323.515 ;
        RECT 98.790 323.285 106.750 323.515 ;
        RECT 107.080 323.285 115.040 323.515 ;
        RECT 124.790 323.285 132.750 323.515 ;
        RECT 133.080 323.285 141.040 323.515 ;
        RECT 150.790 323.285 158.750 323.515 ;
        RECT 159.080 323.285 167.040 323.515 ;
        RECT 176.790 323.285 184.750 323.515 ;
        RECT 185.080 323.285 193.040 323.515 ;
        RECT 202.790 323.285 210.750 323.515 ;
        RECT 211.080 323.285 219.040 323.515 ;
        RECT 228.790 323.285 236.750 323.515 ;
        RECT 237.080 323.285 245.040 323.515 ;
        RECT 254.790 323.285 262.750 323.515 ;
        RECT 263.080 323.285 271.040 323.515 ;
        RECT 280.790 323.285 288.750 323.515 ;
        RECT 289.080 323.285 297.040 323.515 ;
        RECT 46.890 322.975 54.680 323.285 ;
        RECT 55.190 322.975 62.980 323.285 ;
        RECT 72.890 322.975 80.680 323.285 ;
        RECT 81.190 322.975 88.980 323.285 ;
        RECT 98.890 322.975 106.680 323.285 ;
        RECT 107.190 322.975 114.980 323.285 ;
        RECT 124.890 322.975 132.680 323.285 ;
        RECT 133.190 322.975 140.980 323.285 ;
        RECT 150.890 322.975 158.680 323.285 ;
        RECT 159.190 322.975 166.980 323.285 ;
        RECT 176.890 322.975 184.680 323.285 ;
        RECT 185.190 322.975 192.980 323.285 ;
        RECT 202.890 322.975 210.680 323.285 ;
        RECT 211.190 322.975 218.980 323.285 ;
        RECT 228.890 322.975 236.680 323.285 ;
        RECT 237.190 322.975 244.980 323.285 ;
        RECT 254.890 322.975 262.680 323.285 ;
        RECT 263.190 322.975 270.980 323.285 ;
        RECT 280.890 322.975 288.680 323.285 ;
        RECT 289.190 322.975 296.980 323.285 ;
        RECT 46.790 322.745 54.750 322.975 ;
        RECT 55.080 322.745 63.040 322.975 ;
        RECT 72.790 322.745 80.750 322.975 ;
        RECT 81.080 322.745 89.040 322.975 ;
        RECT 98.790 322.745 106.750 322.975 ;
        RECT 107.080 322.745 115.040 322.975 ;
        RECT 124.790 322.745 132.750 322.975 ;
        RECT 133.080 322.745 141.040 322.975 ;
        RECT 150.790 322.745 158.750 322.975 ;
        RECT 159.080 322.745 167.040 322.975 ;
        RECT 176.790 322.745 184.750 322.975 ;
        RECT 185.080 322.745 193.040 322.975 ;
        RECT 202.790 322.745 210.750 322.975 ;
        RECT 211.080 322.745 219.040 322.975 ;
        RECT 228.790 322.745 236.750 322.975 ;
        RECT 237.080 322.745 245.040 322.975 ;
        RECT 254.790 322.745 262.750 322.975 ;
        RECT 263.080 322.745 271.040 322.975 ;
        RECT 280.790 322.745 288.750 322.975 ;
        RECT 289.080 322.745 297.040 322.975 ;
        RECT 46.890 322.740 54.680 322.745 ;
        RECT 72.890 322.740 80.680 322.745 ;
        RECT 98.890 322.740 106.680 322.745 ;
        RECT 124.890 322.740 132.680 322.745 ;
        RECT 150.890 322.740 158.680 322.745 ;
        RECT 176.890 322.740 184.680 322.745 ;
        RECT 202.890 322.740 210.680 322.745 ;
        RECT 228.890 322.740 236.680 322.745 ;
        RECT 254.890 322.740 262.680 322.745 ;
        RECT 280.890 322.740 288.680 322.745 ;
        RECT 47.010 315.335 54.800 315.350 ;
        RECT 55.230 315.335 63.020 315.390 ;
        RECT 73.010 315.335 80.800 315.350 ;
        RECT 81.230 315.335 89.020 315.390 ;
        RECT 99.010 315.335 106.800 315.350 ;
        RECT 107.230 315.335 115.020 315.390 ;
        RECT 125.010 315.335 132.800 315.350 ;
        RECT 133.230 315.335 141.020 315.390 ;
        RECT 151.010 315.335 158.800 315.350 ;
        RECT 159.230 315.335 167.020 315.390 ;
        RECT 177.010 315.335 184.800 315.350 ;
        RECT 185.230 315.335 193.020 315.390 ;
        RECT 203.010 315.335 210.800 315.350 ;
        RECT 211.230 315.335 219.020 315.390 ;
        RECT 229.010 315.335 236.800 315.350 ;
        RECT 237.230 315.335 245.020 315.390 ;
        RECT 255.010 315.335 262.800 315.350 ;
        RECT 263.230 315.335 271.020 315.390 ;
        RECT 281.010 315.335 288.800 315.350 ;
        RECT 289.230 315.335 297.020 315.390 ;
        RECT 46.790 315.105 54.800 315.335 ;
        RECT 55.080 315.105 63.040 315.335 ;
        RECT 72.790 315.105 80.800 315.335 ;
        RECT 81.080 315.105 89.040 315.335 ;
        RECT 98.790 315.105 106.800 315.335 ;
        RECT 107.080 315.105 115.040 315.335 ;
        RECT 124.790 315.105 132.800 315.335 ;
        RECT 133.080 315.105 141.040 315.335 ;
        RECT 150.790 315.105 158.800 315.335 ;
        RECT 159.080 315.105 167.040 315.335 ;
        RECT 176.790 315.105 184.800 315.335 ;
        RECT 185.080 315.105 193.040 315.335 ;
        RECT 202.790 315.105 210.800 315.335 ;
        RECT 211.080 315.105 219.040 315.335 ;
        RECT 228.790 315.105 236.800 315.335 ;
        RECT 237.080 315.105 245.040 315.335 ;
        RECT 254.790 315.105 262.800 315.335 ;
        RECT 263.080 315.105 271.040 315.335 ;
        RECT 280.790 315.105 288.800 315.335 ;
        RECT 289.080 315.105 297.040 315.335 ;
        RECT 47.010 314.795 54.800 315.105 ;
        RECT 55.230 314.795 63.020 315.105 ;
        RECT 73.010 314.795 80.800 315.105 ;
        RECT 81.230 314.795 89.020 315.105 ;
        RECT 99.010 314.795 106.800 315.105 ;
        RECT 107.230 314.795 115.020 315.105 ;
        RECT 125.010 314.795 132.800 315.105 ;
        RECT 133.230 314.795 141.020 315.105 ;
        RECT 151.010 314.795 158.800 315.105 ;
        RECT 159.230 314.795 167.020 315.105 ;
        RECT 177.010 314.795 184.800 315.105 ;
        RECT 185.230 314.795 193.020 315.105 ;
        RECT 203.010 314.795 210.800 315.105 ;
        RECT 211.230 314.795 219.020 315.105 ;
        RECT 229.010 314.795 236.800 315.105 ;
        RECT 237.230 314.795 245.020 315.105 ;
        RECT 255.010 314.795 262.800 315.105 ;
        RECT 263.230 314.795 271.020 315.105 ;
        RECT 281.010 314.795 288.800 315.105 ;
        RECT 289.230 314.795 297.020 315.105 ;
        RECT 46.790 314.565 54.800 314.795 ;
        RECT 55.080 314.565 63.040 314.795 ;
        RECT 72.790 314.565 80.800 314.795 ;
        RECT 81.080 314.565 89.040 314.795 ;
        RECT 98.790 314.565 106.800 314.795 ;
        RECT 107.080 314.565 115.040 314.795 ;
        RECT 124.790 314.565 132.800 314.795 ;
        RECT 133.080 314.565 141.040 314.795 ;
        RECT 150.790 314.565 158.800 314.795 ;
        RECT 159.080 314.565 167.040 314.795 ;
        RECT 176.790 314.565 184.800 314.795 ;
        RECT 185.080 314.565 193.040 314.795 ;
        RECT 202.790 314.565 210.800 314.795 ;
        RECT 211.080 314.565 219.040 314.795 ;
        RECT 228.790 314.565 236.800 314.795 ;
        RECT 237.080 314.565 245.040 314.795 ;
        RECT 254.790 314.565 262.800 314.795 ;
        RECT 263.080 314.565 271.040 314.795 ;
        RECT 280.790 314.565 288.800 314.795 ;
        RECT 289.080 314.565 297.040 314.795 ;
        RECT 47.010 314.560 54.800 314.565 ;
        RECT 73.010 314.560 80.800 314.565 ;
        RECT 99.010 314.560 106.800 314.565 ;
        RECT 125.010 314.560 132.800 314.565 ;
        RECT 151.010 314.560 158.800 314.565 ;
        RECT 177.010 314.560 184.800 314.565 ;
        RECT 203.010 314.560 210.800 314.565 ;
        RECT 229.010 314.560 236.800 314.565 ;
        RECT 255.010 314.560 262.800 314.565 ;
        RECT 281.010 314.560 288.800 314.565 ;
        RECT 46.930 307.155 54.720 307.170 ;
        RECT 55.110 307.155 62.900 307.170 ;
        RECT 72.930 307.155 80.720 307.170 ;
        RECT 81.110 307.155 88.900 307.170 ;
        RECT 98.930 307.155 106.720 307.170 ;
        RECT 107.110 307.155 114.900 307.170 ;
        RECT 124.930 307.155 132.720 307.170 ;
        RECT 133.110 307.155 140.900 307.170 ;
        RECT 150.930 307.155 158.720 307.170 ;
        RECT 159.110 307.155 166.900 307.170 ;
        RECT 176.930 307.155 184.720 307.170 ;
        RECT 185.110 307.155 192.900 307.170 ;
        RECT 202.930 307.155 210.720 307.170 ;
        RECT 211.110 307.155 218.900 307.170 ;
        RECT 228.930 307.155 236.720 307.170 ;
        RECT 237.110 307.155 244.900 307.170 ;
        RECT 254.930 307.155 262.720 307.170 ;
        RECT 263.110 307.155 270.900 307.170 ;
        RECT 280.930 307.155 288.720 307.170 ;
        RECT 289.110 307.155 296.900 307.170 ;
        RECT 46.790 306.925 54.750 307.155 ;
        RECT 55.080 306.925 63.040 307.155 ;
        RECT 72.790 306.925 80.750 307.155 ;
        RECT 81.080 306.925 89.040 307.155 ;
        RECT 98.790 306.925 106.750 307.155 ;
        RECT 107.080 306.925 115.040 307.155 ;
        RECT 124.790 306.925 132.750 307.155 ;
        RECT 133.080 306.925 141.040 307.155 ;
        RECT 150.790 306.925 158.750 307.155 ;
        RECT 159.080 306.925 167.040 307.155 ;
        RECT 176.790 306.925 184.750 307.155 ;
        RECT 185.080 306.925 193.040 307.155 ;
        RECT 202.790 306.925 210.750 307.155 ;
        RECT 211.080 306.925 219.040 307.155 ;
        RECT 228.790 306.925 236.750 307.155 ;
        RECT 237.080 306.925 245.040 307.155 ;
        RECT 254.790 306.925 262.750 307.155 ;
        RECT 263.080 306.925 271.040 307.155 ;
        RECT 280.790 306.925 288.750 307.155 ;
        RECT 289.080 306.925 297.040 307.155 ;
        RECT 46.930 306.615 54.720 306.925 ;
        RECT 55.110 306.615 62.900 306.925 ;
        RECT 72.930 306.615 80.720 306.925 ;
        RECT 81.110 306.615 88.900 306.925 ;
        RECT 98.930 306.615 106.720 306.925 ;
        RECT 107.110 306.615 114.900 306.925 ;
        RECT 124.930 306.615 132.720 306.925 ;
        RECT 133.110 306.615 140.900 306.925 ;
        RECT 150.930 306.615 158.720 306.925 ;
        RECT 159.110 306.615 166.900 306.925 ;
        RECT 176.930 306.615 184.720 306.925 ;
        RECT 185.110 306.615 192.900 306.925 ;
        RECT 202.930 306.615 210.720 306.925 ;
        RECT 211.110 306.615 218.900 306.925 ;
        RECT 228.930 306.615 236.720 306.925 ;
        RECT 237.110 306.615 244.900 306.925 ;
        RECT 254.930 306.615 262.720 306.925 ;
        RECT 263.110 306.615 270.900 306.925 ;
        RECT 280.930 306.615 288.720 306.925 ;
        RECT 289.110 306.615 296.900 306.925 ;
        RECT 46.790 306.385 54.750 306.615 ;
        RECT 55.080 306.385 63.040 306.615 ;
        RECT 72.790 306.385 80.750 306.615 ;
        RECT 81.080 306.385 89.040 306.615 ;
        RECT 98.790 306.385 106.750 306.615 ;
        RECT 107.080 306.385 115.040 306.615 ;
        RECT 124.790 306.385 132.750 306.615 ;
        RECT 133.080 306.385 141.040 306.615 ;
        RECT 150.790 306.385 158.750 306.615 ;
        RECT 159.080 306.385 167.040 306.615 ;
        RECT 176.790 306.385 184.750 306.615 ;
        RECT 185.080 306.385 193.040 306.615 ;
        RECT 202.790 306.385 210.750 306.615 ;
        RECT 211.080 306.385 219.040 306.615 ;
        RECT 228.790 306.385 236.750 306.615 ;
        RECT 237.080 306.385 245.040 306.615 ;
        RECT 254.790 306.385 262.750 306.615 ;
        RECT 263.080 306.385 271.040 306.615 ;
        RECT 280.790 306.385 288.750 306.615 ;
        RECT 289.080 306.385 297.040 306.615 ;
        RECT 46.930 306.380 54.720 306.385 ;
        RECT 55.110 306.380 62.900 306.385 ;
        RECT 72.930 306.380 80.720 306.385 ;
        RECT 81.110 306.380 88.900 306.385 ;
        RECT 98.930 306.380 106.720 306.385 ;
        RECT 107.110 306.380 114.900 306.385 ;
        RECT 124.930 306.380 132.720 306.385 ;
        RECT 133.110 306.380 140.900 306.385 ;
        RECT 150.930 306.380 158.720 306.385 ;
        RECT 159.110 306.380 166.900 306.385 ;
        RECT 176.930 306.380 184.720 306.385 ;
        RECT 185.110 306.380 192.900 306.385 ;
        RECT 202.930 306.380 210.720 306.385 ;
        RECT 211.110 306.380 218.900 306.385 ;
        RECT 228.930 306.380 236.720 306.385 ;
        RECT 237.110 306.380 244.900 306.385 ;
        RECT 254.930 306.380 262.720 306.385 ;
        RECT 263.110 306.380 270.900 306.385 ;
        RECT 280.930 306.380 288.720 306.385 ;
        RECT 289.110 306.380 296.900 306.385 ;
        RECT 46.890 298.975 54.680 299.030 ;
        RECT 55.190 298.975 62.980 299.030 ;
        RECT 72.890 298.975 80.680 299.030 ;
        RECT 81.190 298.975 88.980 299.030 ;
        RECT 98.890 298.975 106.680 299.030 ;
        RECT 107.190 298.975 114.980 299.030 ;
        RECT 124.890 298.975 132.680 299.030 ;
        RECT 133.190 298.975 140.980 299.030 ;
        RECT 150.890 298.975 158.680 299.030 ;
        RECT 159.190 298.975 166.980 299.030 ;
        RECT 176.890 298.975 184.680 299.030 ;
        RECT 185.190 298.975 192.980 299.030 ;
        RECT 202.890 298.975 210.680 299.030 ;
        RECT 211.190 298.975 218.980 299.030 ;
        RECT 228.890 298.975 236.680 299.030 ;
        RECT 237.190 298.975 244.980 299.030 ;
        RECT 254.890 298.975 262.680 299.030 ;
        RECT 263.190 298.975 270.980 299.030 ;
        RECT 280.890 298.975 288.680 299.030 ;
        RECT 289.190 298.975 296.980 299.030 ;
        RECT 46.790 298.745 54.750 298.975 ;
        RECT 55.080 298.745 63.040 298.975 ;
        RECT 72.790 298.745 80.750 298.975 ;
        RECT 81.080 298.745 89.040 298.975 ;
        RECT 98.790 298.745 106.750 298.975 ;
        RECT 107.080 298.745 115.040 298.975 ;
        RECT 124.790 298.745 132.750 298.975 ;
        RECT 133.080 298.745 141.040 298.975 ;
        RECT 150.790 298.745 158.750 298.975 ;
        RECT 159.080 298.745 167.040 298.975 ;
        RECT 176.790 298.745 184.750 298.975 ;
        RECT 185.080 298.745 193.040 298.975 ;
        RECT 202.790 298.745 210.750 298.975 ;
        RECT 211.080 298.745 219.040 298.975 ;
        RECT 228.790 298.745 236.750 298.975 ;
        RECT 237.080 298.745 245.040 298.975 ;
        RECT 254.790 298.745 262.750 298.975 ;
        RECT 263.080 298.745 271.040 298.975 ;
        RECT 280.790 298.745 288.750 298.975 ;
        RECT 289.080 298.745 297.040 298.975 ;
        RECT 46.890 298.435 54.680 298.745 ;
        RECT 55.190 298.435 62.980 298.745 ;
        RECT 72.890 298.435 80.680 298.745 ;
        RECT 81.190 298.435 88.980 298.745 ;
        RECT 98.890 298.435 106.680 298.745 ;
        RECT 107.190 298.435 114.980 298.745 ;
        RECT 124.890 298.435 132.680 298.745 ;
        RECT 133.190 298.435 140.980 298.745 ;
        RECT 150.890 298.435 158.680 298.745 ;
        RECT 159.190 298.435 166.980 298.745 ;
        RECT 176.890 298.435 184.680 298.745 ;
        RECT 185.190 298.435 192.980 298.745 ;
        RECT 202.890 298.435 210.680 298.745 ;
        RECT 211.190 298.435 218.980 298.745 ;
        RECT 228.890 298.435 236.680 298.745 ;
        RECT 237.190 298.435 244.980 298.745 ;
        RECT 254.890 298.435 262.680 298.745 ;
        RECT 263.190 298.435 270.980 298.745 ;
        RECT 280.890 298.435 288.680 298.745 ;
        RECT 289.190 298.435 296.980 298.745 ;
        RECT 46.790 298.205 54.750 298.435 ;
        RECT 55.080 298.205 63.040 298.435 ;
        RECT 72.790 298.205 80.750 298.435 ;
        RECT 81.080 298.205 89.040 298.435 ;
        RECT 98.790 298.205 106.750 298.435 ;
        RECT 107.080 298.205 115.040 298.435 ;
        RECT 124.790 298.205 132.750 298.435 ;
        RECT 133.080 298.205 141.040 298.435 ;
        RECT 150.790 298.205 158.750 298.435 ;
        RECT 159.080 298.205 167.040 298.435 ;
        RECT 176.790 298.205 184.750 298.435 ;
        RECT 185.080 298.205 193.040 298.435 ;
        RECT 202.790 298.205 210.750 298.435 ;
        RECT 211.080 298.205 219.040 298.435 ;
        RECT 228.790 298.205 236.750 298.435 ;
        RECT 237.080 298.205 245.040 298.435 ;
        RECT 254.790 298.205 262.750 298.435 ;
        RECT 263.080 298.205 271.040 298.435 ;
        RECT 280.790 298.205 288.750 298.435 ;
        RECT 289.080 298.205 297.040 298.435 ;
        RECT 46.850 290.795 54.640 290.850 ;
        RECT 55.070 290.795 62.860 290.810 ;
        RECT 72.850 290.795 80.640 290.850 ;
        RECT 81.070 290.795 88.860 290.810 ;
        RECT 98.850 290.795 106.640 290.850 ;
        RECT 107.070 290.795 114.860 290.810 ;
        RECT 124.850 290.795 132.640 290.850 ;
        RECT 133.070 290.795 140.860 290.810 ;
        RECT 150.850 290.795 158.640 290.850 ;
        RECT 159.070 290.795 166.860 290.810 ;
        RECT 176.850 290.795 184.640 290.850 ;
        RECT 185.070 290.795 192.860 290.810 ;
        RECT 202.850 290.795 210.640 290.850 ;
        RECT 211.070 290.795 218.860 290.810 ;
        RECT 228.850 290.795 236.640 290.850 ;
        RECT 237.070 290.795 244.860 290.810 ;
        RECT 254.850 290.795 262.640 290.850 ;
        RECT 263.070 290.795 270.860 290.810 ;
        RECT 280.850 290.795 288.640 290.850 ;
        RECT 289.070 290.795 296.860 290.810 ;
        RECT 46.790 290.565 54.750 290.795 ;
        RECT 55.070 290.565 63.040 290.795 ;
        RECT 72.790 290.565 80.750 290.795 ;
        RECT 81.070 290.565 89.040 290.795 ;
        RECT 98.790 290.565 106.750 290.795 ;
        RECT 107.070 290.565 115.040 290.795 ;
        RECT 124.790 290.565 132.750 290.795 ;
        RECT 133.070 290.565 141.040 290.795 ;
        RECT 150.790 290.565 158.750 290.795 ;
        RECT 159.070 290.565 167.040 290.795 ;
        RECT 176.790 290.565 184.750 290.795 ;
        RECT 185.070 290.565 193.040 290.795 ;
        RECT 202.790 290.565 210.750 290.795 ;
        RECT 211.070 290.565 219.040 290.795 ;
        RECT 228.790 290.565 236.750 290.795 ;
        RECT 237.070 290.565 245.040 290.795 ;
        RECT 254.790 290.565 262.750 290.795 ;
        RECT 263.070 290.565 271.040 290.795 ;
        RECT 280.790 290.565 288.750 290.795 ;
        RECT 289.070 290.565 297.040 290.795 ;
        RECT 46.850 290.255 54.640 290.565 ;
        RECT 55.070 290.255 62.860 290.565 ;
        RECT 72.850 290.255 80.640 290.565 ;
        RECT 81.070 290.255 88.860 290.565 ;
        RECT 98.850 290.255 106.640 290.565 ;
        RECT 107.070 290.255 114.860 290.565 ;
        RECT 124.850 290.255 132.640 290.565 ;
        RECT 133.070 290.255 140.860 290.565 ;
        RECT 150.850 290.255 158.640 290.565 ;
        RECT 159.070 290.255 166.860 290.565 ;
        RECT 176.850 290.255 184.640 290.565 ;
        RECT 185.070 290.255 192.860 290.565 ;
        RECT 202.850 290.255 210.640 290.565 ;
        RECT 211.070 290.255 218.860 290.565 ;
        RECT 228.850 290.255 236.640 290.565 ;
        RECT 237.070 290.255 244.860 290.565 ;
        RECT 254.850 290.255 262.640 290.565 ;
        RECT 263.070 290.255 270.860 290.565 ;
        RECT 280.850 290.255 288.640 290.565 ;
        RECT 289.070 290.255 296.860 290.565 ;
        RECT 46.790 290.025 54.750 290.255 ;
        RECT 55.070 290.025 63.040 290.255 ;
        RECT 72.790 290.025 80.750 290.255 ;
        RECT 81.070 290.025 89.040 290.255 ;
        RECT 98.790 290.025 106.750 290.255 ;
        RECT 107.070 290.025 115.040 290.255 ;
        RECT 124.790 290.025 132.750 290.255 ;
        RECT 133.070 290.025 141.040 290.255 ;
        RECT 150.790 290.025 158.750 290.255 ;
        RECT 159.070 290.025 167.040 290.255 ;
        RECT 176.790 290.025 184.750 290.255 ;
        RECT 185.070 290.025 193.040 290.255 ;
        RECT 202.790 290.025 210.750 290.255 ;
        RECT 211.070 290.025 219.040 290.255 ;
        RECT 228.790 290.025 236.750 290.255 ;
        RECT 237.070 290.025 245.040 290.255 ;
        RECT 254.790 290.025 262.750 290.255 ;
        RECT 263.070 290.025 271.040 290.255 ;
        RECT 280.790 290.025 288.750 290.255 ;
        RECT 289.070 290.025 297.040 290.255 ;
        RECT 55.070 290.020 62.860 290.025 ;
        RECT 81.070 290.020 88.860 290.025 ;
        RECT 107.070 290.020 114.860 290.025 ;
        RECT 133.070 290.020 140.860 290.025 ;
        RECT 159.070 290.020 166.860 290.025 ;
        RECT 185.070 290.020 192.860 290.025 ;
        RECT 211.070 290.020 218.860 290.025 ;
        RECT 237.070 290.020 244.860 290.025 ;
        RECT 263.070 290.020 270.860 290.025 ;
        RECT 289.070 290.020 296.860 290.025 ;
        RECT 46.970 282.615 54.760 282.670 ;
        RECT 55.110 282.615 62.900 282.670 ;
        RECT 72.970 282.615 80.760 282.670 ;
        RECT 81.110 282.615 88.900 282.670 ;
        RECT 98.970 282.615 106.760 282.670 ;
        RECT 107.110 282.615 114.900 282.670 ;
        RECT 124.970 282.615 132.760 282.670 ;
        RECT 133.110 282.615 140.900 282.670 ;
        RECT 150.970 282.615 158.760 282.670 ;
        RECT 159.110 282.615 166.900 282.670 ;
        RECT 176.970 282.615 184.760 282.670 ;
        RECT 185.110 282.615 192.900 282.670 ;
        RECT 202.970 282.615 210.760 282.670 ;
        RECT 211.110 282.615 218.900 282.670 ;
        RECT 228.970 282.615 236.760 282.670 ;
        RECT 237.110 282.615 244.900 282.670 ;
        RECT 254.970 282.615 262.760 282.670 ;
        RECT 263.110 282.615 270.900 282.670 ;
        RECT 280.970 282.615 288.760 282.670 ;
        RECT 289.110 282.615 296.900 282.670 ;
        RECT 46.790 282.385 54.760 282.615 ;
        RECT 55.080 282.385 63.040 282.615 ;
        RECT 72.790 282.385 80.760 282.615 ;
        RECT 81.080 282.385 89.040 282.615 ;
        RECT 98.790 282.385 106.760 282.615 ;
        RECT 107.080 282.385 115.040 282.615 ;
        RECT 124.790 282.385 132.760 282.615 ;
        RECT 133.080 282.385 141.040 282.615 ;
        RECT 150.790 282.385 158.760 282.615 ;
        RECT 159.080 282.385 167.040 282.615 ;
        RECT 176.790 282.385 184.760 282.615 ;
        RECT 185.080 282.385 193.040 282.615 ;
        RECT 202.790 282.385 210.760 282.615 ;
        RECT 211.080 282.385 219.040 282.615 ;
        RECT 228.790 282.385 236.760 282.615 ;
        RECT 237.080 282.385 245.040 282.615 ;
        RECT 254.790 282.385 262.760 282.615 ;
        RECT 263.080 282.385 271.040 282.615 ;
        RECT 280.790 282.385 288.760 282.615 ;
        RECT 289.080 282.385 297.040 282.615 ;
        RECT 46.970 282.075 54.760 282.385 ;
        RECT 55.110 282.075 62.900 282.385 ;
        RECT 72.970 282.075 80.760 282.385 ;
        RECT 81.110 282.075 88.900 282.385 ;
        RECT 98.970 282.075 106.760 282.385 ;
        RECT 107.110 282.075 114.900 282.385 ;
        RECT 124.970 282.075 132.760 282.385 ;
        RECT 133.110 282.075 140.900 282.385 ;
        RECT 150.970 282.075 158.760 282.385 ;
        RECT 159.110 282.075 166.900 282.385 ;
        RECT 176.970 282.075 184.760 282.385 ;
        RECT 185.110 282.075 192.900 282.385 ;
        RECT 202.970 282.075 210.760 282.385 ;
        RECT 211.110 282.075 218.900 282.385 ;
        RECT 228.970 282.075 236.760 282.385 ;
        RECT 237.110 282.075 244.900 282.385 ;
        RECT 254.970 282.075 262.760 282.385 ;
        RECT 263.110 282.075 270.900 282.385 ;
        RECT 280.970 282.075 288.760 282.385 ;
        RECT 289.110 282.075 296.900 282.385 ;
        RECT 46.790 281.880 54.760 282.075 ;
        RECT 46.790 281.845 54.750 281.880 ;
        RECT 55.080 281.845 63.040 282.075 ;
        RECT 72.790 281.880 80.760 282.075 ;
        RECT 72.790 281.845 80.750 281.880 ;
        RECT 81.080 281.845 89.040 282.075 ;
        RECT 98.790 281.880 106.760 282.075 ;
        RECT 98.790 281.845 106.750 281.880 ;
        RECT 107.080 281.845 115.040 282.075 ;
        RECT 124.790 281.880 132.760 282.075 ;
        RECT 124.790 281.845 132.750 281.880 ;
        RECT 133.080 281.845 141.040 282.075 ;
        RECT 150.790 281.880 158.760 282.075 ;
        RECT 150.790 281.845 158.750 281.880 ;
        RECT 159.080 281.845 167.040 282.075 ;
        RECT 176.790 281.880 184.760 282.075 ;
        RECT 176.790 281.845 184.750 281.880 ;
        RECT 185.080 281.845 193.040 282.075 ;
        RECT 202.790 281.880 210.760 282.075 ;
        RECT 202.790 281.845 210.750 281.880 ;
        RECT 211.080 281.845 219.040 282.075 ;
        RECT 228.790 281.880 236.760 282.075 ;
        RECT 228.790 281.845 236.750 281.880 ;
        RECT 237.080 281.845 245.040 282.075 ;
        RECT 254.790 281.880 262.760 282.075 ;
        RECT 254.790 281.845 262.750 281.880 ;
        RECT 263.080 281.845 271.040 282.075 ;
        RECT 280.790 281.880 288.760 282.075 ;
        RECT 280.790 281.845 288.750 281.880 ;
        RECT 289.080 281.845 297.040 282.075 ;
        RECT 46.970 274.435 54.760 274.490 ;
        RECT 55.110 274.435 62.900 274.490 ;
        RECT 72.970 274.435 80.760 274.490 ;
        RECT 81.110 274.435 88.900 274.490 ;
        RECT 98.970 274.435 106.760 274.490 ;
        RECT 107.110 274.435 114.900 274.490 ;
        RECT 124.970 274.435 132.760 274.490 ;
        RECT 133.110 274.435 140.900 274.490 ;
        RECT 150.970 274.435 158.760 274.490 ;
        RECT 159.110 274.435 166.900 274.490 ;
        RECT 176.970 274.435 184.760 274.490 ;
        RECT 185.110 274.435 192.900 274.490 ;
        RECT 202.970 274.435 210.760 274.490 ;
        RECT 211.110 274.435 218.900 274.490 ;
        RECT 228.970 274.435 236.760 274.490 ;
        RECT 237.110 274.435 244.900 274.490 ;
        RECT 254.970 274.435 262.760 274.490 ;
        RECT 263.110 274.435 270.900 274.490 ;
        RECT 280.970 274.435 288.760 274.490 ;
        RECT 289.110 274.435 296.900 274.490 ;
        RECT 46.790 274.205 54.760 274.435 ;
        RECT 55.080 274.205 63.040 274.435 ;
        RECT 72.790 274.205 80.760 274.435 ;
        RECT 81.080 274.205 89.040 274.435 ;
        RECT 98.790 274.205 106.760 274.435 ;
        RECT 107.080 274.205 115.040 274.435 ;
        RECT 124.790 274.205 132.760 274.435 ;
        RECT 133.080 274.205 141.040 274.435 ;
        RECT 150.790 274.205 158.760 274.435 ;
        RECT 159.080 274.205 167.040 274.435 ;
        RECT 176.790 274.205 184.760 274.435 ;
        RECT 185.080 274.205 193.040 274.435 ;
        RECT 202.790 274.205 210.760 274.435 ;
        RECT 211.080 274.205 219.040 274.435 ;
        RECT 228.790 274.205 236.760 274.435 ;
        RECT 237.080 274.205 245.040 274.435 ;
        RECT 254.790 274.205 262.760 274.435 ;
        RECT 263.080 274.205 271.040 274.435 ;
        RECT 280.790 274.205 288.760 274.435 ;
        RECT 289.080 274.205 297.040 274.435 ;
        RECT 46.970 273.895 54.760 274.205 ;
        RECT 55.110 273.895 62.900 274.205 ;
        RECT 72.970 273.895 80.760 274.205 ;
        RECT 81.110 273.895 88.900 274.205 ;
        RECT 98.970 273.895 106.760 274.205 ;
        RECT 107.110 273.895 114.900 274.205 ;
        RECT 124.970 273.895 132.760 274.205 ;
        RECT 133.110 273.895 140.900 274.205 ;
        RECT 150.970 273.895 158.760 274.205 ;
        RECT 159.110 273.895 166.900 274.205 ;
        RECT 176.970 273.895 184.760 274.205 ;
        RECT 185.110 273.895 192.900 274.205 ;
        RECT 202.970 273.895 210.760 274.205 ;
        RECT 211.110 273.895 218.900 274.205 ;
        RECT 228.970 273.895 236.760 274.205 ;
        RECT 237.110 273.895 244.900 274.205 ;
        RECT 254.970 273.895 262.760 274.205 ;
        RECT 263.110 273.895 270.900 274.205 ;
        RECT 280.970 273.895 288.760 274.205 ;
        RECT 289.110 273.895 296.900 274.205 ;
        RECT 46.790 273.700 54.760 273.895 ;
        RECT 46.790 273.665 54.750 273.700 ;
        RECT 55.080 273.665 63.040 273.895 ;
        RECT 72.790 273.700 80.760 273.895 ;
        RECT 72.790 273.665 80.750 273.700 ;
        RECT 81.080 273.665 89.040 273.895 ;
        RECT 98.790 273.700 106.760 273.895 ;
        RECT 98.790 273.665 106.750 273.700 ;
        RECT 107.080 273.665 115.040 273.895 ;
        RECT 124.790 273.700 132.760 273.895 ;
        RECT 124.790 273.665 132.750 273.700 ;
        RECT 133.080 273.665 141.040 273.895 ;
        RECT 150.790 273.700 158.760 273.895 ;
        RECT 150.790 273.665 158.750 273.700 ;
        RECT 159.080 273.665 167.040 273.895 ;
        RECT 176.790 273.700 184.760 273.895 ;
        RECT 176.790 273.665 184.750 273.700 ;
        RECT 185.080 273.665 193.040 273.895 ;
        RECT 202.790 273.700 210.760 273.895 ;
        RECT 202.790 273.665 210.750 273.700 ;
        RECT 211.080 273.665 219.040 273.895 ;
        RECT 228.790 273.700 236.760 273.895 ;
        RECT 228.790 273.665 236.750 273.700 ;
        RECT 237.080 273.665 245.040 273.895 ;
        RECT 254.790 273.700 262.760 273.895 ;
        RECT 254.790 273.665 262.750 273.700 ;
        RECT 263.080 273.665 271.040 273.895 ;
        RECT 280.790 273.700 288.760 273.895 ;
        RECT 280.790 273.665 288.750 273.700 ;
        RECT 289.080 273.665 297.040 273.895 ;
        RECT 46.890 266.255 54.680 266.270 ;
        RECT 55.150 266.255 62.940 266.310 ;
        RECT 72.890 266.255 80.680 266.270 ;
        RECT 81.150 266.255 88.940 266.310 ;
        RECT 98.890 266.255 106.680 266.270 ;
        RECT 107.150 266.255 114.940 266.310 ;
        RECT 124.890 266.255 132.680 266.270 ;
        RECT 133.150 266.255 140.940 266.310 ;
        RECT 150.890 266.255 158.680 266.270 ;
        RECT 159.150 266.255 166.940 266.310 ;
        RECT 176.890 266.255 184.680 266.270 ;
        RECT 185.150 266.255 192.940 266.310 ;
        RECT 202.890 266.255 210.680 266.270 ;
        RECT 211.150 266.255 218.940 266.310 ;
        RECT 228.890 266.255 236.680 266.270 ;
        RECT 237.150 266.255 244.940 266.310 ;
        RECT 254.890 266.255 262.680 266.270 ;
        RECT 263.150 266.255 270.940 266.310 ;
        RECT 280.890 266.255 288.680 266.270 ;
        RECT 289.150 266.255 296.940 266.310 ;
        RECT 46.790 266.025 54.750 266.255 ;
        RECT 55.080 266.025 63.040 266.255 ;
        RECT 72.790 266.025 80.750 266.255 ;
        RECT 81.080 266.025 89.040 266.255 ;
        RECT 98.790 266.025 106.750 266.255 ;
        RECT 107.080 266.025 115.040 266.255 ;
        RECT 124.790 266.025 132.750 266.255 ;
        RECT 133.080 266.025 141.040 266.255 ;
        RECT 150.790 266.025 158.750 266.255 ;
        RECT 159.080 266.025 167.040 266.255 ;
        RECT 176.790 266.025 184.750 266.255 ;
        RECT 185.080 266.025 193.040 266.255 ;
        RECT 202.790 266.025 210.750 266.255 ;
        RECT 211.080 266.025 219.040 266.255 ;
        RECT 228.790 266.025 236.750 266.255 ;
        RECT 237.080 266.025 245.040 266.255 ;
        RECT 254.790 266.025 262.750 266.255 ;
        RECT 263.080 266.025 271.040 266.255 ;
        RECT 280.790 266.025 288.750 266.255 ;
        RECT 289.080 266.025 297.040 266.255 ;
        RECT 46.890 265.715 54.680 266.025 ;
        RECT 55.150 265.715 62.940 266.025 ;
        RECT 72.890 265.715 80.680 266.025 ;
        RECT 81.150 265.715 88.940 266.025 ;
        RECT 98.890 265.715 106.680 266.025 ;
        RECT 107.150 265.715 114.940 266.025 ;
        RECT 124.890 265.715 132.680 266.025 ;
        RECT 133.150 265.715 140.940 266.025 ;
        RECT 150.890 265.715 158.680 266.025 ;
        RECT 159.150 265.715 166.940 266.025 ;
        RECT 176.890 265.715 184.680 266.025 ;
        RECT 185.150 265.715 192.940 266.025 ;
        RECT 202.890 265.715 210.680 266.025 ;
        RECT 211.150 265.715 218.940 266.025 ;
        RECT 228.890 265.715 236.680 266.025 ;
        RECT 237.150 265.715 244.940 266.025 ;
        RECT 254.890 265.715 262.680 266.025 ;
        RECT 263.150 265.715 270.940 266.025 ;
        RECT 280.890 265.715 288.680 266.025 ;
        RECT 289.150 265.715 296.940 266.025 ;
        RECT 46.790 265.485 54.750 265.715 ;
        RECT 55.080 265.485 63.040 265.715 ;
        RECT 72.790 265.485 80.750 265.715 ;
        RECT 81.080 265.485 89.040 265.715 ;
        RECT 98.790 265.485 106.750 265.715 ;
        RECT 107.080 265.485 115.040 265.715 ;
        RECT 124.790 265.485 132.750 265.715 ;
        RECT 133.080 265.485 141.040 265.715 ;
        RECT 150.790 265.485 158.750 265.715 ;
        RECT 159.080 265.485 167.040 265.715 ;
        RECT 176.790 265.485 184.750 265.715 ;
        RECT 185.080 265.485 193.040 265.715 ;
        RECT 202.790 265.485 210.750 265.715 ;
        RECT 211.080 265.485 219.040 265.715 ;
        RECT 228.790 265.485 236.750 265.715 ;
        RECT 237.080 265.485 245.040 265.715 ;
        RECT 254.790 265.485 262.750 265.715 ;
        RECT 263.080 265.485 271.040 265.715 ;
        RECT 280.790 265.485 288.750 265.715 ;
        RECT 289.080 265.485 297.040 265.715 ;
        RECT 46.890 265.480 54.680 265.485 ;
        RECT 72.890 265.480 80.680 265.485 ;
        RECT 98.890 265.480 106.680 265.485 ;
        RECT 124.890 265.480 132.680 265.485 ;
        RECT 150.890 265.480 158.680 265.485 ;
        RECT 176.890 265.480 184.680 265.485 ;
        RECT 202.890 265.480 210.680 265.485 ;
        RECT 228.890 265.480 236.680 265.485 ;
        RECT 254.890 265.480 262.680 265.485 ;
        RECT 280.890 265.480 288.680 265.485 ;
        RECT 46.890 258.075 54.680 258.130 ;
        RECT 55.270 258.075 63.060 258.090 ;
        RECT 72.890 258.075 80.680 258.130 ;
        RECT 81.270 258.075 89.060 258.090 ;
        RECT 98.890 258.075 106.680 258.130 ;
        RECT 107.270 258.075 115.060 258.090 ;
        RECT 124.890 258.075 132.680 258.130 ;
        RECT 133.270 258.075 141.060 258.090 ;
        RECT 150.890 258.075 158.680 258.130 ;
        RECT 159.270 258.075 167.060 258.090 ;
        RECT 176.890 258.075 184.680 258.130 ;
        RECT 185.270 258.075 193.060 258.090 ;
        RECT 202.890 258.075 210.680 258.130 ;
        RECT 211.270 258.075 219.060 258.090 ;
        RECT 228.890 258.075 236.680 258.130 ;
        RECT 237.270 258.075 245.060 258.090 ;
        RECT 254.890 258.075 262.680 258.130 ;
        RECT 263.270 258.075 271.060 258.090 ;
        RECT 280.890 258.075 288.680 258.130 ;
        RECT 289.270 258.075 297.060 258.090 ;
        RECT 46.790 257.845 54.750 258.075 ;
        RECT 55.080 257.845 63.060 258.075 ;
        RECT 72.790 257.845 80.750 258.075 ;
        RECT 81.080 257.845 89.060 258.075 ;
        RECT 98.790 257.845 106.750 258.075 ;
        RECT 107.080 257.845 115.060 258.075 ;
        RECT 124.790 257.845 132.750 258.075 ;
        RECT 133.080 257.845 141.060 258.075 ;
        RECT 150.790 257.845 158.750 258.075 ;
        RECT 159.080 257.845 167.060 258.075 ;
        RECT 176.790 257.845 184.750 258.075 ;
        RECT 185.080 257.845 193.060 258.075 ;
        RECT 202.790 257.845 210.750 258.075 ;
        RECT 211.080 257.845 219.060 258.075 ;
        RECT 228.790 257.845 236.750 258.075 ;
        RECT 237.080 257.845 245.060 258.075 ;
        RECT 254.790 257.845 262.750 258.075 ;
        RECT 263.080 257.845 271.060 258.075 ;
        RECT 280.790 257.845 288.750 258.075 ;
        RECT 289.080 257.845 297.060 258.075 ;
        RECT 46.890 257.535 54.680 257.845 ;
        RECT 55.270 257.535 63.060 257.845 ;
        RECT 72.890 257.535 80.680 257.845 ;
        RECT 81.270 257.535 89.060 257.845 ;
        RECT 98.890 257.535 106.680 257.845 ;
        RECT 107.270 257.535 115.060 257.845 ;
        RECT 124.890 257.535 132.680 257.845 ;
        RECT 133.270 257.535 141.060 257.845 ;
        RECT 150.890 257.535 158.680 257.845 ;
        RECT 159.270 257.535 167.060 257.845 ;
        RECT 176.890 257.535 184.680 257.845 ;
        RECT 185.270 257.535 193.060 257.845 ;
        RECT 202.890 257.535 210.680 257.845 ;
        RECT 211.270 257.535 219.060 257.845 ;
        RECT 228.890 257.535 236.680 257.845 ;
        RECT 237.270 257.535 245.060 257.845 ;
        RECT 254.890 257.535 262.680 257.845 ;
        RECT 263.270 257.535 271.060 257.845 ;
        RECT 280.890 257.535 288.680 257.845 ;
        RECT 289.270 257.535 297.060 257.845 ;
        RECT 46.790 257.305 54.750 257.535 ;
        RECT 55.080 257.305 63.060 257.535 ;
        RECT 72.790 257.305 80.750 257.535 ;
        RECT 81.080 257.305 89.060 257.535 ;
        RECT 98.790 257.305 106.750 257.535 ;
        RECT 107.080 257.305 115.060 257.535 ;
        RECT 124.790 257.305 132.750 257.535 ;
        RECT 133.080 257.305 141.060 257.535 ;
        RECT 150.790 257.305 158.750 257.535 ;
        RECT 159.080 257.305 167.060 257.535 ;
        RECT 176.790 257.305 184.750 257.535 ;
        RECT 185.080 257.305 193.060 257.535 ;
        RECT 202.790 257.305 210.750 257.535 ;
        RECT 211.080 257.305 219.060 257.535 ;
        RECT 228.790 257.305 236.750 257.535 ;
        RECT 237.080 257.305 245.060 257.535 ;
        RECT 254.790 257.305 262.750 257.535 ;
        RECT 263.080 257.305 271.060 257.535 ;
        RECT 280.790 257.305 288.750 257.535 ;
        RECT 289.080 257.305 297.060 257.535 ;
        RECT 55.270 257.300 63.060 257.305 ;
        RECT 81.270 257.300 89.060 257.305 ;
        RECT 107.270 257.300 115.060 257.305 ;
        RECT 133.270 257.300 141.060 257.305 ;
        RECT 159.270 257.300 167.060 257.305 ;
        RECT 185.270 257.300 193.060 257.305 ;
        RECT 211.270 257.300 219.060 257.305 ;
        RECT 237.270 257.300 245.060 257.305 ;
        RECT 263.270 257.300 271.060 257.305 ;
        RECT 289.270 257.300 297.060 257.305 ;
        RECT 46.970 249.895 54.760 249.910 ;
        RECT 55.310 249.895 63.100 249.910 ;
        RECT 72.970 249.895 80.760 249.910 ;
        RECT 81.310 249.895 89.100 249.910 ;
        RECT 98.970 249.895 106.760 249.910 ;
        RECT 107.310 249.895 115.100 249.910 ;
        RECT 124.970 249.895 132.760 249.910 ;
        RECT 133.310 249.895 141.100 249.910 ;
        RECT 150.970 249.895 158.760 249.910 ;
        RECT 159.310 249.895 167.100 249.910 ;
        RECT 176.970 249.895 184.760 249.910 ;
        RECT 185.310 249.895 193.100 249.910 ;
        RECT 202.970 249.895 210.760 249.910 ;
        RECT 211.310 249.895 219.100 249.910 ;
        RECT 228.970 249.895 236.760 249.910 ;
        RECT 237.310 249.895 245.100 249.910 ;
        RECT 254.970 249.895 262.760 249.910 ;
        RECT 263.310 249.895 271.100 249.910 ;
        RECT 280.970 249.895 288.760 249.910 ;
        RECT 289.310 249.895 297.100 249.910 ;
        RECT 46.790 249.665 54.760 249.895 ;
        RECT 55.080 249.665 63.100 249.895 ;
        RECT 72.790 249.665 80.760 249.895 ;
        RECT 81.080 249.665 89.100 249.895 ;
        RECT 98.790 249.665 106.760 249.895 ;
        RECT 107.080 249.665 115.100 249.895 ;
        RECT 124.790 249.665 132.760 249.895 ;
        RECT 133.080 249.665 141.100 249.895 ;
        RECT 150.790 249.665 158.760 249.895 ;
        RECT 159.080 249.665 167.100 249.895 ;
        RECT 176.790 249.665 184.760 249.895 ;
        RECT 185.080 249.665 193.100 249.895 ;
        RECT 202.790 249.665 210.760 249.895 ;
        RECT 211.080 249.665 219.100 249.895 ;
        RECT 228.790 249.665 236.760 249.895 ;
        RECT 237.080 249.665 245.100 249.895 ;
        RECT 254.790 249.665 262.760 249.895 ;
        RECT 263.080 249.665 271.100 249.895 ;
        RECT 280.790 249.665 288.760 249.895 ;
        RECT 289.080 249.665 297.100 249.895 ;
        RECT 46.970 249.355 54.760 249.665 ;
        RECT 55.310 249.355 63.100 249.665 ;
        RECT 72.970 249.355 80.760 249.665 ;
        RECT 81.310 249.355 89.100 249.665 ;
        RECT 98.970 249.355 106.760 249.665 ;
        RECT 107.310 249.355 115.100 249.665 ;
        RECT 124.970 249.355 132.760 249.665 ;
        RECT 133.310 249.355 141.100 249.665 ;
        RECT 150.970 249.355 158.760 249.665 ;
        RECT 159.310 249.355 167.100 249.665 ;
        RECT 176.970 249.355 184.760 249.665 ;
        RECT 185.310 249.355 193.100 249.665 ;
        RECT 202.970 249.355 210.760 249.665 ;
        RECT 211.310 249.355 219.100 249.665 ;
        RECT 228.970 249.355 236.760 249.665 ;
        RECT 237.310 249.355 245.100 249.665 ;
        RECT 254.970 249.355 262.760 249.665 ;
        RECT 263.310 249.355 271.100 249.665 ;
        RECT 280.970 249.355 288.760 249.665 ;
        RECT 289.310 249.355 297.100 249.665 ;
        RECT 46.790 249.125 54.760 249.355 ;
        RECT 55.080 249.125 63.100 249.355 ;
        RECT 72.790 249.125 80.760 249.355 ;
        RECT 81.080 249.125 89.100 249.355 ;
        RECT 98.790 249.125 106.760 249.355 ;
        RECT 107.080 249.125 115.100 249.355 ;
        RECT 124.790 249.125 132.760 249.355 ;
        RECT 133.080 249.125 141.100 249.355 ;
        RECT 150.790 249.125 158.760 249.355 ;
        RECT 159.080 249.125 167.100 249.355 ;
        RECT 176.790 249.125 184.760 249.355 ;
        RECT 185.080 249.125 193.100 249.355 ;
        RECT 202.790 249.125 210.760 249.355 ;
        RECT 211.080 249.125 219.100 249.355 ;
        RECT 228.790 249.125 236.760 249.355 ;
        RECT 237.080 249.125 245.100 249.355 ;
        RECT 254.790 249.125 262.760 249.355 ;
        RECT 263.080 249.125 271.100 249.355 ;
        RECT 280.790 249.125 288.760 249.355 ;
        RECT 289.080 249.125 297.100 249.355 ;
        RECT 46.970 249.120 54.760 249.125 ;
        RECT 55.310 249.120 63.100 249.125 ;
        RECT 72.970 249.120 80.760 249.125 ;
        RECT 81.310 249.120 89.100 249.125 ;
        RECT 98.970 249.120 106.760 249.125 ;
        RECT 107.310 249.120 115.100 249.125 ;
        RECT 124.970 249.120 132.760 249.125 ;
        RECT 133.310 249.120 141.100 249.125 ;
        RECT 150.970 249.120 158.760 249.125 ;
        RECT 159.310 249.120 167.100 249.125 ;
        RECT 176.970 249.120 184.760 249.125 ;
        RECT 185.310 249.120 193.100 249.125 ;
        RECT 202.970 249.120 210.760 249.125 ;
        RECT 211.310 249.120 219.100 249.125 ;
        RECT 228.970 249.120 236.760 249.125 ;
        RECT 237.310 249.120 245.100 249.125 ;
        RECT 254.970 249.120 262.760 249.125 ;
        RECT 263.310 249.120 271.100 249.125 ;
        RECT 280.970 249.120 288.760 249.125 ;
        RECT 289.310 249.120 297.100 249.125 ;
        RECT 46.890 241.715 54.680 241.730 ;
        RECT 55.270 241.715 63.060 241.770 ;
        RECT 72.890 241.715 80.680 241.730 ;
        RECT 81.270 241.715 89.060 241.770 ;
        RECT 98.890 241.715 106.680 241.730 ;
        RECT 107.270 241.715 115.060 241.770 ;
        RECT 124.890 241.715 132.680 241.730 ;
        RECT 133.270 241.715 141.060 241.770 ;
        RECT 150.890 241.715 158.680 241.730 ;
        RECT 159.270 241.715 167.060 241.770 ;
        RECT 176.890 241.715 184.680 241.730 ;
        RECT 185.270 241.715 193.060 241.770 ;
        RECT 202.890 241.715 210.680 241.730 ;
        RECT 211.270 241.715 219.060 241.770 ;
        RECT 228.890 241.715 236.680 241.730 ;
        RECT 237.270 241.715 245.060 241.770 ;
        RECT 254.890 241.715 262.680 241.730 ;
        RECT 263.270 241.715 271.060 241.770 ;
        RECT 280.890 241.715 288.680 241.730 ;
        RECT 289.270 241.715 297.060 241.770 ;
        RECT 46.790 241.485 54.750 241.715 ;
        RECT 55.080 241.485 63.060 241.715 ;
        RECT 72.790 241.485 80.750 241.715 ;
        RECT 81.080 241.485 89.060 241.715 ;
        RECT 98.790 241.485 106.750 241.715 ;
        RECT 107.080 241.485 115.060 241.715 ;
        RECT 124.790 241.485 132.750 241.715 ;
        RECT 133.080 241.485 141.060 241.715 ;
        RECT 150.790 241.485 158.750 241.715 ;
        RECT 159.080 241.485 167.060 241.715 ;
        RECT 176.790 241.485 184.750 241.715 ;
        RECT 185.080 241.485 193.060 241.715 ;
        RECT 202.790 241.485 210.750 241.715 ;
        RECT 211.080 241.485 219.060 241.715 ;
        RECT 228.790 241.485 236.750 241.715 ;
        RECT 237.080 241.485 245.060 241.715 ;
        RECT 254.790 241.485 262.750 241.715 ;
        RECT 263.080 241.485 271.060 241.715 ;
        RECT 280.790 241.485 288.750 241.715 ;
        RECT 289.080 241.485 297.060 241.715 ;
        RECT 46.890 241.175 54.680 241.485 ;
        RECT 55.270 241.175 63.060 241.485 ;
        RECT 72.890 241.175 80.680 241.485 ;
        RECT 81.270 241.175 89.060 241.485 ;
        RECT 98.890 241.175 106.680 241.485 ;
        RECT 107.270 241.175 115.060 241.485 ;
        RECT 124.890 241.175 132.680 241.485 ;
        RECT 133.270 241.175 141.060 241.485 ;
        RECT 150.890 241.175 158.680 241.485 ;
        RECT 159.270 241.175 167.060 241.485 ;
        RECT 176.890 241.175 184.680 241.485 ;
        RECT 185.270 241.175 193.060 241.485 ;
        RECT 202.890 241.175 210.680 241.485 ;
        RECT 211.270 241.175 219.060 241.485 ;
        RECT 228.890 241.175 236.680 241.485 ;
        RECT 237.270 241.175 245.060 241.485 ;
        RECT 254.890 241.175 262.680 241.485 ;
        RECT 263.270 241.175 271.060 241.485 ;
        RECT 280.890 241.175 288.680 241.485 ;
        RECT 289.270 241.175 297.060 241.485 ;
        RECT 46.790 240.945 54.750 241.175 ;
        RECT 55.080 240.980 63.060 241.175 ;
        RECT 55.080 240.945 63.040 240.980 ;
        RECT 72.790 240.945 80.750 241.175 ;
        RECT 81.080 240.980 89.060 241.175 ;
        RECT 81.080 240.945 89.040 240.980 ;
        RECT 98.790 240.945 106.750 241.175 ;
        RECT 107.080 240.980 115.060 241.175 ;
        RECT 107.080 240.945 115.040 240.980 ;
        RECT 124.790 240.945 132.750 241.175 ;
        RECT 133.080 240.980 141.060 241.175 ;
        RECT 133.080 240.945 141.040 240.980 ;
        RECT 150.790 240.945 158.750 241.175 ;
        RECT 159.080 240.980 167.060 241.175 ;
        RECT 159.080 240.945 167.040 240.980 ;
        RECT 176.790 240.945 184.750 241.175 ;
        RECT 185.080 240.980 193.060 241.175 ;
        RECT 185.080 240.945 193.040 240.980 ;
        RECT 202.790 240.945 210.750 241.175 ;
        RECT 211.080 240.980 219.060 241.175 ;
        RECT 211.080 240.945 219.040 240.980 ;
        RECT 228.790 240.945 236.750 241.175 ;
        RECT 237.080 240.980 245.060 241.175 ;
        RECT 237.080 240.945 245.040 240.980 ;
        RECT 254.790 240.945 262.750 241.175 ;
        RECT 263.080 240.980 271.060 241.175 ;
        RECT 263.080 240.945 271.040 240.980 ;
        RECT 280.790 240.945 288.750 241.175 ;
        RECT 289.080 240.980 297.060 241.175 ;
        RECT 289.080 240.945 297.040 240.980 ;
        RECT 46.890 240.940 54.680 240.945 ;
        RECT 72.890 240.940 80.680 240.945 ;
        RECT 98.890 240.940 106.680 240.945 ;
        RECT 124.890 240.940 132.680 240.945 ;
        RECT 150.890 240.940 158.680 240.945 ;
        RECT 176.890 240.940 184.680 240.945 ;
        RECT 202.890 240.940 210.680 240.945 ;
        RECT 228.890 240.940 236.680 240.945 ;
        RECT 254.890 240.940 262.680 240.945 ;
        RECT 280.890 240.940 288.680 240.945 ;
        RECT 47.010 233.535 54.800 233.550 ;
        RECT 55.150 233.535 62.940 233.590 ;
        RECT 73.010 233.535 80.800 233.550 ;
        RECT 81.150 233.535 88.940 233.590 ;
        RECT 99.010 233.535 106.800 233.550 ;
        RECT 107.150 233.535 114.940 233.590 ;
        RECT 125.010 233.535 132.800 233.550 ;
        RECT 133.150 233.535 140.940 233.590 ;
        RECT 151.010 233.535 158.800 233.550 ;
        RECT 159.150 233.535 166.940 233.590 ;
        RECT 177.010 233.535 184.800 233.550 ;
        RECT 185.150 233.535 192.940 233.590 ;
        RECT 203.010 233.535 210.800 233.550 ;
        RECT 211.150 233.535 218.940 233.590 ;
        RECT 229.010 233.535 236.800 233.550 ;
        RECT 237.150 233.535 244.940 233.590 ;
        RECT 255.010 233.535 262.800 233.550 ;
        RECT 263.150 233.535 270.940 233.590 ;
        RECT 281.010 233.535 288.800 233.550 ;
        RECT 289.150 233.535 296.940 233.590 ;
        RECT 46.790 233.305 54.800 233.535 ;
        RECT 55.080 233.305 63.040 233.535 ;
        RECT 72.790 233.305 80.800 233.535 ;
        RECT 81.080 233.305 89.040 233.535 ;
        RECT 98.790 233.305 106.800 233.535 ;
        RECT 107.080 233.305 115.040 233.535 ;
        RECT 124.790 233.305 132.800 233.535 ;
        RECT 133.080 233.305 141.040 233.535 ;
        RECT 150.790 233.305 158.800 233.535 ;
        RECT 159.080 233.305 167.040 233.535 ;
        RECT 176.790 233.305 184.800 233.535 ;
        RECT 185.080 233.305 193.040 233.535 ;
        RECT 202.790 233.305 210.800 233.535 ;
        RECT 211.080 233.305 219.040 233.535 ;
        RECT 228.790 233.305 236.800 233.535 ;
        RECT 237.080 233.305 245.040 233.535 ;
        RECT 254.790 233.305 262.800 233.535 ;
        RECT 263.080 233.305 271.040 233.535 ;
        RECT 280.790 233.305 288.800 233.535 ;
        RECT 289.080 233.305 297.040 233.535 ;
        RECT 47.010 232.995 54.800 233.305 ;
        RECT 55.150 232.995 62.940 233.305 ;
        RECT 73.010 232.995 80.800 233.305 ;
        RECT 81.150 232.995 88.940 233.305 ;
        RECT 99.010 232.995 106.800 233.305 ;
        RECT 107.150 232.995 114.940 233.305 ;
        RECT 125.010 232.995 132.800 233.305 ;
        RECT 133.150 232.995 140.940 233.305 ;
        RECT 151.010 232.995 158.800 233.305 ;
        RECT 159.150 232.995 166.940 233.305 ;
        RECT 177.010 232.995 184.800 233.305 ;
        RECT 185.150 232.995 192.940 233.305 ;
        RECT 203.010 232.995 210.800 233.305 ;
        RECT 211.150 232.995 218.940 233.305 ;
        RECT 229.010 232.995 236.800 233.305 ;
        RECT 237.150 232.995 244.940 233.305 ;
        RECT 255.010 232.995 262.800 233.305 ;
        RECT 263.150 232.995 270.940 233.305 ;
        RECT 281.010 232.995 288.800 233.305 ;
        RECT 289.150 232.995 296.940 233.305 ;
        RECT 46.790 232.765 54.800 232.995 ;
        RECT 55.080 232.765 63.040 232.995 ;
        RECT 72.790 232.765 80.800 232.995 ;
        RECT 81.080 232.765 89.040 232.995 ;
        RECT 98.790 232.765 106.800 232.995 ;
        RECT 107.080 232.765 115.040 232.995 ;
        RECT 124.790 232.765 132.800 232.995 ;
        RECT 133.080 232.765 141.040 232.995 ;
        RECT 150.790 232.765 158.800 232.995 ;
        RECT 159.080 232.765 167.040 232.995 ;
        RECT 176.790 232.765 184.800 232.995 ;
        RECT 185.080 232.765 193.040 232.995 ;
        RECT 202.790 232.765 210.800 232.995 ;
        RECT 211.080 232.765 219.040 232.995 ;
        RECT 228.790 232.765 236.800 232.995 ;
        RECT 237.080 232.765 245.040 232.995 ;
        RECT 254.790 232.765 262.800 232.995 ;
        RECT 263.080 232.765 271.040 232.995 ;
        RECT 280.790 232.765 288.800 232.995 ;
        RECT 289.080 232.765 297.040 232.995 ;
        RECT 47.010 232.760 54.800 232.765 ;
        RECT 73.010 232.760 80.800 232.765 ;
        RECT 99.010 232.760 106.800 232.765 ;
        RECT 125.010 232.760 132.800 232.765 ;
        RECT 151.010 232.760 158.800 232.765 ;
        RECT 177.010 232.760 184.800 232.765 ;
        RECT 203.010 232.760 210.800 232.765 ;
        RECT 229.010 232.760 236.800 232.765 ;
        RECT 255.010 232.760 262.800 232.765 ;
        RECT 281.010 232.760 288.800 232.765 ;
        RECT 46.970 225.420 54.660 225.450 ;
        RECT 72.970 225.420 80.660 225.450 ;
        RECT 98.970 225.420 106.660 225.450 ;
        RECT 124.970 225.420 132.660 225.450 ;
        RECT 150.970 225.420 158.660 225.450 ;
        RECT 176.970 225.420 184.660 225.450 ;
        RECT 202.970 225.420 210.660 225.450 ;
        RECT 228.970 225.420 236.660 225.450 ;
        RECT 254.970 225.420 262.660 225.450 ;
        RECT 280.970 225.420 288.660 225.450 ;
        RECT 46.970 225.355 54.760 225.420 ;
        RECT 55.310 225.355 63.100 225.410 ;
        RECT 72.970 225.355 80.760 225.420 ;
        RECT 81.310 225.355 89.100 225.410 ;
        RECT 98.970 225.355 106.760 225.420 ;
        RECT 107.310 225.355 115.100 225.410 ;
        RECT 124.970 225.355 132.760 225.420 ;
        RECT 133.310 225.355 141.100 225.410 ;
        RECT 150.970 225.355 158.760 225.420 ;
        RECT 159.310 225.355 167.100 225.410 ;
        RECT 176.970 225.355 184.760 225.420 ;
        RECT 185.310 225.355 193.100 225.410 ;
        RECT 202.970 225.355 210.760 225.420 ;
        RECT 211.310 225.355 219.100 225.410 ;
        RECT 228.970 225.355 236.760 225.420 ;
        RECT 237.310 225.355 245.100 225.410 ;
        RECT 254.970 225.355 262.760 225.420 ;
        RECT 263.310 225.355 271.100 225.410 ;
        RECT 280.970 225.355 288.760 225.420 ;
        RECT 289.310 225.355 297.100 225.410 ;
        RECT 46.790 225.125 54.760 225.355 ;
        RECT 55.080 225.125 63.100 225.355 ;
        RECT 72.790 225.125 80.760 225.355 ;
        RECT 81.080 225.125 89.100 225.355 ;
        RECT 98.790 225.125 106.760 225.355 ;
        RECT 107.080 225.125 115.100 225.355 ;
        RECT 124.790 225.125 132.760 225.355 ;
        RECT 133.080 225.125 141.100 225.355 ;
        RECT 150.790 225.125 158.760 225.355 ;
        RECT 159.080 225.125 167.100 225.355 ;
        RECT 176.790 225.125 184.760 225.355 ;
        RECT 185.080 225.125 193.100 225.355 ;
        RECT 202.790 225.125 210.760 225.355 ;
        RECT 211.080 225.125 219.100 225.355 ;
        RECT 228.790 225.125 236.760 225.355 ;
        RECT 237.080 225.125 245.100 225.355 ;
        RECT 254.790 225.125 262.760 225.355 ;
        RECT 263.080 225.125 271.100 225.355 ;
        RECT 280.790 225.125 288.760 225.355 ;
        RECT 289.080 225.125 297.100 225.355 ;
        RECT 46.970 224.815 54.760 225.125 ;
        RECT 55.310 224.815 63.100 225.125 ;
        RECT 72.970 224.815 80.760 225.125 ;
        RECT 81.310 224.815 89.100 225.125 ;
        RECT 98.970 224.815 106.760 225.125 ;
        RECT 107.310 224.815 115.100 225.125 ;
        RECT 124.970 224.815 132.760 225.125 ;
        RECT 133.310 224.815 141.100 225.125 ;
        RECT 150.970 224.815 158.760 225.125 ;
        RECT 159.310 224.815 167.100 225.125 ;
        RECT 176.970 224.815 184.760 225.125 ;
        RECT 185.310 224.815 193.100 225.125 ;
        RECT 202.970 224.815 210.760 225.125 ;
        RECT 211.310 224.815 219.100 225.125 ;
        RECT 228.970 224.815 236.760 225.125 ;
        RECT 237.310 224.815 245.100 225.125 ;
        RECT 254.970 224.815 262.760 225.125 ;
        RECT 263.310 224.815 271.100 225.125 ;
        RECT 280.970 224.815 288.760 225.125 ;
        RECT 289.310 224.815 297.100 225.125 ;
        RECT 46.790 224.660 54.760 224.815 ;
        RECT 46.790 224.585 54.750 224.660 ;
        RECT 55.080 224.620 63.100 224.815 ;
        RECT 72.790 224.660 80.760 224.815 ;
        RECT 55.080 224.585 63.040 224.620 ;
        RECT 72.790 224.585 80.750 224.660 ;
        RECT 81.080 224.620 89.100 224.815 ;
        RECT 98.790 224.660 106.760 224.815 ;
        RECT 81.080 224.585 89.040 224.620 ;
        RECT 98.790 224.585 106.750 224.660 ;
        RECT 107.080 224.620 115.100 224.815 ;
        RECT 124.790 224.660 132.760 224.815 ;
        RECT 107.080 224.585 115.040 224.620 ;
        RECT 124.790 224.585 132.750 224.660 ;
        RECT 133.080 224.620 141.100 224.815 ;
        RECT 150.790 224.660 158.760 224.815 ;
        RECT 133.080 224.585 141.040 224.620 ;
        RECT 150.790 224.585 158.750 224.660 ;
        RECT 159.080 224.620 167.100 224.815 ;
        RECT 176.790 224.660 184.760 224.815 ;
        RECT 159.080 224.585 167.040 224.620 ;
        RECT 176.790 224.585 184.750 224.660 ;
        RECT 185.080 224.620 193.100 224.815 ;
        RECT 202.790 224.660 210.760 224.815 ;
        RECT 185.080 224.585 193.040 224.620 ;
        RECT 202.790 224.585 210.750 224.660 ;
        RECT 211.080 224.620 219.100 224.815 ;
        RECT 228.790 224.660 236.760 224.815 ;
        RECT 211.080 224.585 219.040 224.620 ;
        RECT 228.790 224.585 236.750 224.660 ;
        RECT 237.080 224.620 245.100 224.815 ;
        RECT 254.790 224.660 262.760 224.815 ;
        RECT 237.080 224.585 245.040 224.620 ;
        RECT 254.790 224.585 262.750 224.660 ;
        RECT 263.080 224.620 271.100 224.815 ;
        RECT 280.790 224.660 288.760 224.815 ;
        RECT 263.080 224.585 271.040 224.620 ;
        RECT 280.790 224.585 288.750 224.660 ;
        RECT 289.080 224.620 297.100 224.815 ;
        RECT 289.080 224.585 297.040 224.620 ;
        RECT 46.970 217.175 54.760 217.190 ;
        RECT 55.190 217.175 62.980 217.230 ;
        RECT 72.970 217.175 80.760 217.190 ;
        RECT 81.190 217.175 88.980 217.230 ;
        RECT 98.970 217.175 106.760 217.190 ;
        RECT 107.190 217.175 114.980 217.230 ;
        RECT 124.970 217.175 132.760 217.190 ;
        RECT 133.190 217.175 140.980 217.230 ;
        RECT 150.970 217.175 158.760 217.190 ;
        RECT 159.190 217.175 166.980 217.230 ;
        RECT 176.970 217.175 184.760 217.190 ;
        RECT 185.190 217.175 192.980 217.230 ;
        RECT 202.970 217.175 210.760 217.190 ;
        RECT 211.190 217.175 218.980 217.230 ;
        RECT 228.970 217.175 236.760 217.190 ;
        RECT 237.190 217.175 244.980 217.230 ;
        RECT 254.970 217.175 262.760 217.190 ;
        RECT 263.190 217.175 270.980 217.230 ;
        RECT 280.970 217.175 288.760 217.190 ;
        RECT 289.190 217.175 296.980 217.230 ;
        RECT 46.790 216.945 54.760 217.175 ;
        RECT 55.080 216.945 63.040 217.175 ;
        RECT 72.790 216.945 80.760 217.175 ;
        RECT 81.080 216.945 89.040 217.175 ;
        RECT 98.790 216.945 106.760 217.175 ;
        RECT 107.080 216.945 115.040 217.175 ;
        RECT 124.790 216.945 132.760 217.175 ;
        RECT 133.080 216.945 141.040 217.175 ;
        RECT 150.790 216.945 158.760 217.175 ;
        RECT 159.080 216.945 167.040 217.175 ;
        RECT 176.790 216.945 184.760 217.175 ;
        RECT 185.080 216.945 193.040 217.175 ;
        RECT 202.790 216.945 210.760 217.175 ;
        RECT 211.080 216.945 219.040 217.175 ;
        RECT 228.790 216.945 236.760 217.175 ;
        RECT 237.080 216.945 245.040 217.175 ;
        RECT 254.790 216.945 262.760 217.175 ;
        RECT 263.080 216.945 271.040 217.175 ;
        RECT 280.790 216.945 288.760 217.175 ;
        RECT 289.080 216.945 297.040 217.175 ;
        RECT 46.970 216.635 54.760 216.945 ;
        RECT 55.190 216.635 62.980 216.945 ;
        RECT 72.970 216.635 80.760 216.945 ;
        RECT 81.190 216.635 88.980 216.945 ;
        RECT 98.970 216.635 106.760 216.945 ;
        RECT 107.190 216.635 114.980 216.945 ;
        RECT 124.970 216.635 132.760 216.945 ;
        RECT 133.190 216.635 140.980 216.945 ;
        RECT 150.970 216.635 158.760 216.945 ;
        RECT 159.190 216.635 166.980 216.945 ;
        RECT 176.970 216.635 184.760 216.945 ;
        RECT 185.190 216.635 192.980 216.945 ;
        RECT 202.970 216.635 210.760 216.945 ;
        RECT 211.190 216.635 218.980 216.945 ;
        RECT 228.970 216.635 236.760 216.945 ;
        RECT 237.190 216.635 244.980 216.945 ;
        RECT 254.970 216.635 262.760 216.945 ;
        RECT 263.190 216.635 270.980 216.945 ;
        RECT 280.970 216.635 288.760 216.945 ;
        RECT 289.190 216.635 296.980 216.945 ;
        RECT 46.790 216.405 54.760 216.635 ;
        RECT 55.080 216.405 63.040 216.635 ;
        RECT 72.790 216.405 80.760 216.635 ;
        RECT 81.080 216.405 89.040 216.635 ;
        RECT 98.790 216.405 106.760 216.635 ;
        RECT 107.080 216.405 115.040 216.635 ;
        RECT 124.790 216.405 132.760 216.635 ;
        RECT 133.080 216.405 141.040 216.635 ;
        RECT 150.790 216.405 158.760 216.635 ;
        RECT 159.080 216.405 167.040 216.635 ;
        RECT 176.790 216.405 184.760 216.635 ;
        RECT 185.080 216.405 193.040 216.635 ;
        RECT 202.790 216.405 210.760 216.635 ;
        RECT 211.080 216.405 219.040 216.635 ;
        RECT 228.790 216.405 236.760 216.635 ;
        RECT 237.080 216.405 245.040 216.635 ;
        RECT 254.790 216.405 262.760 216.635 ;
        RECT 263.080 216.405 271.040 216.635 ;
        RECT 280.790 216.405 288.760 216.635 ;
        RECT 289.080 216.405 297.040 216.635 ;
        RECT 46.970 216.400 54.760 216.405 ;
        RECT 72.970 216.400 80.760 216.405 ;
        RECT 98.970 216.400 106.760 216.405 ;
        RECT 124.970 216.400 132.760 216.405 ;
        RECT 150.970 216.400 158.760 216.405 ;
        RECT 176.970 216.400 184.760 216.405 ;
        RECT 202.970 216.400 210.760 216.405 ;
        RECT 228.970 216.400 236.760 216.405 ;
        RECT 254.970 216.400 262.760 216.405 ;
        RECT 280.970 216.400 288.760 216.405 ;
        RECT 46.970 208.995 54.760 209.010 ;
        RECT 55.270 208.995 63.060 209.050 ;
        RECT 72.970 208.995 80.760 209.010 ;
        RECT 81.270 208.995 89.060 209.050 ;
        RECT 98.970 208.995 106.760 209.010 ;
        RECT 107.270 208.995 115.060 209.050 ;
        RECT 124.970 208.995 132.760 209.010 ;
        RECT 133.270 208.995 141.060 209.050 ;
        RECT 150.970 208.995 158.760 209.010 ;
        RECT 159.270 208.995 167.060 209.050 ;
        RECT 176.970 208.995 184.760 209.010 ;
        RECT 185.270 208.995 193.060 209.050 ;
        RECT 202.970 208.995 210.760 209.010 ;
        RECT 211.270 208.995 219.060 209.050 ;
        RECT 228.970 208.995 236.760 209.010 ;
        RECT 237.270 208.995 245.060 209.050 ;
        RECT 254.970 208.995 262.760 209.010 ;
        RECT 263.270 208.995 271.060 209.050 ;
        RECT 280.970 208.995 288.760 209.010 ;
        RECT 289.270 208.995 297.060 209.050 ;
        RECT 46.790 208.765 54.760 208.995 ;
        RECT 55.080 208.765 63.060 208.995 ;
        RECT 72.790 208.765 80.760 208.995 ;
        RECT 81.080 208.765 89.060 208.995 ;
        RECT 98.790 208.765 106.760 208.995 ;
        RECT 107.080 208.765 115.060 208.995 ;
        RECT 124.790 208.765 132.760 208.995 ;
        RECT 133.080 208.765 141.060 208.995 ;
        RECT 150.790 208.765 158.760 208.995 ;
        RECT 159.080 208.765 167.060 208.995 ;
        RECT 176.790 208.765 184.760 208.995 ;
        RECT 185.080 208.765 193.060 208.995 ;
        RECT 202.790 208.765 210.760 208.995 ;
        RECT 211.080 208.765 219.060 208.995 ;
        RECT 228.790 208.765 236.760 208.995 ;
        RECT 237.080 208.765 245.060 208.995 ;
        RECT 254.790 208.765 262.760 208.995 ;
        RECT 263.080 208.765 271.060 208.995 ;
        RECT 280.790 208.765 288.760 208.995 ;
        RECT 289.080 208.765 297.060 208.995 ;
        RECT 586.510 208.810 592.150 208.890 ;
        RECT 46.970 208.455 54.760 208.765 ;
        RECT 55.270 208.455 63.060 208.765 ;
        RECT 72.970 208.455 80.760 208.765 ;
        RECT 81.270 208.455 89.060 208.765 ;
        RECT 98.970 208.455 106.760 208.765 ;
        RECT 107.270 208.455 115.060 208.765 ;
        RECT 124.970 208.455 132.760 208.765 ;
        RECT 133.270 208.455 141.060 208.765 ;
        RECT 150.970 208.455 158.760 208.765 ;
        RECT 159.270 208.455 167.060 208.765 ;
        RECT 176.970 208.455 184.760 208.765 ;
        RECT 185.270 208.455 193.060 208.765 ;
        RECT 202.970 208.455 210.760 208.765 ;
        RECT 211.270 208.455 219.060 208.765 ;
        RECT 228.970 208.455 236.760 208.765 ;
        RECT 237.270 208.455 245.060 208.765 ;
        RECT 254.970 208.455 262.760 208.765 ;
        RECT 263.270 208.455 271.060 208.765 ;
        RECT 280.970 208.455 288.760 208.765 ;
        RECT 289.270 208.455 297.060 208.765 ;
        RECT 46.790 208.225 54.760 208.455 ;
        RECT 55.080 208.260 63.060 208.455 ;
        RECT 55.080 208.225 63.040 208.260 ;
        RECT 72.790 208.225 80.760 208.455 ;
        RECT 81.080 208.260 89.060 208.455 ;
        RECT 81.080 208.225 89.040 208.260 ;
        RECT 98.790 208.225 106.760 208.455 ;
        RECT 107.080 208.260 115.060 208.455 ;
        RECT 107.080 208.225 115.040 208.260 ;
        RECT 124.790 208.225 132.760 208.455 ;
        RECT 133.080 208.260 141.060 208.455 ;
        RECT 133.080 208.225 141.040 208.260 ;
        RECT 150.790 208.225 158.760 208.455 ;
        RECT 159.080 208.260 167.060 208.455 ;
        RECT 159.080 208.225 167.040 208.260 ;
        RECT 176.790 208.225 184.760 208.455 ;
        RECT 185.080 208.260 193.060 208.455 ;
        RECT 185.080 208.225 193.040 208.260 ;
        RECT 202.790 208.225 210.760 208.455 ;
        RECT 211.080 208.260 219.060 208.455 ;
        RECT 211.080 208.225 219.040 208.260 ;
        RECT 228.790 208.225 236.760 208.455 ;
        RECT 237.080 208.260 245.060 208.455 ;
        RECT 237.080 208.225 245.040 208.260 ;
        RECT 254.790 208.225 262.760 208.455 ;
        RECT 263.080 208.260 271.060 208.455 ;
        RECT 263.080 208.225 271.040 208.260 ;
        RECT 280.790 208.225 288.760 208.455 ;
        RECT 289.080 208.260 297.060 208.455 ;
        RECT 558.080 208.320 592.150 208.810 ;
        RECT 289.080 208.225 297.040 208.260 ;
        RECT 46.970 208.220 54.760 208.225 ;
        RECT 72.970 208.220 80.760 208.225 ;
        RECT 98.970 208.220 106.760 208.225 ;
        RECT 124.970 208.220 132.760 208.225 ;
        RECT 150.970 208.220 158.760 208.225 ;
        RECT 176.970 208.220 184.760 208.225 ;
        RECT 202.970 208.220 210.760 208.225 ;
        RECT 228.970 208.220 236.760 208.225 ;
        RECT 254.970 208.220 262.760 208.225 ;
        RECT 280.970 208.220 288.760 208.225 ;
        RECT 448.030 205.240 592.150 208.320 ;
        RECT 46.970 200.880 54.660 200.910 ;
        RECT 46.970 200.815 54.760 200.880 ;
        RECT 55.190 200.815 62.980 200.910 ;
        RECT 72.970 200.880 80.660 200.910 ;
        RECT 72.970 200.815 80.760 200.880 ;
        RECT 81.190 200.815 88.980 200.910 ;
        RECT 98.970 200.880 106.660 200.910 ;
        RECT 98.970 200.815 106.760 200.880 ;
        RECT 107.190 200.815 114.980 200.910 ;
        RECT 124.970 200.880 132.660 200.910 ;
        RECT 124.970 200.815 132.760 200.880 ;
        RECT 133.190 200.815 140.980 200.910 ;
        RECT 150.970 200.880 158.660 200.910 ;
        RECT 150.970 200.815 158.760 200.880 ;
        RECT 159.190 200.815 166.980 200.910 ;
        RECT 176.970 200.880 184.660 200.910 ;
        RECT 176.970 200.815 184.760 200.880 ;
        RECT 185.190 200.815 192.980 200.910 ;
        RECT 202.970 200.880 210.660 200.910 ;
        RECT 202.970 200.815 210.760 200.880 ;
        RECT 211.190 200.815 218.980 200.910 ;
        RECT 228.970 200.880 236.660 200.910 ;
        RECT 228.970 200.815 236.760 200.880 ;
        RECT 237.190 200.815 244.980 200.910 ;
        RECT 254.970 200.880 262.660 200.910 ;
        RECT 254.970 200.815 262.760 200.880 ;
        RECT 263.190 200.815 270.980 200.910 ;
        RECT 280.970 200.880 288.660 200.910 ;
        RECT 280.970 200.815 288.760 200.880 ;
        RECT 289.190 200.815 296.980 200.910 ;
        RECT 46.790 200.585 54.760 200.815 ;
        RECT 55.080 200.585 63.040 200.815 ;
        RECT 72.790 200.585 80.760 200.815 ;
        RECT 81.080 200.585 89.040 200.815 ;
        RECT 98.790 200.585 106.760 200.815 ;
        RECT 107.080 200.585 115.040 200.815 ;
        RECT 124.790 200.585 132.760 200.815 ;
        RECT 133.080 200.585 141.040 200.815 ;
        RECT 150.790 200.585 158.760 200.815 ;
        RECT 159.080 200.585 167.040 200.815 ;
        RECT 176.790 200.585 184.760 200.815 ;
        RECT 185.080 200.585 193.040 200.815 ;
        RECT 202.790 200.585 210.760 200.815 ;
        RECT 211.080 200.585 219.040 200.815 ;
        RECT 228.790 200.585 236.760 200.815 ;
        RECT 237.080 200.585 245.040 200.815 ;
        RECT 254.790 200.585 262.760 200.815 ;
        RECT 263.080 200.585 271.040 200.815 ;
        RECT 280.790 200.585 288.760 200.815 ;
        RECT 289.080 200.585 297.040 200.815 ;
        RECT 46.970 200.275 54.760 200.585 ;
        RECT 55.190 200.275 62.980 200.585 ;
        RECT 72.970 200.275 80.760 200.585 ;
        RECT 81.190 200.275 88.980 200.585 ;
        RECT 98.970 200.275 106.760 200.585 ;
        RECT 107.190 200.275 114.980 200.585 ;
        RECT 124.970 200.275 132.760 200.585 ;
        RECT 133.190 200.275 140.980 200.585 ;
        RECT 150.970 200.275 158.760 200.585 ;
        RECT 159.190 200.275 166.980 200.585 ;
        RECT 176.970 200.275 184.760 200.585 ;
        RECT 185.190 200.275 192.980 200.585 ;
        RECT 202.970 200.275 210.760 200.585 ;
        RECT 211.190 200.275 218.980 200.585 ;
        RECT 228.970 200.275 236.760 200.585 ;
        RECT 237.190 200.275 244.980 200.585 ;
        RECT 254.970 200.275 262.760 200.585 ;
        RECT 263.190 200.275 270.980 200.585 ;
        RECT 280.970 200.275 288.760 200.585 ;
        RECT 289.190 200.275 296.980 200.585 ;
        RECT 46.790 200.120 54.760 200.275 ;
        RECT 46.790 200.045 54.750 200.120 ;
        RECT 55.080 200.045 63.040 200.275 ;
        RECT 72.790 200.120 80.760 200.275 ;
        RECT 72.790 200.045 80.750 200.120 ;
        RECT 81.080 200.045 89.040 200.275 ;
        RECT 98.790 200.120 106.760 200.275 ;
        RECT 98.790 200.045 106.750 200.120 ;
        RECT 107.080 200.045 115.040 200.275 ;
        RECT 124.790 200.120 132.760 200.275 ;
        RECT 124.790 200.045 132.750 200.120 ;
        RECT 133.080 200.045 141.040 200.275 ;
        RECT 150.790 200.120 158.760 200.275 ;
        RECT 150.790 200.045 158.750 200.120 ;
        RECT 159.080 200.045 167.040 200.275 ;
        RECT 176.790 200.120 184.760 200.275 ;
        RECT 176.790 200.045 184.750 200.120 ;
        RECT 185.080 200.045 193.040 200.275 ;
        RECT 202.790 200.120 210.760 200.275 ;
        RECT 202.790 200.045 210.750 200.120 ;
        RECT 211.080 200.045 219.040 200.275 ;
        RECT 228.790 200.120 236.760 200.275 ;
        RECT 228.790 200.045 236.750 200.120 ;
        RECT 237.080 200.045 245.040 200.275 ;
        RECT 254.790 200.120 262.760 200.275 ;
        RECT 254.790 200.045 262.750 200.120 ;
        RECT 263.080 200.045 271.040 200.275 ;
        RECT 280.790 200.120 288.760 200.275 ;
        RECT 280.790 200.045 288.750 200.120 ;
        RECT 289.080 200.045 297.040 200.275 ;
        RECT 475.070 195.000 541.600 197.460 ;
        RECT 55.170 192.700 62.860 192.730 ;
        RECT 81.170 192.700 88.860 192.730 ;
        RECT 107.170 192.700 114.860 192.730 ;
        RECT 133.170 192.700 140.860 192.730 ;
        RECT 159.170 192.700 166.860 192.730 ;
        RECT 185.170 192.700 192.860 192.730 ;
        RECT 211.170 192.700 218.860 192.730 ;
        RECT 237.170 192.700 244.860 192.730 ;
        RECT 263.170 192.700 270.860 192.730 ;
        RECT 289.170 192.700 296.860 192.730 ;
        RECT 46.890 192.635 54.680 192.690 ;
        RECT 55.070 192.635 62.860 192.700 ;
        RECT 72.890 192.635 80.680 192.690 ;
        RECT 81.070 192.635 88.860 192.700 ;
        RECT 98.890 192.635 106.680 192.690 ;
        RECT 107.070 192.635 114.860 192.700 ;
        RECT 124.890 192.635 132.680 192.690 ;
        RECT 133.070 192.635 140.860 192.700 ;
        RECT 150.890 192.635 158.680 192.690 ;
        RECT 159.070 192.635 166.860 192.700 ;
        RECT 176.890 192.635 184.680 192.690 ;
        RECT 185.070 192.635 192.860 192.700 ;
        RECT 202.890 192.635 210.680 192.690 ;
        RECT 211.070 192.635 218.860 192.700 ;
        RECT 228.890 192.635 236.680 192.690 ;
        RECT 237.070 192.635 244.860 192.700 ;
        RECT 254.890 192.635 262.680 192.690 ;
        RECT 263.070 192.635 270.860 192.700 ;
        RECT 280.890 192.635 288.680 192.690 ;
        RECT 289.070 192.635 296.860 192.700 ;
        RECT 46.790 192.405 54.750 192.635 ;
        RECT 55.070 192.405 63.040 192.635 ;
        RECT 72.790 192.405 80.750 192.635 ;
        RECT 81.070 192.405 89.040 192.635 ;
        RECT 98.790 192.405 106.750 192.635 ;
        RECT 107.070 192.405 115.040 192.635 ;
        RECT 124.790 192.405 132.750 192.635 ;
        RECT 133.070 192.405 141.040 192.635 ;
        RECT 150.790 192.405 158.750 192.635 ;
        RECT 159.070 192.405 167.040 192.635 ;
        RECT 176.790 192.405 184.750 192.635 ;
        RECT 185.070 192.405 193.040 192.635 ;
        RECT 202.790 192.405 210.750 192.635 ;
        RECT 211.070 192.405 219.040 192.635 ;
        RECT 228.790 192.405 236.750 192.635 ;
        RECT 237.070 192.405 245.040 192.635 ;
        RECT 254.790 192.405 262.750 192.635 ;
        RECT 263.070 192.405 271.040 192.635 ;
        RECT 280.790 192.405 288.750 192.635 ;
        RECT 289.070 192.405 297.040 192.635 ;
        RECT 46.890 192.095 54.680 192.405 ;
        RECT 55.070 192.095 62.860 192.405 ;
        RECT 72.890 192.095 80.680 192.405 ;
        RECT 81.070 192.095 88.860 192.405 ;
        RECT 98.890 192.095 106.680 192.405 ;
        RECT 107.070 192.095 114.860 192.405 ;
        RECT 124.890 192.095 132.680 192.405 ;
        RECT 133.070 192.095 140.860 192.405 ;
        RECT 150.890 192.095 158.680 192.405 ;
        RECT 159.070 192.095 166.860 192.405 ;
        RECT 176.890 192.095 184.680 192.405 ;
        RECT 185.070 192.095 192.860 192.405 ;
        RECT 202.890 192.095 210.680 192.405 ;
        RECT 211.070 192.095 218.860 192.405 ;
        RECT 228.890 192.095 236.680 192.405 ;
        RECT 237.070 192.095 244.860 192.405 ;
        RECT 254.890 192.095 262.680 192.405 ;
        RECT 263.070 192.095 270.860 192.405 ;
        RECT 280.890 192.095 288.680 192.405 ;
        RECT 289.070 192.095 296.860 192.405 ;
        RECT 46.790 191.865 54.750 192.095 ;
        RECT 55.070 191.940 63.040 192.095 ;
        RECT 55.080 191.865 63.040 191.940 ;
        RECT 72.790 191.865 80.750 192.095 ;
        RECT 81.070 191.940 89.040 192.095 ;
        RECT 81.080 191.865 89.040 191.940 ;
        RECT 98.790 191.865 106.750 192.095 ;
        RECT 107.070 191.940 115.040 192.095 ;
        RECT 107.080 191.865 115.040 191.940 ;
        RECT 124.790 191.865 132.750 192.095 ;
        RECT 133.070 191.940 141.040 192.095 ;
        RECT 133.080 191.865 141.040 191.940 ;
        RECT 150.790 191.865 158.750 192.095 ;
        RECT 159.070 191.940 167.040 192.095 ;
        RECT 159.080 191.865 167.040 191.940 ;
        RECT 176.790 191.865 184.750 192.095 ;
        RECT 185.070 191.940 193.040 192.095 ;
        RECT 185.080 191.865 193.040 191.940 ;
        RECT 202.790 191.865 210.750 192.095 ;
        RECT 211.070 191.940 219.040 192.095 ;
        RECT 211.080 191.865 219.040 191.940 ;
        RECT 228.790 191.865 236.750 192.095 ;
        RECT 237.070 191.940 245.040 192.095 ;
        RECT 237.080 191.865 245.040 191.940 ;
        RECT 254.790 191.865 262.750 192.095 ;
        RECT 263.070 191.940 271.040 192.095 ;
        RECT 263.080 191.865 271.040 191.940 ;
        RECT 280.790 191.865 288.750 192.095 ;
        RECT 289.070 191.940 297.040 192.095 ;
        RECT 289.080 191.865 297.040 191.940 ;
        RECT 46.970 184.455 54.760 184.510 ;
        RECT 55.150 184.455 62.940 184.510 ;
        RECT 72.970 184.455 80.760 184.510 ;
        RECT 81.150 184.455 88.940 184.510 ;
        RECT 98.970 184.455 106.760 184.510 ;
        RECT 107.150 184.455 114.940 184.510 ;
        RECT 124.970 184.455 132.760 184.510 ;
        RECT 133.150 184.455 140.940 184.510 ;
        RECT 150.970 184.455 158.760 184.510 ;
        RECT 159.150 184.455 166.940 184.510 ;
        RECT 176.970 184.455 184.760 184.510 ;
        RECT 185.150 184.455 192.940 184.510 ;
        RECT 202.970 184.455 210.760 184.510 ;
        RECT 211.150 184.455 218.940 184.510 ;
        RECT 228.970 184.455 236.760 184.510 ;
        RECT 237.150 184.455 244.940 184.510 ;
        RECT 254.970 184.455 262.760 184.510 ;
        RECT 263.150 184.455 270.940 184.510 ;
        RECT 280.970 184.455 288.760 184.510 ;
        RECT 289.150 184.455 296.940 184.510 ;
        RECT 46.790 184.225 54.760 184.455 ;
        RECT 55.080 184.225 63.040 184.455 ;
        RECT 72.790 184.225 80.760 184.455 ;
        RECT 81.080 184.225 89.040 184.455 ;
        RECT 98.790 184.225 106.760 184.455 ;
        RECT 107.080 184.225 115.040 184.455 ;
        RECT 124.790 184.225 132.760 184.455 ;
        RECT 133.080 184.225 141.040 184.455 ;
        RECT 150.790 184.225 158.760 184.455 ;
        RECT 159.080 184.225 167.040 184.455 ;
        RECT 176.790 184.225 184.760 184.455 ;
        RECT 185.080 184.225 193.040 184.455 ;
        RECT 202.790 184.225 210.760 184.455 ;
        RECT 211.080 184.225 219.040 184.455 ;
        RECT 228.790 184.225 236.760 184.455 ;
        RECT 237.080 184.225 245.040 184.455 ;
        RECT 254.790 184.225 262.760 184.455 ;
        RECT 263.080 184.225 271.040 184.455 ;
        RECT 280.790 184.225 288.760 184.455 ;
        RECT 289.080 184.225 297.040 184.455 ;
        RECT 46.970 183.915 54.760 184.225 ;
        RECT 55.150 183.915 62.940 184.225 ;
        RECT 72.970 183.915 80.760 184.225 ;
        RECT 81.150 183.915 88.940 184.225 ;
        RECT 98.970 183.915 106.760 184.225 ;
        RECT 107.150 183.915 114.940 184.225 ;
        RECT 124.970 183.915 132.760 184.225 ;
        RECT 133.150 183.915 140.940 184.225 ;
        RECT 150.970 183.915 158.760 184.225 ;
        RECT 159.150 183.915 166.940 184.225 ;
        RECT 176.970 183.915 184.760 184.225 ;
        RECT 185.150 183.915 192.940 184.225 ;
        RECT 202.970 183.915 210.760 184.225 ;
        RECT 211.150 183.915 218.940 184.225 ;
        RECT 228.970 183.915 236.760 184.225 ;
        RECT 237.150 183.915 244.940 184.225 ;
        RECT 254.970 183.915 262.760 184.225 ;
        RECT 263.150 183.915 270.940 184.225 ;
        RECT 280.970 183.915 288.760 184.225 ;
        RECT 289.150 183.915 296.940 184.225 ;
        RECT 46.790 183.720 54.760 183.915 ;
        RECT 46.790 183.685 54.750 183.720 ;
        RECT 55.080 183.685 63.040 183.915 ;
        RECT 72.790 183.720 80.760 183.915 ;
        RECT 72.790 183.685 80.750 183.720 ;
        RECT 81.080 183.685 89.040 183.915 ;
        RECT 98.790 183.720 106.760 183.915 ;
        RECT 98.790 183.685 106.750 183.720 ;
        RECT 107.080 183.685 115.040 183.915 ;
        RECT 124.790 183.720 132.760 183.915 ;
        RECT 124.790 183.685 132.750 183.720 ;
        RECT 133.080 183.685 141.040 183.915 ;
        RECT 150.790 183.720 158.760 183.915 ;
        RECT 150.790 183.685 158.750 183.720 ;
        RECT 159.080 183.685 167.040 183.915 ;
        RECT 176.790 183.720 184.760 183.915 ;
        RECT 176.790 183.685 184.750 183.720 ;
        RECT 185.080 183.685 193.040 183.915 ;
        RECT 202.790 183.720 210.760 183.915 ;
        RECT 202.790 183.685 210.750 183.720 ;
        RECT 211.080 183.685 219.040 183.915 ;
        RECT 228.790 183.720 236.760 183.915 ;
        RECT 228.790 183.685 236.750 183.720 ;
        RECT 237.080 183.685 245.040 183.915 ;
        RECT 254.790 183.720 262.760 183.915 ;
        RECT 254.790 183.685 262.750 183.720 ;
        RECT 263.080 183.685 271.040 183.915 ;
        RECT 280.790 183.720 288.760 183.915 ;
        RECT 280.790 183.685 288.750 183.720 ;
        RECT 289.080 183.685 297.040 183.915 ;
        RECT 46.850 176.275 54.640 176.330 ;
        RECT 55.190 176.275 62.980 176.330 ;
        RECT 72.850 176.275 80.640 176.330 ;
        RECT 81.190 176.275 88.980 176.330 ;
        RECT 98.850 176.275 106.640 176.330 ;
        RECT 107.190 176.275 114.980 176.330 ;
        RECT 124.850 176.275 132.640 176.330 ;
        RECT 133.190 176.275 140.980 176.330 ;
        RECT 150.850 176.275 158.640 176.330 ;
        RECT 159.190 176.275 166.980 176.330 ;
        RECT 176.850 176.275 184.640 176.330 ;
        RECT 185.190 176.275 192.980 176.330 ;
        RECT 202.850 176.275 210.640 176.330 ;
        RECT 211.190 176.275 218.980 176.330 ;
        RECT 228.850 176.275 236.640 176.330 ;
        RECT 237.190 176.275 244.980 176.330 ;
        RECT 254.850 176.275 262.640 176.330 ;
        RECT 263.190 176.275 270.980 176.330 ;
        RECT 280.850 176.275 288.640 176.330 ;
        RECT 289.190 176.275 296.980 176.330 ;
        RECT 46.790 176.045 54.750 176.275 ;
        RECT 55.080 176.045 63.040 176.275 ;
        RECT 72.790 176.045 80.750 176.275 ;
        RECT 81.080 176.045 89.040 176.275 ;
        RECT 98.790 176.045 106.750 176.275 ;
        RECT 107.080 176.045 115.040 176.275 ;
        RECT 124.790 176.045 132.750 176.275 ;
        RECT 133.080 176.045 141.040 176.275 ;
        RECT 150.790 176.045 158.750 176.275 ;
        RECT 159.080 176.045 167.040 176.275 ;
        RECT 176.790 176.045 184.750 176.275 ;
        RECT 185.080 176.045 193.040 176.275 ;
        RECT 202.790 176.045 210.750 176.275 ;
        RECT 211.080 176.045 219.040 176.275 ;
        RECT 228.790 176.045 236.750 176.275 ;
        RECT 237.080 176.045 245.040 176.275 ;
        RECT 254.790 176.045 262.750 176.275 ;
        RECT 263.080 176.045 271.040 176.275 ;
        RECT 280.790 176.045 288.750 176.275 ;
        RECT 289.080 176.045 297.040 176.275 ;
        RECT 46.850 175.735 54.640 176.045 ;
        RECT 55.190 175.735 62.980 176.045 ;
        RECT 72.850 175.735 80.640 176.045 ;
        RECT 81.190 175.735 88.980 176.045 ;
        RECT 98.850 175.735 106.640 176.045 ;
        RECT 107.190 175.735 114.980 176.045 ;
        RECT 124.850 175.735 132.640 176.045 ;
        RECT 133.190 175.735 140.980 176.045 ;
        RECT 150.850 175.735 158.640 176.045 ;
        RECT 159.190 175.735 166.980 176.045 ;
        RECT 176.850 175.735 184.640 176.045 ;
        RECT 185.190 175.735 192.980 176.045 ;
        RECT 202.850 175.735 210.640 176.045 ;
        RECT 211.190 175.735 218.980 176.045 ;
        RECT 228.850 175.735 236.640 176.045 ;
        RECT 237.190 175.735 244.980 176.045 ;
        RECT 254.850 175.735 262.640 176.045 ;
        RECT 263.190 175.735 270.980 176.045 ;
        RECT 280.850 175.735 288.640 176.045 ;
        RECT 289.190 175.735 296.980 176.045 ;
        RECT 46.790 175.505 54.750 175.735 ;
        RECT 55.080 175.505 63.040 175.735 ;
        RECT 72.790 175.505 80.750 175.735 ;
        RECT 81.080 175.505 89.040 175.735 ;
        RECT 98.790 175.505 106.750 175.735 ;
        RECT 107.080 175.505 115.040 175.735 ;
        RECT 124.790 175.505 132.750 175.735 ;
        RECT 133.080 175.505 141.040 175.735 ;
        RECT 150.790 175.505 158.750 175.735 ;
        RECT 159.080 175.505 167.040 175.735 ;
        RECT 176.790 175.505 184.750 175.735 ;
        RECT 185.080 175.505 193.040 175.735 ;
        RECT 202.790 175.505 210.750 175.735 ;
        RECT 211.080 175.505 219.040 175.735 ;
        RECT 228.790 175.505 236.750 175.735 ;
        RECT 237.080 175.505 245.040 175.735 ;
        RECT 254.790 175.505 262.750 175.735 ;
        RECT 263.080 175.505 271.040 175.735 ;
        RECT 280.790 175.505 288.750 175.735 ;
        RECT 289.080 175.505 297.040 175.735 ;
        RECT 176.590 168.150 297.120 168.160 ;
        RECT 46.780 168.110 169.920 168.120 ;
        RECT 46.780 167.240 170.060 168.110 ;
        RECT 173.520 167.350 297.120 168.150 ;
        RECT 173.520 167.330 176.660 167.350 ;
        RECT 169.710 163.180 170.060 167.240 ;
        RECT 173.530 163.180 173.890 167.330 ;
        RECT 169.690 162.930 170.060 163.180 ;
        RECT 168.360 162.690 170.060 162.930 ;
        RECT 173.520 162.930 173.920 163.180 ;
        RECT 173.520 162.690 173.930 162.930 ;
        RECT 168.360 162.260 170.050 162.690 ;
        RECT 168.360 160.610 168.740 162.260 ;
        RECT 171.960 161.100 172.270 161.270 ;
        RECT 173.550 161.100 173.930 162.690 ;
        RECT 171.960 161.060 174.200 161.100 ;
        RECT 170.530 160.860 174.200 161.060 ;
        RECT 170.540 160.840 174.200 160.860 ;
        RECT 170.540 160.700 170.690 160.840 ;
        RECT 171.770 160.820 174.200 160.840 ;
        RECT 171.770 160.800 172.280 160.820 ;
        RECT 170.530 160.690 170.690 160.700 ;
        RECT 168.330 160.460 169.690 160.610 ;
        RECT 168.330 160.430 168.740 160.460 ;
        RECT 168.330 160.130 168.710 160.430 ;
        RECT 169.550 160.260 169.690 160.460 ;
        RECT 170.530 160.260 170.680 160.690 ;
        RECT 169.070 160.250 169.300 160.260 ;
        RECT 168.440 157.350 168.690 160.130 ;
        RECT 168.870 158.260 169.300 160.250 ;
        RECT 169.550 158.260 169.780 160.260 ;
        RECT 170.030 158.260 170.260 160.260 ;
        RECT 170.510 158.260 170.740 160.260 ;
        RECT 170.990 158.270 171.470 160.260 ;
        RECT 170.990 158.260 171.370 158.270 ;
        RECT 169.050 158.030 169.230 158.260 ;
        RECT 168.850 157.860 169.230 158.030 ;
        RECT 168.850 157.640 169.260 157.860 ;
        RECT 170.030 157.650 170.210 158.260 ;
        RECT 168.850 157.520 169.880 157.640 ;
        RECT 168.930 157.490 169.880 157.520 ;
        RECT 170.030 157.510 171.000 157.650 ;
        RECT 170.030 157.500 170.460 157.510 ;
        RECT 170.030 157.490 170.260 157.500 ;
        RECT 168.440 157.210 169.400 157.350 ;
        RECT 169.260 157.040 169.400 157.210 ;
        RECT 169.740 157.040 169.880 157.490 ;
        RECT 170.820 157.040 171.000 157.510 ;
        RECT 168.830 157.020 169.060 157.040 ;
        RECT 168.660 156.060 169.060 157.020 ;
        RECT 168.830 156.040 169.060 156.060 ;
        RECT 169.260 156.040 169.540 157.040 ;
        RECT 169.740 156.060 170.020 157.040 ;
        RECT 169.790 156.040 170.020 156.060 ;
        RECT 170.270 156.110 170.500 157.040 ;
        RECT 170.750 157.020 171.000 157.040 ;
        RECT 170.270 156.040 170.530 156.110 ;
        RECT 170.750 156.070 171.160 157.020 ;
        RECT 170.750 156.040 170.980 156.070 ;
        RECT 170.330 155.680 170.530 156.040 ;
        RECT 171.970 155.700 172.280 160.800 ;
        RECT 174.360 160.360 174.890 160.870 ;
        RECT 354.670 156.010 358.460 156.030 ;
        RECT 372.150 156.010 373.300 156.140 ;
        RECT 171.950 155.690 172.290 155.700 ;
        RECT 171.780 155.680 172.290 155.690 ;
        RECT 170.330 155.450 172.290 155.680 ;
        RECT 173.020 155.500 173.540 156.010 ;
        RECT 171.780 155.430 172.290 155.450 ;
        RECT 171.780 155.420 171.980 155.430 ;
        RECT 354.670 154.540 373.300 156.010 ;
        RECT 354.670 154.500 358.850 154.540 ;
        RECT 354.670 154.490 358.460 154.500 ;
        RECT 372.150 152.870 373.300 154.540 ;
        RECT 375.000 156.010 376.470 156.020 ;
        RECT 375.000 155.990 385.960 156.010 ;
        RECT 386.190 155.990 387.060 156.010 ;
        RECT 375.000 155.970 387.060 155.990 ;
        RECT 387.800 155.970 388.730 156.010 ;
        RECT 375.000 154.540 388.800 155.970 ;
        RECT 375.000 154.530 378.030 154.540 ;
        RECT 375.000 153.900 376.470 154.530 ;
        RECT 384.720 154.450 388.800 154.540 ;
        RECT 385.790 154.340 385.960 154.450 ;
        RECT 386.190 154.340 387.060 154.450 ;
        RECT 372.150 151.790 374.380 152.870 ;
        RECT 372.250 151.730 374.380 151.790 ;
        RECT 374.930 151.450 376.470 153.900 ;
        RECT 387.800 153.730 388.730 154.450 ;
        RECT 386.010 152.840 386.950 152.910 ;
        RECT 378.150 151.820 387.020 152.840 ;
        RECT 378.150 151.790 380.460 151.820 ;
        RECT 374.980 150.290 376.390 151.450 ;
        RECT 386.010 151.170 386.950 151.820 ;
        RECT 116.690 134.070 118.090 139.790 ;
        RECT 126.770 137.530 129.810 137.590 ;
        RECT 126.750 137.130 129.810 137.530 ;
        RECT 118.950 134.340 124.890 136.660 ;
        RECT 126.750 136.130 127.180 137.130 ;
        RECT 129.540 136.660 131.300 136.690 ;
        RECT 126.730 135.720 127.180 136.130 ;
        RECT 129.530 135.800 131.300 136.660 ;
        RECT 129.530 135.760 129.760 135.800 ;
        RECT 126.730 135.550 127.170 135.720 ;
        RECT 121.310 134.330 123.020 134.340 ;
        RECT 116.040 133.490 118.090 134.070 ;
        RECT 116.010 133.330 118.090 133.490 ;
        RECT 121.490 133.330 122.400 134.330 ;
        RECT 116.010 132.750 122.400 133.330 ;
        RECT 126.770 133.180 127.170 135.550 ;
        RECT 131.050 134.950 131.300 135.800 ;
        RECT 135.040 134.950 136.720 134.960 ;
        RECT 131.020 133.290 136.720 134.950 ;
        RECT 138.590 133.670 139.990 139.350 ;
        RECT 148.670 137.090 151.710 137.150 ;
        RECT 148.650 136.690 151.710 137.090 ;
        RECT 140.850 133.900 146.790 136.220 ;
        RECT 148.650 135.280 149.080 136.690 ;
        RECT 151.440 136.220 153.200 136.250 ;
        RECT 151.430 135.360 153.200 136.220 ;
        RECT 151.430 135.320 151.660 135.360 ;
        RECT 143.210 133.890 144.920 133.900 ;
        RECT 116.010 132.710 122.380 132.750 ;
        RECT 126.750 132.720 129.760 133.180 ;
        RECT 116.010 132.680 118.090 132.710 ;
        RECT 116.010 132.650 117.290 132.680 ;
        RECT 116.010 122.410 117.120 132.650 ;
        RECT 126.750 131.210 127.210 132.720 ;
        RECT 131.050 132.560 131.300 133.290 ;
        RECT 135.040 133.270 136.720 133.290 ;
        RECT 129.440 132.540 131.300 132.560 ;
        RECT 129.430 132.250 131.300 132.540 ;
        RECT 129.430 132.220 129.710 132.250 ;
        RECT 131.050 132.220 131.300 132.250 ;
        RECT 137.420 132.890 139.990 133.670 ;
        RECT 143.390 132.890 144.300 133.890 ;
        RECT 137.420 132.310 144.300 132.890 ;
        RECT 148.670 132.740 149.070 135.280 ;
        RECT 152.950 133.870 153.200 135.360 ;
        RECT 153.760 133.870 156.920 134.050 ;
        RECT 152.940 133.400 156.920 133.870 ;
        RECT 159.380 133.640 160.780 139.120 ;
        RECT 169.460 136.860 172.500 136.920 ;
        RECT 169.440 136.460 172.500 136.860 ;
        RECT 161.640 133.670 167.580 135.990 ;
        RECT 169.440 135.520 169.870 136.460 ;
        RECT 172.230 135.990 173.990 136.020 ;
        RECT 169.320 134.870 169.970 135.520 ;
        RECT 172.220 135.130 173.990 135.990 ;
        RECT 172.220 135.090 172.450 135.130 ;
        RECT 164.000 133.660 165.710 133.670 ;
        RECT 137.420 132.270 144.280 132.310 ;
        RECT 148.650 132.280 151.660 132.740 ;
        RECT 137.420 132.240 139.990 132.270 ;
        RECT 129.200 132.010 129.480 132.070 ;
        RECT 129.200 131.780 129.490 132.010 ;
        RECT 129.200 131.750 129.480 131.780 ;
        RECT 122.520 131.180 127.210 131.210 ;
        RECT 121.390 128.810 127.210 131.180 ;
        RECT 121.390 127.080 127.190 128.810 ;
        RECT 121.400 127.040 122.200 127.080 ;
        RECT 122.520 127.070 127.190 127.080 ;
        RECT 121.630 125.090 122.240 125.550 ;
        RECT 116.010 122.290 128.840 122.410 ;
        RECT 116.010 121.390 128.920 122.290 ;
        RECT 114.460 115.230 117.110 117.050 ;
        RECT 117.450 116.440 123.250 116.950 ;
        RECT 114.460 114.900 120.420 115.230 ;
        RECT 114.410 114.690 120.420 114.900 ;
        RECT 114.380 114.580 120.420 114.690 ;
        RECT 114.380 114.540 117.610 114.580 ;
        RECT 114.380 112.830 117.400 114.540 ;
        RECT 114.380 112.600 117.610 112.830 ;
        RECT 114.380 112.510 117.400 112.600 ;
        RECT 116.060 110.940 116.380 112.510 ;
        RECT 115.860 110.560 116.460 110.940 ;
        RECT 116.060 110.360 116.380 110.560 ;
        RECT 115.850 109.920 122.780 110.060 ;
        RECT 114.590 109.550 122.780 109.920 ;
        RECT 114.630 108.960 115.310 109.550 ;
        RECT 116.160 109.270 116.390 109.280 ;
        RECT 116.090 107.670 116.390 109.270 ;
        RECT 118.240 108.580 118.880 109.410 ;
        RECT 116.900 108.065 117.940 108.295 ;
        RECT 119.190 108.065 120.230 108.295 ;
        RECT 120.710 108.100 121.010 109.310 ;
        RECT 122.840 108.580 123.480 109.410 ;
        RECT 120.710 107.740 120.990 108.100 ;
        RECT 121.480 108.065 122.520 108.295 ;
        RECT 120.650 107.670 120.990 107.740 ;
        RECT 116.090 107.420 120.990 107.670 ;
        RECT 115.520 104.655 117.560 104.885 ;
        RECT 115.410 102.660 117.910 103.270 ;
        RECT 127.930 103.210 128.920 121.390 ;
        RECT 137.420 118.920 138.940 132.240 ;
        RECT 148.650 130.770 149.110 132.280 ;
        RECT 152.950 132.120 153.200 133.400 ;
        RECT 153.760 133.120 156.920 133.400 ;
        RECT 151.340 132.100 153.200 132.120 ;
        RECT 151.330 131.810 153.200 132.100 ;
        RECT 151.330 131.780 151.610 131.810 ;
        RECT 152.950 131.780 153.200 131.810 ;
        RECT 158.110 132.660 160.780 133.640 ;
        RECT 164.180 132.660 165.090 133.660 ;
        RECT 158.110 132.080 165.090 132.660 ;
        RECT 169.460 132.510 169.860 134.870 ;
        RECT 173.740 133.640 173.990 135.130 ;
        RECT 174.660 133.640 177.820 133.880 ;
        RECT 173.730 133.170 177.820 133.640 ;
        RECT 340.880 133.310 342.750 133.420 ;
        RECT 158.110 132.040 165.070 132.080 ;
        RECT 169.440 132.050 172.450 132.510 ;
        RECT 158.110 132.010 160.780 132.040 ;
        RECT 158.110 131.980 160.180 132.010 ;
        RECT 151.100 131.570 151.380 131.630 ;
        RECT 151.100 131.340 151.390 131.570 ;
        RECT 151.100 131.310 151.380 131.340 ;
        RECT 144.420 130.740 149.110 130.770 ;
        RECT 143.290 128.370 149.110 130.740 ;
        RECT 143.290 126.640 149.090 128.370 ;
        RECT 143.300 126.600 144.100 126.640 ;
        RECT 144.420 126.630 149.090 126.640 ;
        RECT 143.530 124.650 144.140 125.110 ;
        RECT 158.110 119.380 159.710 131.980 ;
        RECT 169.440 130.540 169.900 132.050 ;
        RECT 173.740 131.890 173.990 133.170 ;
        RECT 174.660 132.950 177.820 133.170 ;
        RECT 339.260 133.090 343.400 133.310 ;
        RECT 339.260 133.055 345.200 133.090 ;
        RECT 375.020 133.055 376.370 150.290 ;
        RECT 386.090 148.850 386.910 151.170 ;
        RECT 386.240 148.840 386.890 148.850 ;
        RECT 387.800 148.790 388.680 153.730 ;
        RECT 530.570 153.030 531.910 195.000 ;
        RECT 530.340 153.020 531.910 153.030 ;
        RECT 475.090 147.940 476.140 151.010 ;
        RECT 530.340 150.300 531.320 153.020 ;
        RECT 531.550 150.290 531.910 153.020 ;
        RECT 557.920 147.990 559.370 205.240 ;
        RECT 586.510 202.910 592.150 205.240 ;
        RECT 172.130 131.870 173.990 131.890 ;
        RECT 172.120 131.580 173.990 131.870 ;
        RECT 311.510 131.690 311.880 132.030 ;
        RECT 318.320 131.850 318.700 132.180 ;
        RECT 320.320 131.930 320.640 132.410 ;
        RECT 323.350 131.930 323.750 132.250 ;
        RECT 320.320 131.750 323.750 131.930 ;
        RECT 172.120 131.550 172.400 131.580 ;
        RECT 173.740 131.550 173.990 131.580 ;
        RECT 171.890 131.340 172.170 131.400 ;
        RECT 171.890 131.110 172.180 131.340 ;
        RECT 171.890 131.080 172.170 131.110 ;
        RECT 320.320 131.050 320.640 131.750 ;
        RECT 325.200 131.730 325.580 132.050 ;
        RECT 333.990 132.020 334.370 132.440 ;
        RECT 339.260 132.375 376.370 133.055 ;
        RECT 339.260 132.180 345.200 132.375 ;
        RECT 375.020 132.350 376.370 132.375 ;
        RECT 337.270 132.170 338.580 132.180 ;
        RECT 336.990 132.020 338.650 132.170 ;
        RECT 333.990 131.420 338.650 132.020 ;
        RECT 332.010 130.980 332.420 131.400 ;
        RECT 333.990 131.070 334.370 131.420 ;
        RECT 336.990 131.200 338.650 131.420 ;
        RECT 339.260 131.970 343.400 132.180 ;
        RECT 165.210 130.510 169.900 130.540 ;
        RECT 164.080 128.140 169.900 130.510 ;
        RECT 164.080 126.410 169.880 128.140 ;
        RECT 339.260 126.780 340.210 131.970 ;
        RECT 340.880 131.750 342.750 131.970 ;
        RECT 164.090 126.370 164.890 126.410 ;
        RECT 165.210 126.400 169.880 126.410 ;
        RECT 321.460 125.680 321.930 126.160 ;
        RECT 330.160 126.110 330.500 126.560 ;
        RECT 323.300 125.600 323.720 125.960 ;
        RECT 330.060 125.680 330.520 126.110 ;
        RECT 332.100 125.730 332.460 126.310 ;
        RECT 339.260 125.780 340.250 126.780 ;
        RECT 342.690 126.480 346.530 129.000 ;
        RECT 333.260 125.730 340.250 125.780 ;
        RECT 330.160 124.930 330.500 125.680 ;
        RECT 332.100 125.470 340.250 125.730 ;
        RECT 332.100 124.970 332.460 125.470 ;
        RECT 333.260 125.450 340.250 125.470 ;
        RECT 339.260 125.050 340.250 125.450 ;
        RECT 339.280 125.040 340.250 125.050 ;
        RECT 330.160 124.920 330.470 124.930 ;
        RECT 164.320 124.420 164.930 124.880 ;
        RECT 343.010 123.510 344.980 126.480 ;
        RECT 386.330 125.400 386.760 125.420 ;
        RECT 386.330 125.250 386.810 125.400 ;
        RECT 339.590 123.220 344.980 123.510 ;
        RECT 329.760 122.230 344.980 123.220 ;
        RECT 339.590 121.710 344.980 122.230 ;
        RECT 339.590 121.680 344.370 121.710 ;
        RECT 386.340 121.630 386.810 125.250 ;
        RECT 387.890 121.990 388.420 125.420 ;
        RECT 407.560 121.990 408.970 122.790 ;
        RECT 387.890 121.770 408.970 121.990 ;
        RECT 387.890 121.740 391.190 121.770 ;
        RECT 387.890 121.720 388.420 121.740 ;
        RECT 383.140 121.590 386.810 121.630 ;
        RECT 377.800 121.330 386.810 121.590 ;
        RECT 391.340 121.520 391.550 121.530 ;
        RECT 391.340 121.370 397.400 121.520 ;
        RECT 391.340 121.360 393.750 121.370 ;
        RECT 377.810 119.530 378.210 121.330 ;
        RECT 383.140 121.320 386.750 121.330 ;
        RECT 137.420 117.200 144.490 118.920 ;
        RECT 152.520 118.280 159.710 119.380 ;
        RECT 152.500 117.660 159.710 118.280 ;
        RECT 131.360 105.435 133.400 105.665 ;
        RECT 142.280 104.930 144.370 117.200 ;
        RECT 131.370 104.025 133.480 104.060 ;
        RECT 131.360 103.795 133.480 104.025 ;
        RECT 127.930 103.200 130.770 103.210 ;
        RECT 131.370 103.200 133.480 103.795 ;
        RECT 127.930 102.790 133.480 103.200 ;
        RECT 127.930 102.750 130.770 102.790 ;
        RECT 116.700 101.200 117.335 102.660 ;
        RECT 130.085 101.215 130.710 102.750 ;
        RECT 142.280 102.700 144.370 103.640 ;
        RECT 106.280 101.060 108.240 101.090 ;
        RECT 116.700 101.060 117.340 101.200 ;
        RECT 106.280 100.380 117.340 101.060 ;
        RECT 122.870 100.440 123.300 100.920 ;
        RECT 130.065 100.495 130.710 101.215 ;
        RECT 143.360 101.030 143.995 102.700 ;
        RECT 152.500 101.760 154.050 117.660 ;
        RECT 158.110 117.640 159.710 117.660 ;
        RECT 377.820 109.640 378.210 119.530 ;
        RECT 378.620 119.240 383.170 119.270 ;
        RECT 386.210 119.240 386.670 119.260 ;
        RECT 378.620 119.020 386.670 119.240 ;
        RECT 378.620 118.930 384.180 119.020 ;
        RECT 385.340 118.930 386.670 119.020 ;
        RECT 378.620 118.920 383.170 118.930 ;
        RECT 378.620 118.840 381.800 118.920 ;
        RECT 377.800 109.010 378.210 109.640 ;
        RECT 234.210 105.830 236.460 107.890 ;
        RECT 255.660 107.380 257.930 107.910 ;
        RECT 255.650 104.220 257.930 106.300 ;
        RECT 260.200 104.250 262.470 104.720 ;
        RECT 281.610 104.200 283.900 107.890 ;
        RECT 106.280 93.560 108.240 100.380 ;
        RECT 110.635 100.180 111.435 100.185 ;
        RECT 116.700 100.180 117.330 100.380 ;
        RECT 122.885 100.180 123.685 100.185 ;
        RECT 110.635 99.685 123.685 100.180 ;
        RECT 110.635 98.540 111.435 99.685 ;
        RECT 122.885 98.540 123.685 99.685 ;
        RECT 110.635 97.585 123.685 98.540 ;
        RECT 110.635 96.490 111.435 97.585 ;
        RECT 122.885 96.490 123.685 97.585 ;
        RECT 110.635 95.535 123.685 96.490 ;
        RECT 110.635 94.340 111.435 95.535 ;
        RECT 122.885 94.340 123.685 95.535 ;
        RECT 110.635 93.385 123.685 94.340 ;
        RECT 110.635 92.290 111.435 93.385 ;
        RECT 122.885 92.290 123.685 93.385 ;
        RECT 110.635 91.335 123.685 92.290 ;
        RECT 110.635 90.190 111.435 91.335 ;
        RECT 122.885 90.190 123.685 91.335 ;
        RECT 110.635 89.235 123.685 90.190 ;
        RECT 110.635 88.140 111.435 89.235 ;
        RECT 122.885 88.140 123.685 89.235 ;
        RECT 110.635 87.185 123.685 88.140 ;
        RECT 110.635 86.035 111.435 87.185 ;
        RECT 122.885 86.035 123.685 87.185 ;
        RECT 110.635 85.385 123.685 86.035 ;
        RECT 123.985 100.180 124.785 100.185 ;
        RECT 130.080 100.180 130.710 100.495 ;
        RECT 135.480 100.370 136.090 100.890 ;
        RECT 143.360 100.495 144.060 101.030 ;
        RECT 145.640 100.500 146.210 101.000 ;
        RECT 137.300 100.185 138.100 100.190 ;
        RECT 143.360 100.185 143.990 100.495 ;
        RECT 149.570 100.490 154.050 101.760 ;
        RECT 152.500 100.460 154.050 100.490 ;
        RECT 149.550 100.185 150.350 100.190 ;
        RECT 136.235 100.180 137.035 100.185 ;
        RECT 123.985 99.685 137.035 100.180 ;
        RECT 123.985 98.540 124.785 99.685 ;
        RECT 136.235 98.540 137.035 99.685 ;
        RECT 123.985 97.585 137.035 98.540 ;
        RECT 123.985 96.490 124.785 97.585 ;
        RECT 136.235 96.490 137.035 97.585 ;
        RECT 123.985 95.535 137.035 96.490 ;
        RECT 123.985 94.340 124.785 95.535 ;
        RECT 136.235 94.340 137.035 95.535 ;
        RECT 123.985 93.385 137.035 94.340 ;
        RECT 123.985 92.290 124.785 93.385 ;
        RECT 136.235 92.290 137.035 93.385 ;
        RECT 123.985 91.335 137.035 92.290 ;
        RECT 123.985 90.190 124.785 91.335 ;
        RECT 136.235 90.190 137.035 91.335 ;
        RECT 123.985 89.235 137.035 90.190 ;
        RECT 123.985 88.140 124.785 89.235 ;
        RECT 136.235 88.140 137.035 89.235 ;
        RECT 123.985 87.185 137.035 88.140 ;
        RECT 123.985 86.035 124.785 87.185 ;
        RECT 136.235 86.035 137.035 87.185 ;
        RECT 123.985 85.385 137.035 86.035 ;
        RECT 137.300 99.690 150.350 100.185 ;
        RECT 137.300 98.545 138.100 99.690 ;
        RECT 149.550 98.545 150.350 99.690 ;
        RECT 234.240 99.460 236.480 99.920 ;
        RECT 255.620 99.450 257.900 103.150 ;
        RECT 260.210 101.060 262.440 103.120 ;
        RECT 281.650 102.660 283.890 103.110 ;
        RECT 281.650 99.470 283.880 101.530 ;
        RECT 137.300 97.590 150.350 98.545 ;
        RECT 137.300 96.495 138.100 97.590 ;
        RECT 149.550 96.495 150.350 97.590 ;
        RECT 234.210 98.300 236.460 98.340 ;
        RECT 137.300 95.540 150.350 96.495 ;
        RECT 137.300 94.345 138.100 95.540 ;
        RECT 149.550 94.345 150.350 95.540 ;
        RECT 137.300 93.390 150.350 94.345 ;
        RECT 137.300 92.295 138.100 93.390 ;
        RECT 149.550 92.295 150.350 93.390 ;
        RECT 137.300 91.340 150.350 92.295 ;
        RECT 137.300 90.195 138.100 91.340 ;
        RECT 149.550 90.195 150.350 91.340 ;
        RECT 137.300 89.240 150.350 90.195 ;
        RECT 137.300 88.145 138.100 89.240 ;
        RECT 149.550 88.145 150.350 89.240 ;
        RECT 137.300 87.190 150.350 88.145 ;
        RECT 137.300 86.040 138.100 87.190 ;
        RECT 149.550 86.040 150.350 87.190 ;
        RECT 137.300 85.390 150.350 86.040 ;
        RECT 116.220 84.270 118.140 85.385 ;
        RECT 130.190 84.990 132.110 85.385 ;
        RECT 130.200 84.620 132.110 84.990 ;
        RECT 116.220 83.800 116.970 84.270 ;
        RECT 130.190 83.840 132.110 84.620 ;
        RECT 143.210 84.200 145.130 85.390 ;
        RECT 143.210 83.830 144.410 84.200 ;
        RECT 117.120 83.140 117.620 83.700 ;
        RECT 131.790 83.270 132.190 83.670 ;
        RECT 144.280 83.190 146.510 83.690 ;
        RECT 116.410 82.830 116.950 83.060 ;
        RECT 131.070 82.870 131.610 83.100 ;
        RECT 143.630 82.870 144.170 83.100 ;
        RECT 20.030 80.900 21.150 80.950 ;
        RECT 20.030 79.650 39.440 80.900 ;
        RECT 20.030 71.260 21.150 79.650 ;
        RECT 24.760 74.160 25.690 75.130 ;
        RECT 18.700 71.060 19.720 71.230 ;
        RECT 24.840 71.060 25.530 74.160 ;
        RECT 18.700 70.390 25.530 71.060 ;
        RECT 18.700 70.270 19.720 70.390 ;
        RECT 24.840 70.370 25.530 70.390 ;
        RECT 22.390 69.600 23.130 69.760 ;
        RECT 21.130 69.210 27.470 69.600 ;
        RECT 21.150 64.680 21.480 69.210 ;
        RECT 22.390 68.960 23.130 69.210 ;
        RECT 27.210 69.190 27.450 69.210 ;
        RECT 29.530 69.200 29.770 69.550 ;
        RECT 24.670 67.030 25.410 67.150 ;
        RECT 24.670 66.640 27.540 67.030 ;
        RECT 29.560 66.670 29.800 67.020 ;
        RECT 24.670 66.350 25.410 66.640 ;
        RECT 24.860 64.800 25.270 66.350 ;
        RECT 21.140 63.580 21.490 64.680 ;
        RECT 21.150 61.640 21.480 63.580 ;
        RECT 24.850 63.470 25.270 64.800 ;
        RECT 27.020 63.990 27.520 64.490 ;
        RECT 29.550 64.080 29.790 64.430 ;
        RECT 38.300 64.070 39.400 79.650 ;
        RECT 152.820 77.720 153.960 96.990 ;
        RECT 234.210 96.330 236.470 98.300 ;
        RECT 260.220 97.880 262.490 98.350 ;
        RECT 234.210 96.280 236.460 96.330 ;
        RECT 255.670 94.690 257.910 95.160 ;
        RECT 260.200 94.660 262.470 96.790 ;
        RECT 377.800 96.420 378.170 109.010 ;
        RECT 377.800 96.220 378.190 96.420 ;
        RECT 226.990 89.580 227.830 90.290 ;
        RECT 227.290 87.300 227.490 89.580 ;
        RECT 243.900 88.750 244.950 89.680 ;
        RECT 226.870 86.440 227.940 87.300 ;
        RECT 244.240 84.790 244.440 88.750 ;
        RECT 245.530 88.550 245.910 89.250 ;
        RECT 246.410 88.590 246.840 89.250 ;
        RECT 250.050 88.590 250.550 89.340 ;
        RECT 258.930 88.620 259.520 89.510 ;
        RECT 246.910 87.650 248.070 87.830 ;
        RECT 256.850 87.650 257.840 87.770 ;
        RECT 246.910 87.450 257.840 87.650 ;
        RECT 271.260 87.560 271.800 88.140 ;
        RECT 278.420 87.640 278.910 88.020 ;
        RECT 279.770 87.690 280.030 87.950 ;
        RECT 281.320 87.910 281.810 88.390 ;
        RECT 246.910 87.350 248.070 87.450 ;
        RECT 244.640 87.090 245.340 87.320 ;
        RECT 253.540 87.090 254.470 87.310 ;
        RECT 244.640 86.850 254.470 87.090 ;
        RECT 256.850 86.880 257.840 87.450 ;
        RECT 279.780 86.860 280.020 87.690 ;
        RECT 244.640 86.840 247.350 86.850 ;
        RECT 244.640 86.700 245.340 86.840 ;
        RECT 253.540 86.620 254.470 86.850 ;
        RECT 259.630 86.440 260.210 86.640 ;
        RECT 251.600 86.410 260.210 86.440 ;
        RECT 260.960 86.410 261.490 86.510 ;
        RECT 251.600 86.210 261.490 86.410 ;
        RECT 275.320 86.320 280.070 86.860 ;
        RECT 281.440 86.780 281.640 87.910 ;
        RECT 288.550 87.650 289.840 87.830 ;
        RECT 288.550 87.460 298.750 87.650 ;
        RECT 288.550 87.330 289.840 87.460 ;
        RECT 289.100 86.850 289.950 87.170 ;
        RECT 251.600 86.190 260.210 86.210 ;
        RECT 251.610 85.850 251.800 86.190 ;
        RECT 250.700 85.835 251.800 85.850 ;
        RECT 250.680 85.605 251.800 85.835 ;
        RECT 259.630 85.680 260.210 86.190 ;
        RECT 260.960 86.160 261.490 86.210 ;
        RECT 261.790 85.690 262.320 85.750 ;
        RECT 261.460 85.680 262.390 85.690 ;
        RECT 250.700 85.600 251.800 85.605 ;
        RECT 259.590 85.440 262.390 85.680 ;
        RECT 261.460 85.370 262.390 85.440 ;
        RECT 261.790 85.230 262.320 85.370 ;
        RECT 275.390 84.980 275.980 86.320 ;
        RECT 279.780 85.140 280.020 86.320 ;
        RECT 281.240 85.780 281.810 86.780 ;
        RECT 279.220 84.840 283.220 85.140 ;
        RECT 238.840 84.690 239.490 84.750 ;
        RECT 243.120 84.690 243.590 84.770 ;
        RECT 238.840 84.450 243.590 84.690 ;
        RECT 238.840 84.310 239.490 84.450 ;
        RECT 243.120 84.370 243.590 84.450 ;
        RECT 244.230 84.330 244.450 84.790 ;
        RECT 244.890 84.690 245.360 84.770 ;
        RECT 244.890 84.450 264.600 84.690 ;
        RECT 244.890 84.370 245.360 84.450 ;
        RECT 213.400 83.320 216.340 83.330 ;
        RECT 213.400 83.150 218.720 83.320 ;
        RECT 213.400 83.130 216.340 83.150 ;
        RECT 213.400 82.320 213.670 83.130 ;
        RECT 216.090 83.120 216.340 83.130 ;
        RECT 212.290 80.310 213.010 82.320 ;
        RECT 213.240 82.310 213.670 82.320 ;
        RECT 213.220 80.320 213.670 82.310 ;
        RECT 213.950 82.810 215.790 82.980 ;
        RECT 213.950 82.300 214.110 82.810 ;
        RECT 215.540 82.800 215.790 82.810 ;
        RECT 215.590 82.320 215.790 82.800 ;
        RECT 213.220 80.310 213.490 80.320 ;
        RECT 212.730 79.780 212.950 80.310 ;
        RECT 213.940 80.300 214.170 82.300 ;
        RECT 214.360 80.300 214.720 82.300 ;
        RECT 213.970 79.800 214.110 80.300 ;
        RECT 214.860 80.290 215.310 82.320 ;
        RECT 215.590 82.290 215.900 82.320 ;
        RECT 216.140 82.300 216.340 83.120 ;
        RECT 216.620 82.300 217.000 82.310 ;
        RECT 216.140 82.290 216.400 82.300 ;
        RECT 215.520 82.280 215.900 82.290 ;
        RECT 215.480 81.470 215.900 82.280 ;
        RECT 215.520 81.130 215.900 81.470 ;
        RECT 215.480 80.300 215.900 81.130 ;
        RECT 216.170 80.300 216.400 82.290 ;
        RECT 216.610 80.300 217.000 82.300 ;
        RECT 212.730 79.640 213.670 79.780 ;
        RECT 213.970 79.660 214.750 79.800 ;
        RECT 213.530 79.120 213.670 79.640 ;
        RECT 214.570 79.140 214.750 79.660 ;
        RECT 215.040 79.790 215.230 80.290 ;
        RECT 215.480 80.280 215.860 80.300 ;
        RECT 215.040 79.650 215.830 79.790 ;
        RECT 214.570 79.130 214.990 79.140 ;
        RECT 215.650 79.130 215.830 79.650 ;
        RECT 216.170 79.780 216.340 80.300 ;
        RECT 216.170 79.640 216.970 79.780 ;
        RECT 213.980 79.120 214.210 79.130 ;
        RECT 212.900 79.070 213.130 79.120 ;
        RECT 212.710 78.130 213.130 79.070 ;
        RECT 212.900 78.120 213.130 78.130 ;
        RECT 213.340 78.130 214.210 79.120 ;
        RECT 214.420 79.120 215.300 79.130 ;
        RECT 215.510 79.120 216.180 79.130 ;
        RECT 216.770 79.120 216.970 79.640 ;
        RECT 214.420 78.150 215.310 79.120 ;
        RECT 214.420 78.140 215.300 78.150 ;
        RECT 214.420 78.130 214.650 78.140 ;
        RECT 214.980 78.130 215.300 78.140 ;
        RECT 215.510 78.140 216.410 79.120 ;
        RECT 215.510 78.130 215.740 78.140 ;
        RECT 213.340 78.120 214.140 78.130 ;
        RECT 214.980 78.120 215.180 78.130 ;
        RECT 216.180 78.120 216.410 78.140 ;
        RECT 216.620 78.150 217.010 79.120 ;
        RECT 216.620 78.120 216.850 78.150 ;
        RECT 214.540 77.980 214.800 77.990 ;
        RECT 218.540 77.980 218.720 83.150 ;
        RECT 239.330 83.220 242.270 83.420 ;
        RECT 239.330 82.410 239.600 83.220 ;
        RECT 242.020 83.210 242.270 83.220 ;
        RECT 238.220 80.400 238.940 82.410 ;
        RECT 239.170 82.400 239.600 82.410 ;
        RECT 239.150 80.410 239.600 82.400 ;
        RECT 239.880 82.900 241.720 83.070 ;
        RECT 239.880 82.390 240.040 82.900 ;
        RECT 241.470 82.890 241.720 82.900 ;
        RECT 241.520 82.410 241.720 82.890 ;
        RECT 239.150 80.400 239.420 80.410 ;
        RECT 238.660 79.870 238.880 80.400 ;
        RECT 239.870 80.390 240.100 82.390 ;
        RECT 240.290 80.390 240.650 82.390 ;
        RECT 239.900 79.890 240.040 80.390 ;
        RECT 240.790 80.380 241.240 82.410 ;
        RECT 241.520 82.380 241.830 82.410 ;
        RECT 242.070 82.390 242.270 83.210 ;
        RECT 242.550 82.390 242.930 82.400 ;
        RECT 242.070 82.380 242.330 82.390 ;
        RECT 241.450 82.370 241.830 82.380 ;
        RECT 241.410 81.560 241.830 82.370 ;
        RECT 241.450 81.220 241.830 81.560 ;
        RECT 241.410 80.390 241.830 81.220 ;
        RECT 242.100 80.390 242.330 82.380 ;
        RECT 242.540 82.070 242.930 82.390 ;
        RECT 244.240 82.090 244.440 84.330 ;
        RECT 251.490 84.180 251.750 84.210 ;
        RECT 244.240 82.070 246.830 82.090 ;
        RECT 242.540 81.870 246.830 82.070 ;
        RECT 242.540 81.850 244.440 81.870 ;
        RECT 242.540 80.390 242.930 81.850 ;
        RECT 238.660 79.730 239.600 79.870 ;
        RECT 239.900 79.750 240.680 79.890 ;
        RECT 239.460 79.210 239.600 79.730 ;
        RECT 240.500 79.230 240.680 79.750 ;
        RECT 240.970 79.880 241.160 80.380 ;
        RECT 241.410 80.370 241.790 80.390 ;
        RECT 240.970 79.740 241.760 79.880 ;
        RECT 240.500 79.220 240.920 79.230 ;
        RECT 241.580 79.220 241.760 79.740 ;
        RECT 242.100 79.870 242.270 80.390 ;
        RECT 246.610 79.920 246.810 81.870 ;
        RECT 250.190 81.620 250.420 84.180 ;
        RECT 251.480 81.620 251.750 84.180 ;
        RECT 252.450 83.700 255.585 84.240 ;
        RECT 246.610 79.890 248.290 79.920 ;
        RECT 251.490 79.890 251.750 81.620 ;
        RECT 252.455 81.450 255.585 83.700 ;
        RECT 255.745 81.460 258.875 84.250 ;
        RECT 264.290 84.120 264.600 84.450 ;
        RECT 259.160 81.490 259.390 84.050 ;
        RECT 260.450 81.490 260.680 84.050 ;
        RECT 264.290 83.990 264.950 84.120 ;
        RECT 274.040 83.990 274.280 84.010 ;
        RECT 262.110 83.440 262.990 83.740 ;
        RECT 264.290 83.710 274.280 83.990 ;
        RECT 264.290 83.590 264.950 83.710 ;
        RECT 265.210 83.440 268.150 83.480 ;
        RECT 262.110 83.280 268.150 83.440 ;
        RECT 262.110 83.230 265.480 83.280 ;
        RECT 267.900 83.270 268.150 83.280 ;
        RECT 262.110 82.990 262.990 83.230 ;
        RECT 265.210 82.470 265.480 83.230 ;
        RECT 264.100 80.460 264.820 82.470 ;
        RECT 265.050 82.460 265.480 82.470 ;
        RECT 265.030 80.470 265.480 82.460 ;
        RECT 265.760 82.960 267.600 83.130 ;
        RECT 265.760 82.450 265.920 82.960 ;
        RECT 267.350 82.950 267.600 82.960 ;
        RECT 267.400 82.470 267.600 82.950 ;
        RECT 265.030 80.460 265.300 80.470 ;
        RECT 242.100 79.730 242.900 79.870 ;
        RECT 242.700 79.560 242.900 79.730 ;
        RECT 246.610 79.720 251.750 79.890 ;
        RECT 246.640 79.700 251.750 79.720 ;
        RECT 247.540 79.690 251.750 79.700 ;
        RECT 244.680 79.560 244.940 79.570 ;
        RECT 242.700 79.330 244.940 79.560 ;
        RECT 239.910 79.210 240.140 79.220 ;
        RECT 238.830 79.160 239.060 79.210 ;
        RECT 225.590 77.980 226.910 78.560 ;
        RECT 238.640 78.220 239.060 79.160 ;
        RECT 238.830 78.210 239.060 78.220 ;
        RECT 239.270 78.220 240.140 79.210 ;
        RECT 240.350 79.210 241.230 79.220 ;
        RECT 241.440 79.210 242.110 79.220 ;
        RECT 242.700 79.210 242.940 79.330 ;
        RECT 240.350 78.240 241.240 79.210 ;
        RECT 240.350 78.230 241.230 78.240 ;
        RECT 240.350 78.220 240.580 78.230 ;
        RECT 240.910 78.220 241.230 78.230 ;
        RECT 241.440 78.230 242.340 79.210 ;
        RECT 241.440 78.220 241.670 78.230 ;
        RECT 239.270 78.210 240.070 78.220 ;
        RECT 240.910 78.210 241.110 78.220 ;
        RECT 242.110 78.210 242.340 78.230 ;
        RECT 242.550 78.240 242.940 79.210 ;
        RECT 244.680 78.740 244.940 79.330 ;
        RECT 247.060 79.370 247.850 79.490 ;
        RECT 253.520 79.370 254.530 80.040 ;
        RECT 263.340 79.940 263.920 80.070 ;
        RECT 264.540 79.940 264.760 80.460 ;
        RECT 265.750 80.450 265.980 82.450 ;
        RECT 266.170 80.450 266.530 82.450 ;
        RECT 263.340 79.930 264.760 79.940 ;
        RECT 265.780 79.950 265.920 80.450 ;
        RECT 266.670 80.440 267.120 82.470 ;
        RECT 267.400 82.440 267.710 82.470 ;
        RECT 267.950 82.450 268.150 83.270 ;
        RECT 268.430 82.450 268.810 82.460 ;
        RECT 267.950 82.440 268.210 82.450 ;
        RECT 267.330 82.430 267.710 82.440 ;
        RECT 267.290 81.620 267.710 82.430 ;
        RECT 267.330 81.280 267.710 81.620 ;
        RECT 267.290 80.450 267.710 81.280 ;
        RECT 267.980 80.450 268.210 82.440 ;
        RECT 268.420 82.380 268.810 82.450 ;
        RECT 268.420 82.150 270.590 82.380 ;
        RECT 268.420 80.450 268.810 82.150 ;
        RECT 263.340 79.790 265.480 79.930 ;
        RECT 265.780 79.810 266.560 79.950 ;
        RECT 263.340 79.770 264.700 79.790 ;
        RECT 263.340 79.560 263.920 79.770 ;
        RECT 247.060 79.320 254.530 79.370 ;
        RECT 247.060 79.210 254.110 79.320 ;
        RECT 265.340 79.270 265.480 79.790 ;
        RECT 266.380 79.290 266.560 79.810 ;
        RECT 266.850 79.940 267.040 80.440 ;
        RECT 267.290 80.430 267.670 80.450 ;
        RECT 266.850 79.800 267.640 79.940 ;
        RECT 266.380 79.280 266.800 79.290 ;
        RECT 267.460 79.280 267.640 79.800 ;
        RECT 267.980 79.930 268.150 80.450 ;
        RECT 267.980 79.790 268.780 79.930 ;
        RECT 265.790 79.270 266.020 79.280 ;
        RECT 264.710 79.220 264.940 79.270 ;
        RECT 247.060 79.090 247.850 79.210 ;
        RECT 258.380 78.740 258.700 79.030 ;
        RECT 244.670 78.560 258.700 78.740 ;
        RECT 258.380 78.520 258.700 78.560 ;
        RECT 259.880 78.270 261.220 78.600 ;
        RECT 264.520 78.280 264.940 79.220 ;
        RECT 264.710 78.270 264.940 78.280 ;
        RECT 265.150 78.280 266.020 79.270 ;
        RECT 266.230 79.270 267.110 79.280 ;
        RECT 267.320 79.270 267.990 79.280 ;
        RECT 268.580 79.270 268.780 79.790 ;
        RECT 266.230 78.300 267.120 79.270 ;
        RECT 266.230 78.290 267.110 78.300 ;
        RECT 266.230 78.280 266.460 78.290 ;
        RECT 266.790 78.280 267.110 78.290 ;
        RECT 267.320 78.290 268.220 79.270 ;
        RECT 267.320 78.280 267.550 78.290 ;
        RECT 265.150 78.270 265.950 78.280 ;
        RECT 266.790 78.270 266.990 78.280 ;
        RECT 267.990 78.270 268.220 78.290 ;
        RECT 268.430 78.300 268.820 79.270 ;
        RECT 268.430 78.270 268.660 78.300 ;
        RECT 247.360 78.260 261.220 78.270 ;
        RECT 242.550 78.210 242.780 78.240 ;
        RECT 214.420 77.750 216.190 77.980 ;
        RECT 218.540 77.750 226.910 77.980 ;
        RECT 214.540 77.740 214.800 77.750 ;
        RECT 215.910 77.720 216.190 77.750 ;
        RECT 115.890 76.685 117.930 76.915 ;
        RECT 129.600 76.805 131.640 77.035 ;
        RECT 142.780 76.845 144.820 77.075 ;
        RECT 134.330 75.730 135.070 76.330 ;
        RECT 44.460 71.650 44.980 72.240 ;
        RECT 47.110 71.270 47.720 71.830 ;
        RECT 47.130 71.260 47.720 71.270 ;
        RECT 45.730 70.460 47.410 70.520 ;
        RECT 45.730 70.290 47.920 70.460 ;
        RECT 45.730 70.230 47.410 70.290 ;
        RECT 46.830 70.220 47.410 70.230 ;
        RECT 43.650 69.700 44.430 70.030 ;
        RECT 44.020 69.440 44.210 69.700 ;
        RECT 45.910 69.440 47.620 69.490 ;
        RECT 47.760 69.440 47.920 70.290 ;
        RECT 44.020 69.430 47.920 69.440 ;
        RECT 43.950 69.260 47.920 69.430 ;
        RECT 43.950 69.230 44.290 69.260 ;
        RECT 45.910 69.240 47.920 69.260 ;
        RECT 45.910 69.210 47.620 69.240 ;
        RECT 47.760 69.230 47.920 69.240 ;
        RECT 47.010 68.200 47.620 68.760 ;
        RECT 68.800 68.670 70.200 74.560 ;
        RECT 115.840 74.190 118.120 75.330 ;
        RECT 118.890 74.360 120.320 75.430 ;
        RECT 129.390 74.420 131.670 75.560 ;
        RECT 142.520 75.435 144.800 75.540 ;
        RECT 145.560 75.480 146.310 76.550 ;
        RECT 152.800 76.450 153.960 77.720 ;
        RECT 225.590 77.310 226.910 77.750 ;
        RECT 236.540 77.190 237.240 77.430 ;
        RECT 239.600 77.190 239.800 78.210 ;
        RECT 240.470 78.070 240.730 78.080 ;
        RECT 240.350 77.840 242.120 78.070 ;
        RECT 240.470 77.830 240.730 77.840 ;
        RECT 241.840 77.810 242.120 77.840 ;
        RECT 247.290 78.020 261.220 78.260 ;
        RECT 266.350 78.130 266.610 78.140 ;
        RECT 218.390 76.450 218.990 76.630 ;
        RECT 230.620 76.450 231.940 77.140 ;
        RECT 236.540 77.090 239.820 77.190 ;
        RECT 247.290 77.090 247.560 78.020 ;
        RECT 259.880 77.650 261.220 78.020 ;
        RECT 266.230 77.900 268.000 78.130 ;
        RECT 266.350 77.890 266.610 77.900 ;
        RECT 267.720 77.870 268.000 77.900 ;
        RECT 236.540 76.900 247.560 77.090 ;
        RECT 236.540 76.790 237.240 76.900 ;
        RECT 239.360 76.880 247.490 76.900 ;
        RECT 239.600 76.870 239.800 76.880 ;
        RECT 218.390 76.220 231.940 76.450 ;
        RECT 218.390 76.050 218.990 76.220 ;
        RECT 230.620 75.890 231.940 76.220 ;
        RECT 240.730 75.910 241.390 76.480 ;
        RECT 211.910 75.500 212.510 75.630 ;
        RECT 237.970 75.500 238.550 75.620 ;
        RECT 142.520 75.205 144.820 75.435 ;
        RECT 211.910 75.260 238.550 75.500 ;
        RECT 78.880 72.300 81.920 72.360 ;
        RECT 78.860 71.900 81.920 72.300 ;
        RECT 71.060 69.110 77.000 71.430 ;
        RECT 78.860 70.490 79.290 71.900 ;
        RECT 106.510 71.840 111.630 72.940 ;
        RECT 116.700 72.660 117.330 74.190 ;
        RECT 130.080 72.660 130.710 74.420 ;
        RECT 142.520 74.400 144.800 75.205 ;
        RECT 211.910 75.090 212.510 75.260 ;
        RECT 237.970 75.150 238.550 75.260 ;
        RECT 210.660 74.600 211.470 75.070 ;
        RECT 237.530 74.600 238.010 74.670 ;
        RECT 106.510 71.460 107.690 71.840 ;
        RECT 116.700 71.800 124.940 72.660 ;
        RECT 130.080 72.445 137.860 72.660 ;
        RECT 130.065 71.910 137.860 72.445 ;
        RECT 110.635 71.595 111.435 71.600 ;
        RECT 116.700 71.595 117.330 71.800 ;
        RECT 130.080 71.780 137.860 71.910 ;
        RECT 143.360 72.610 143.990 74.400 ;
        RECT 210.660 74.310 238.010 74.600 ;
        RECT 152.820 72.610 153.960 72.950 ;
        RECT 143.360 71.910 153.960 72.610 ;
        RECT 143.360 71.900 152.810 71.910 ;
        RECT 122.885 71.595 123.685 71.600 ;
        RECT 110.635 71.590 122.170 71.595 ;
        RECT 122.450 71.590 123.685 71.595 ;
        RECT 81.650 71.430 83.410 71.460 ;
        RECT 81.640 70.570 83.410 71.430 ;
        RECT 81.640 70.530 81.870 70.570 ;
        RECT 73.420 69.100 75.130 69.110 ;
        RECT 68.120 68.530 70.200 68.670 ;
        RECT 68.120 68.100 71.720 68.530 ;
        RECT 73.600 68.100 74.510 69.100 ;
        RECT 68.120 67.520 74.510 68.100 ;
        RECT 78.880 67.950 79.280 70.490 ;
        RECT 83.160 69.080 83.410 70.570 ;
        RECT 110.635 71.100 123.685 71.590 ;
        RECT 110.635 69.955 111.435 71.100 ;
        RECT 122.885 69.955 123.685 71.100 ;
        RECT 84.130 69.080 86.500 69.120 ;
        RECT 83.150 68.610 86.500 69.080 ;
        RECT 110.635 69.000 123.685 69.955 ;
        RECT 68.120 67.480 74.490 67.520 ;
        RECT 78.860 67.490 81.870 67.950 ;
        RECT 45.770 67.400 47.450 67.460 ;
        RECT 45.770 67.230 47.960 67.400 ;
        RECT 45.770 67.170 47.450 67.230 ;
        RECT 46.870 67.160 47.450 67.170 ;
        RECT 43.710 66.650 44.460 66.960 ;
        RECT 44.060 66.380 44.250 66.650 ;
        RECT 45.950 66.380 47.660 66.430 ;
        RECT 47.800 66.380 47.960 67.230 ;
        RECT 44.060 66.340 47.960 66.380 ;
        RECT 43.970 66.200 47.960 66.340 ;
        RECT 43.970 66.140 44.310 66.200 ;
        RECT 45.950 66.180 47.960 66.200 ;
        RECT 45.950 66.150 47.660 66.180 ;
        RECT 47.800 66.170 47.960 66.180 ;
        RECT 68.120 67.360 71.720 67.480 ;
        RECT 47.030 65.300 47.640 65.860 ;
        RECT 45.750 64.510 47.430 64.570 ;
        RECT 45.750 64.340 47.940 64.510 ;
        RECT 45.750 64.280 47.430 64.340 ;
        RECT 46.850 64.270 47.430 64.280 ;
        RECT 38.300 64.050 44.440 64.070 ;
        RECT 38.300 63.790 44.480 64.050 ;
        RECT 38.850 63.780 44.480 63.790 ;
        RECT 39.700 63.760 44.480 63.780 ;
        RECT 43.700 63.750 44.440 63.760 ;
        RECT 24.860 61.830 25.270 63.470 ;
        RECT 44.040 63.490 44.230 63.750 ;
        RECT 45.930 63.490 47.640 63.540 ;
        RECT 47.780 63.490 47.940 64.340 ;
        RECT 44.040 63.450 47.940 63.490 ;
        RECT 43.960 63.310 47.940 63.450 ;
        RECT 43.960 63.250 44.300 63.310 ;
        RECT 45.930 63.290 47.940 63.310 ;
        RECT 45.930 63.260 47.640 63.290 ;
        RECT 47.780 63.280 47.940 63.290 ;
        RECT 47.060 62.430 47.670 62.990 ;
        RECT 25.820 61.970 26.620 62.220 ;
        RECT 21.150 61.030 21.470 61.640 ;
        RECT 21.150 60.840 21.480 61.030 ;
        RECT 24.870 60.580 25.270 61.830 ;
        RECT 25.440 61.520 27.470 61.970 ;
        RECT 29.550 61.530 29.790 61.880 ;
        RECT 45.790 61.640 47.470 61.700 ;
        RECT 25.440 61.470 27.460 61.520 ;
        RECT 45.790 61.470 47.980 61.640 ;
        RECT 24.930 60.430 25.270 60.580 ;
        RECT 25.450 61.380 26.620 61.470 ;
        RECT 45.790 61.410 47.470 61.470 ;
        RECT 46.890 61.400 47.470 61.410 ;
        RECT 20.820 59.920 21.410 60.350 ;
        RECT 20.950 59.900 21.410 59.920 ;
        RECT 25.450 59.910 25.870 61.380 ;
        RECT 43.740 61.170 44.490 61.200 ;
        RECT 43.740 60.950 44.500 61.170 ;
        RECT 43.740 60.890 44.490 60.950 ;
        RECT 44.080 60.620 44.270 60.890 ;
        RECT 45.970 60.620 47.680 60.670 ;
        RECT 47.820 60.620 47.980 61.470 ;
        RECT 44.080 60.600 47.980 60.620 ;
        RECT 44.040 60.590 47.980 60.600 ;
        RECT 43.990 60.440 47.980 60.590 ;
        RECT 43.990 60.390 44.330 60.440 ;
        RECT 45.970 60.420 47.980 60.440 ;
        RECT 45.970 60.390 47.680 60.420 ;
        RECT 47.820 60.410 47.980 60.420 ;
        RECT 24.920 59.530 25.870 59.910 ;
        RECT 47.050 59.540 47.660 60.100 ;
        RECT 24.950 59.510 25.870 59.530 ;
        RECT 21.130 59.360 21.430 59.410 ;
        RECT 21.100 58.960 27.510 59.360 ;
        RECT 29.550 58.980 29.790 59.330 ;
        RECT 21.130 58.920 21.430 58.960 ;
        RECT 24.910 58.800 25.440 58.820 ;
        RECT 21.140 58.000 21.500 58.450 ;
        RECT 24.910 58.430 25.900 58.800 ;
        RECT 21.130 57.130 21.460 57.460 ;
        RECT 21.130 57.080 21.430 57.130 ;
        RECT 21.150 56.680 21.430 57.080 ;
        RECT 21.150 54.270 21.460 56.680 ;
        RECT 24.950 54.380 25.260 57.950 ;
        RECT 25.570 56.900 25.900 58.430 ;
        RECT 39.680 58.450 40.890 58.760 ;
        RECT 45.790 58.750 47.470 58.810 ;
        RECT 45.790 58.580 47.980 58.750 ;
        RECT 45.790 58.520 47.470 58.580 ;
        RECT 46.890 58.510 47.470 58.520 ;
        RECT 39.680 58.370 41.480 58.450 ;
        RECT 39.680 58.330 42.090 58.370 ;
        RECT 39.680 58.310 43.480 58.330 ;
        RECT 39.680 58.270 44.480 58.310 ;
        RECT 39.680 58.040 44.500 58.270 ;
        RECT 39.680 58.000 44.480 58.040 ;
        RECT 39.680 57.980 41.480 58.000 ;
        RECT 39.680 57.430 40.890 57.980 ;
        RECT 44.070 57.730 44.270 58.000 ;
        RECT 45.970 57.730 47.680 57.780 ;
        RECT 47.820 57.730 47.980 58.580 ;
        RECT 68.120 58.360 69.030 67.360 ;
        RECT 78.860 65.980 79.320 67.490 ;
        RECT 83.160 67.330 83.410 68.610 ;
        RECT 81.550 67.310 83.410 67.330 ;
        RECT 81.540 67.020 83.410 67.310 ;
        RECT 81.540 66.990 81.820 67.020 ;
        RECT 83.160 66.990 83.410 67.020 ;
        RECT 81.310 66.780 81.590 66.840 ;
        RECT 81.310 66.550 81.600 66.780 ;
        RECT 81.310 66.520 81.590 66.550 ;
        RECT 74.630 65.950 79.320 65.980 ;
        RECT 73.500 63.580 79.320 65.950 ;
        RECT 73.500 61.850 79.300 63.580 ;
        RECT 73.510 61.810 74.310 61.850 ;
        RECT 74.630 61.840 79.300 61.850 ;
        RECT 73.740 59.860 74.350 60.320 ;
        RECT 44.070 57.570 47.980 57.730 ;
        RECT 44.080 57.550 47.980 57.570 ;
        RECT 45.970 57.530 47.980 57.550 ;
        RECT 45.970 57.500 47.680 57.530 ;
        RECT 47.820 57.520 47.980 57.530 ;
        RECT 25.570 56.790 26.520 56.900 ;
        RECT 25.570 56.410 27.520 56.790 ;
        RECT 29.550 56.430 29.790 56.780 ;
        RECT 47.040 56.650 47.650 57.210 ;
        RECT 25.590 56.400 27.520 56.410 ;
        RECT 25.590 55.880 26.520 56.400 ;
        RECT 45.790 55.860 47.470 55.920 ;
        RECT 39.240 55.350 40.280 55.730 ;
        RECT 45.790 55.690 47.980 55.860 ;
        RECT 45.790 55.630 47.470 55.690 ;
        RECT 46.890 55.620 47.470 55.630 ;
        RECT 43.740 55.390 44.480 55.420 ;
        RECT 40.960 55.350 44.500 55.390 ;
        RECT 39.240 55.100 44.500 55.350 ;
        RECT 39.240 55.080 41.550 55.100 ;
        RECT 39.240 54.530 40.280 55.080 ;
        RECT 44.080 54.840 44.270 55.100 ;
        RECT 45.970 54.840 47.680 54.890 ;
        RECT 47.820 54.840 47.980 55.690 ;
        RECT 44.080 54.660 47.980 54.840 ;
        RECT 45.970 54.640 47.980 54.660 ;
        RECT 45.970 54.610 47.680 54.640 ;
        RECT 47.820 54.630 47.980 54.640 ;
        RECT 67.950 55.510 69.090 58.360 ;
        RECT 21.140 53.790 21.470 54.270 ;
        RECT 21.150 52.140 21.460 53.790 ;
        RECT 21.130 49.150 21.460 52.140 ;
        RECT 24.950 53.670 25.250 54.380 ;
        RECT 27.030 54.300 27.490 54.310 ;
        RECT 27.030 53.800 27.520 54.300 ;
        RECT 29.550 53.880 29.790 54.230 ;
        RECT 27.030 53.790 27.490 53.800 ;
        RECT 47.150 53.730 47.760 54.290 ;
        RECT 67.950 54.050 86.220 55.510 ;
        RECT 24.950 51.980 25.260 53.670 ;
        RECT 45.810 52.950 47.490 53.010 ;
        RECT 39.310 52.460 40.410 52.910 ;
        RECT 45.810 52.780 48.000 52.950 ;
        RECT 45.810 52.720 47.490 52.780 ;
        RECT 46.910 52.710 47.490 52.720 ;
        RECT 43.760 52.460 44.500 52.510 ;
        RECT 39.310 52.170 44.560 52.460 ;
        RECT 24.860 51.860 25.680 51.980 ;
        RECT 24.780 51.720 25.680 51.860 ;
        RECT 24.780 51.300 27.490 51.720 ;
        RECT 29.550 51.330 29.790 51.680 ;
        RECT 39.310 51.560 40.410 52.170 ;
        RECT 44.100 51.930 44.290 52.170 ;
        RECT 45.990 51.930 47.700 51.980 ;
        RECT 47.840 51.930 48.000 52.780 ;
        RECT 44.100 51.890 48.000 51.930 ;
        RECT 44.060 51.750 48.000 51.890 ;
        RECT 44.060 51.720 44.350 51.750 ;
        RECT 45.990 51.730 48.000 51.750 ;
        RECT 45.990 51.700 47.700 51.730 ;
        RECT 47.840 51.720 48.000 51.730 ;
        RECT 24.780 51.280 25.680 51.300 ;
        RECT 24.860 51.210 25.680 51.280 ;
        RECT 47.130 50.860 47.740 51.420 ;
        RECT 68.060 50.630 85.900 51.710 ;
        RECT 45.790 50.070 47.470 50.130 ;
        RECT 45.790 49.900 47.980 50.070 ;
        RECT 45.790 49.840 47.470 49.900 ;
        RECT 46.890 49.830 47.470 49.840 ;
        RECT 39.650 49.620 41.440 49.740 ;
        RECT 43.740 49.620 44.480 49.630 ;
        RECT 25.950 49.150 26.840 49.450 ;
        RECT 39.650 49.340 44.500 49.620 ;
        RECT 39.650 49.230 41.440 49.340 ;
        RECT 43.740 49.320 44.480 49.340 ;
        RECT 21.090 48.760 27.520 49.150 ;
        RECT 29.550 48.780 29.790 49.130 ;
        RECT 21.130 48.730 21.460 48.760 ;
        RECT 25.950 48.550 26.840 48.760 ;
        RECT 24.760 45.870 25.640 46.790 ;
        RECT 24.890 45.740 25.640 45.870 ;
        RECT 32.860 45.740 34.570 45.770 ;
        RECT 39.650 45.740 40.500 49.230 ;
        RECT 44.080 49.050 44.270 49.320 ;
        RECT 45.970 49.050 47.680 49.100 ;
        RECT 47.820 49.050 47.980 49.900 ;
        RECT 44.080 49.020 47.980 49.050 ;
        RECT 44.060 48.870 47.980 49.020 ;
        RECT 44.060 48.850 44.350 48.870 ;
        RECT 45.970 48.850 47.980 48.870 ;
        RECT 45.970 48.820 47.680 48.850 ;
        RECT 47.820 48.840 47.980 48.850 ;
        RECT 69.090 48.810 70.430 50.630 ;
        RECT 43.370 48.350 43.840 48.800 ;
        RECT 69.090 48.320 70.590 48.810 ;
        RECT 45.770 47.220 47.450 47.280 ;
        RECT 45.770 47.050 47.960 47.220 ;
        RECT 45.770 46.990 47.450 47.050 ;
        RECT 46.870 46.980 47.450 46.990 ;
        RECT 43.710 46.470 44.470 46.790 ;
        RECT 44.060 46.200 44.250 46.470 ;
        RECT 45.950 46.200 47.660 46.250 ;
        RECT 47.800 46.200 47.960 47.050 ;
        RECT 44.060 46.020 47.960 46.200 ;
        RECT 44.060 45.980 44.350 46.020 ;
        RECT 45.950 46.000 47.960 46.020 ;
        RECT 45.950 45.970 47.660 46.000 ;
        RECT 47.800 45.990 47.960 46.000 ;
        RECT 24.890 45.690 25.940 45.740 ;
        RECT 32.860 45.690 40.500 45.740 ;
        RECT 24.890 45.160 40.500 45.690 ;
        RECT 24.900 44.920 40.500 45.160 ;
        RECT 24.900 44.880 40.240 44.920 ;
        RECT 24.900 44.870 33.480 44.880 ;
        RECT 25.760 44.850 33.480 44.870 ;
        RECT 69.190 42.350 70.590 48.320 ;
        RECT 79.270 46.550 82.310 46.610 ;
        RECT 106.550 46.550 107.690 67.960 ;
        RECT 110.635 67.905 111.435 69.000 ;
        RECT 122.885 67.905 123.685 69.000 ;
        RECT 110.635 66.950 123.685 67.905 ;
        RECT 110.635 65.755 111.435 66.950 ;
        RECT 122.885 65.755 123.685 66.950 ;
        RECT 110.635 64.800 123.685 65.755 ;
        RECT 110.635 63.705 111.435 64.800 ;
        RECT 122.885 63.705 123.685 64.800 ;
        RECT 110.635 62.750 123.685 63.705 ;
        RECT 110.635 61.605 111.435 62.750 ;
        RECT 122.885 61.605 123.685 62.750 ;
        RECT 110.635 60.650 123.685 61.605 ;
        RECT 110.635 59.555 111.435 60.650 ;
        RECT 122.885 59.555 123.685 60.650 ;
        RECT 110.635 58.600 123.685 59.555 ;
        RECT 110.635 57.450 111.435 58.600 ;
        RECT 122.885 57.450 123.685 58.600 ;
        RECT 110.635 56.820 123.685 57.450 ;
        RECT 110.635 56.800 117.120 56.820 ;
        RECT 117.480 56.800 123.685 56.820 ;
        RECT 123.985 71.595 124.785 71.600 ;
        RECT 130.080 71.595 130.710 71.780 ;
        RECT 137.300 71.600 138.100 71.605 ;
        RECT 143.360 71.600 143.990 71.900 ;
        RECT 235.190 71.720 238.170 72.160 ;
        RECT 149.550 71.600 150.350 71.605 ;
        RECT 136.235 71.595 137.035 71.600 ;
        RECT 123.985 71.590 135.540 71.595 ;
        RECT 135.810 71.590 137.035 71.595 ;
        RECT 123.985 71.100 137.035 71.590 ;
        RECT 123.985 69.955 124.785 71.100 ;
        RECT 136.235 69.955 137.035 71.100 ;
        RECT 123.985 69.000 137.035 69.955 ;
        RECT 123.985 67.905 124.785 69.000 ;
        RECT 136.235 67.905 137.035 69.000 ;
        RECT 123.985 66.950 137.035 67.905 ;
        RECT 123.985 65.755 124.785 66.950 ;
        RECT 136.235 65.755 137.035 66.950 ;
        RECT 123.985 64.800 137.035 65.755 ;
        RECT 123.985 63.705 124.785 64.800 ;
        RECT 136.235 63.705 137.035 64.800 ;
        RECT 123.985 62.750 137.035 63.705 ;
        RECT 123.985 61.605 124.785 62.750 ;
        RECT 136.235 61.605 137.035 62.750 ;
        RECT 123.985 60.650 137.035 61.605 ;
        RECT 123.985 59.555 124.785 60.650 ;
        RECT 136.235 59.555 137.035 60.650 ;
        RECT 123.985 58.600 137.035 59.555 ;
        RECT 123.985 57.450 124.785 58.600 ;
        RECT 136.235 57.450 137.035 58.600 ;
        RECT 123.985 56.800 137.035 57.450 ;
        RECT 137.300 71.105 150.350 71.600 ;
        RECT 137.300 69.960 138.100 71.105 ;
        RECT 149.550 69.960 150.350 71.105 ;
        RECT 227.620 71.500 238.170 71.720 ;
        RECT 227.620 70.260 227.850 71.500 ;
        RECT 235.190 71.140 238.170 71.500 ;
        RECT 137.300 69.005 150.350 69.960 ;
        RECT 224.110 69.900 231.140 70.260 ;
        RECT 137.300 67.910 138.100 69.005 ;
        RECT 149.550 67.910 150.350 69.005 ;
        RECT 137.300 66.955 150.350 67.910 ;
        RECT 137.300 65.760 138.100 66.955 ;
        RECT 149.550 65.760 150.350 66.955 ;
        RECT 240.870 66.260 241.210 75.910 ;
        RECT 249.875 75.115 255.610 76.275 ;
        RECT 259.890 76.270 261.180 77.130 ;
        RECT 265.650 76.550 266.320 77.200 ;
        RECT 256.080 76.220 261.180 76.270 ;
        RECT 256.080 75.115 260.680 76.220 ;
        RECT 261.000 75.610 261.880 76.050 ;
        RECT 251.160 70.840 255.610 75.115 ;
        RECT 256.230 70.840 260.680 75.115 ;
        RECT 265.750 73.440 266.200 76.550 ;
        RECT 265.750 73.200 266.220 73.440 ;
        RECT 265.760 72.340 266.220 73.200 ;
        RECT 250.060 69.700 251.850 70.020 ;
        RECT 251.620 67.030 251.850 69.700 ;
        RECT 255.380 70.010 256.300 70.260 ;
        RECT 261.010 70.010 261.740 70.160 ;
        RECT 255.380 69.780 261.740 70.010 ;
        RECT 255.380 69.270 256.300 69.780 ;
        RECT 261.010 69.740 261.740 69.780 ;
        RECT 262.020 69.710 262.970 69.990 ;
        RECT 270.380 69.710 270.590 82.150 ;
        RECT 274.040 77.930 274.280 83.710 ;
        RECT 289.750 78.940 289.930 86.850 ;
        RECT 295.140 82.880 295.820 83.420 ;
        RECT 290.630 82.430 291.320 82.790 ;
        RECT 293.490 82.430 296.430 82.440 ;
        RECT 290.630 82.240 296.430 82.430 ;
        RECT 290.630 82.010 291.320 82.240 ;
        RECT 293.490 81.430 293.760 82.240 ;
        RECT 296.180 82.230 296.430 82.240 ;
        RECT 292.380 79.420 293.100 81.430 ;
        RECT 293.330 81.420 293.760 81.430 ;
        RECT 293.310 79.430 293.760 81.420 ;
        RECT 294.040 81.920 295.880 82.090 ;
        RECT 294.040 81.410 294.200 81.920 ;
        RECT 295.630 81.910 295.880 81.920 ;
        RECT 295.680 81.430 295.880 81.910 ;
        RECT 293.310 79.420 293.580 79.430 ;
        RECT 292.820 78.940 293.040 79.420 ;
        RECT 294.030 79.410 294.260 81.410 ;
        RECT 294.450 79.410 294.810 81.410 ;
        RECT 289.750 78.890 293.040 78.940 ;
        RECT 294.060 78.910 294.200 79.410 ;
        RECT 294.950 79.400 295.400 81.430 ;
        RECT 295.680 81.400 295.990 81.430 ;
        RECT 296.230 81.410 296.430 82.230 ;
        RECT 296.710 81.410 297.090 81.420 ;
        RECT 296.230 81.400 296.490 81.410 ;
        RECT 295.610 81.390 295.990 81.400 ;
        RECT 295.570 80.580 295.990 81.390 ;
        RECT 295.610 80.240 295.990 80.580 ;
        RECT 295.570 79.410 295.990 80.240 ;
        RECT 296.260 79.410 296.490 81.400 ;
        RECT 296.700 81.350 297.090 81.410 ;
        RECT 298.510 81.350 298.700 87.460 ;
        RECT 377.820 83.520 378.190 96.220 ;
        RECT 377.820 83.000 378.220 83.520 ;
        RECT 296.700 81.160 298.700 81.350 ;
        RECT 296.700 79.410 297.090 81.160 ;
        RECT 298.510 81.100 298.700 81.160 ;
        RECT 289.750 78.760 293.760 78.890 ;
        RECT 294.060 78.770 294.840 78.910 ;
        RECT 292.820 78.750 293.760 78.760 ;
        RECT 293.620 78.230 293.760 78.750 ;
        RECT 294.660 78.250 294.840 78.770 ;
        RECT 295.130 78.900 295.320 79.400 ;
        RECT 295.570 79.390 295.950 79.410 ;
        RECT 295.130 78.760 295.920 78.900 ;
        RECT 294.660 78.240 295.080 78.250 ;
        RECT 295.740 78.240 295.920 78.760 ;
        RECT 296.260 78.890 296.430 79.410 ;
        RECT 296.260 78.750 297.060 78.890 ;
        RECT 294.070 78.230 294.300 78.240 ;
        RECT 292.990 78.180 293.220 78.230 ;
        RECT 287.250 77.930 287.840 78.000 ;
        RECT 274.040 77.650 287.840 77.930 ;
        RECT 287.250 77.550 287.840 77.650 ;
        RECT 270.850 77.010 271.220 77.190 ;
        RECT 291.330 77.020 291.840 77.250 ;
        RECT 292.800 77.240 293.220 78.180 ;
        RECT 292.990 77.230 293.220 77.240 ;
        RECT 293.430 77.240 294.300 78.230 ;
        RECT 294.510 78.230 295.390 78.240 ;
        RECT 295.600 78.230 296.270 78.240 ;
        RECT 296.860 78.230 297.060 78.750 ;
        RECT 294.510 77.260 295.400 78.230 ;
        RECT 294.510 77.250 295.390 77.260 ;
        RECT 294.510 77.240 294.740 77.250 ;
        RECT 295.070 77.240 295.390 77.250 ;
        RECT 295.600 77.250 296.500 78.230 ;
        RECT 295.600 77.240 295.830 77.250 ;
        RECT 293.430 77.230 294.230 77.240 ;
        RECT 295.070 77.230 295.270 77.240 ;
        RECT 296.270 77.230 296.500 77.250 ;
        RECT 296.710 77.260 297.100 78.230 ;
        RECT 296.710 77.230 296.940 77.260 ;
        RECT 294.630 77.090 294.890 77.100 ;
        RECT 280.870 77.010 291.840 77.020 ;
        RECT 270.850 76.780 291.840 77.010 ;
        RECT 294.510 76.860 296.280 77.090 ;
        RECT 294.630 76.850 294.890 76.860 ;
        RECT 296.000 76.830 296.280 76.860 ;
        RECT 270.850 76.770 281.030 76.780 ;
        RECT 290.580 76.770 291.840 76.780 ;
        RECT 270.850 76.630 271.220 76.770 ;
        RECT 291.330 76.760 291.840 76.770 ;
        RECT 304.700 76.410 305.300 76.780 ;
        RECT 271.690 74.500 272.980 74.700 ;
        RECT 271.690 74.280 283.080 74.500 ;
        RECT 271.690 74.130 272.980 74.280 ;
        RECT 270.780 73.960 271.320 74.100 ;
        RECT 270.780 73.940 274.050 73.960 ;
        RECT 270.780 73.730 278.150 73.940 ;
        RECT 270.780 73.690 274.050 73.730 ;
        RECT 270.780 73.430 271.320 73.690 ;
        RECT 277.960 72.600 278.150 73.730 ;
        RECT 277.110 72.470 278.150 72.600 ;
        RECT 282.870 72.490 283.080 74.280 ;
        RECT 282.130 72.470 283.080 72.490 ;
        RECT 277.110 72.130 280.390 72.470 ;
        RECT 282.130 72.130 285.400 72.470 ;
        RECT 262.020 69.500 270.650 69.710 ;
        RECT 262.020 69.290 262.970 69.500 ;
        RECT 265.580 69.490 266.620 69.500 ;
        RECT 251.610 67.020 253.730 67.030 ;
        RECT 251.610 66.710 258.920 67.020 ;
        RECT 252.970 66.690 258.920 66.710 ;
        RECT 253.580 66.660 258.920 66.690 ;
        RECT 240.870 66.250 256.590 66.260 ;
        RECT 265.750 66.250 266.200 68.980 ;
        RECT 268.800 67.440 269.940 68.470 ;
        RECT 277.110 67.720 278.000 72.130 ;
        RECT 277.110 67.380 280.400 67.720 ;
        RECT 282.130 67.700 283.020 72.130 ;
        RECT 377.850 70.660 378.220 83.000 ;
        RECT 377.820 70.100 378.220 70.660 ;
        RECT 240.870 65.990 266.230 66.250 ;
        RECT 240.880 65.970 266.230 65.990 ;
        RECT 250.520 65.960 266.230 65.970 ;
        RECT 137.300 64.805 150.350 65.760 ;
        RECT 137.300 63.710 138.100 64.805 ;
        RECT 149.550 63.710 150.350 64.805 ;
        RECT 137.300 62.755 150.350 63.710 ;
        RECT 137.300 61.610 138.100 62.755 ;
        RECT 149.550 61.610 150.350 62.755 ;
        RECT 277.110 62.950 278.000 67.380 ;
        RECT 282.130 67.360 285.400 67.700 ;
        RECT 277.110 62.610 280.410 62.950 ;
        RECT 282.130 62.930 283.020 67.360 ;
        RECT 277.110 62.480 278.000 62.610 ;
        RECT 282.130 62.590 285.400 62.930 ;
        RECT 282.130 62.370 283.020 62.590 ;
        RECT 137.300 60.655 150.350 61.610 ;
        RECT 137.300 59.560 138.100 60.655 ;
        RECT 149.550 59.560 150.350 60.655 ;
        RECT 137.300 58.605 150.350 59.560 ;
        RECT 137.300 57.455 138.100 58.605 ;
        RECT 149.550 57.455 150.350 58.605 ;
        RECT 137.300 56.805 150.350 57.455 ;
        RECT 116.290 55.800 117.120 56.800 ;
        RECT 116.290 55.270 116.960 55.800 ;
        RECT 130.050 55.480 131.290 56.800 ;
        RECT 116.320 55.260 116.860 55.270 ;
        RECT 116.320 54.290 116.860 54.520 ;
        RECT 117.020 54.480 117.500 55.140 ;
        RECT 130.050 54.920 131.170 55.480 ;
        RECT 142.690 55.180 143.190 56.805 ;
        RECT 143.550 56.800 144.100 56.805 ;
        RECT 184.990 55.410 186.390 58.410 ;
        RECT 377.820 57.240 378.190 70.100 ;
        RECT 378.640 57.920 379.170 118.840 ;
        RECT 386.210 116.600 386.670 118.930 ;
        RECT 387.800 119.200 388.280 119.210 ;
        RECT 391.340 119.200 391.550 121.360 ;
        RECT 396.010 119.590 397.400 121.370 ;
        RECT 407.560 120.780 408.970 121.770 ;
        RECT 387.800 119.030 391.730 119.200 ;
        RECT 387.800 119.000 389.410 119.030 ;
        RECT 390.320 119.000 391.730 119.030 ;
        RECT 387.800 116.610 388.280 119.000 ;
        RECT 380.410 95.310 386.790 95.340 ;
        RECT 380.410 94.750 386.840 95.310 ;
        RECT 380.460 91.780 381.890 94.750 ;
        RECT 386.160 90.730 386.840 94.750 ;
        RECT 387.640 93.160 388.480 93.170 ;
        RECT 386.260 90.710 386.660 90.730 ;
        RECT 382.000 89.650 382.930 89.700 ;
        RECT 382.000 89.470 383.410 89.650 ;
        RECT 386.260 89.570 386.660 89.640 ;
        RECT 387.610 89.570 388.530 93.160 ;
        RECT 386.260 89.470 388.530 89.570 ;
        RECT 382.000 89.210 388.530 89.470 ;
        RECT 382.000 89.200 386.690 89.210 ;
        RECT 387.610 89.200 388.530 89.210 ;
        RECT 382.000 88.920 383.410 89.200 ;
        RECT 382.000 88.000 382.930 88.920 ;
        RECT 382.000 87.070 382.870 88.000 ;
        RECT 382.000 86.970 382.860 87.070 ;
        RECT 380.030 74.180 381.090 74.570 ;
        RECT 381.970 74.180 382.860 86.970 ;
        RECT 380.030 73.710 382.860 74.180 ;
        RECT 380.030 73.200 381.090 73.710 ;
        RECT 381.970 73.580 382.860 73.710 ;
        RECT 454.830 69.630 457.670 109.980 ;
        RECT 482.630 82.440 485.800 110.250 ;
        RECT 512.290 109.870 515.910 110.180 ;
        RECT 510.540 109.810 515.910 109.870 ;
        RECT 510.500 108.080 515.910 109.810 ;
        RECT 521.120 109.260 525.010 110.640 ;
        RECT 538.080 110.190 541.590 110.530 ;
        RECT 482.270 82.190 486.990 82.440 ;
        RECT 482.180 81.740 489.520 82.190 ;
        RECT 481.720 76.710 489.520 81.740 ;
        RECT 510.500 77.710 514.190 108.080 ;
        RECT 510.620 77.140 514.170 77.710 ;
        RECT 481.720 76.470 487.350 76.710 ;
        RECT 454.710 60.530 457.750 69.630 ;
        RECT 378.640 57.370 379.180 57.920 ;
        RECT 195.070 56.150 198.110 56.210 ;
        RECT 142.690 54.950 143.250 55.180 ;
        RECT 130.600 54.000 131.140 54.230 ;
        RECT 131.310 54.170 131.840 54.890 ;
        RECT 143.410 54.280 143.950 54.920 ;
        RECT 142.710 53.980 143.250 54.210 ;
        RECT 179.490 53.970 186.390 55.410 ;
        RECT 195.050 55.750 198.110 56.150 ;
        RECT 184.990 51.950 186.390 53.970 ;
        RECT 187.250 52.960 193.190 55.280 ;
        RECT 195.050 54.340 195.480 55.750 ;
        RECT 197.840 55.280 199.600 55.310 ;
        RECT 197.830 54.420 199.600 55.280 ;
        RECT 293.970 55.170 296.640 57.220 ;
        RECT 197.830 54.380 198.060 54.420 ;
        RECT 189.610 52.950 191.320 52.960 ;
        RECT 189.790 51.950 190.700 52.950 ;
        RECT 184.990 51.370 190.700 51.950 ;
        RECT 195.070 51.800 195.470 54.340 ;
        RECT 199.350 52.930 199.600 54.420 ;
        RECT 293.940 53.380 304.270 55.170 ;
        RECT 293.970 53.110 296.640 53.380 ;
        RECT 200.520 52.930 204.470 52.940 ;
        RECT 199.340 52.460 204.470 52.930 ;
        RECT 184.990 51.330 190.680 51.370 ;
        RECT 195.050 51.340 198.060 51.800 ;
        RECT 184.990 51.300 186.390 51.330 ;
        RECT 195.050 49.830 195.510 51.340 ;
        RECT 199.350 51.180 199.600 52.460 ;
        RECT 197.740 51.160 199.600 51.180 ;
        RECT 197.730 50.870 199.600 51.160 ;
        RECT 197.730 50.840 198.010 50.870 ;
        RECT 199.350 50.840 199.600 50.870 ;
        RECT 197.500 50.630 197.780 50.690 ;
        RECT 197.500 50.400 197.790 50.630 ;
        RECT 197.500 50.370 197.780 50.400 ;
        RECT 190.820 49.800 195.510 49.830 ;
        RECT 129.870 47.455 131.910 47.685 ;
        RECT 116.170 47.215 118.210 47.445 ;
        RECT 142.550 47.225 144.590 47.455 ;
        RECT 189.690 47.430 195.510 49.800 ;
        RECT 79.250 46.150 82.310 46.550 ;
        RECT 71.450 43.360 77.390 45.680 ;
        RECT 79.250 45.320 79.680 46.150 ;
        RECT 82.040 45.680 83.800 45.710 ;
        RECT 79.110 44.480 79.690 45.320 ;
        RECT 82.030 44.820 83.800 45.680 ;
        RECT 116.060 45.390 118.450 46.020 ;
        RECT 118.880 45.880 119.860 46.980 ;
        RECT 129.640 45.390 132.070 46.320 ;
        RECT 132.770 46.040 133.750 47.140 ;
        RECT 145.390 46.060 146.370 47.160 ;
        RECT 116.060 44.950 118.490 45.390 ;
        RECT 129.330 45.050 132.070 45.390 ;
        RECT 129.640 45.040 132.070 45.050 ;
        RECT 82.030 44.780 82.260 44.820 ;
        RECT 73.810 43.350 75.520 43.360 ;
        RECT 73.990 42.350 74.900 43.350 ;
        RECT 69.190 41.770 74.900 42.350 ;
        RECT 79.270 42.200 79.670 44.480 ;
        RECT 83.550 43.330 83.800 44.820 ;
        RECT 116.290 44.710 118.490 44.950 ;
        RECT 116.705 43.440 117.335 44.710 ;
        RECT 84.250 43.330 86.620 43.350 ;
        RECT 83.540 42.860 86.620 43.330 ;
        RECT 69.190 41.730 74.880 41.770 ;
        RECT 79.250 41.740 82.260 42.200 ;
        RECT 69.190 41.700 70.590 41.730 ;
        RECT 79.250 40.230 79.710 41.740 ;
        RECT 83.550 41.580 83.800 42.860 ;
        RECT 84.250 42.840 86.620 42.860 ;
        RECT 106.550 43.225 117.335 43.440 ;
        RECT 130.085 43.235 130.715 45.040 ;
        RECT 142.470 44.690 144.900 45.970 ;
        RECT 189.690 45.700 195.490 47.430 ;
        RECT 189.700 45.660 190.500 45.700 ;
        RECT 190.820 45.690 195.490 45.700 ;
        RECT 106.550 42.390 117.330 43.225 ;
        RECT 130.080 43.135 130.715 43.235 ;
        RECT 130.080 42.925 130.710 43.135 ;
        RECT 130.065 42.390 130.710 42.925 ;
        RECT 110.630 42.075 111.460 42.090 ;
        RECT 116.700 42.075 117.330 42.390 ;
        RECT 122.885 42.075 123.685 42.080 ;
        RECT 110.630 41.585 123.685 42.075 ;
        RECT 81.940 41.560 83.800 41.580 ;
        RECT 81.930 41.270 83.800 41.560 ;
        RECT 81.930 41.240 82.210 41.270 ;
        RECT 83.550 41.240 83.800 41.270 ;
        RECT 110.635 41.580 123.685 41.585 ;
        RECT 81.700 41.030 81.980 41.090 ;
        RECT 81.700 40.800 81.990 41.030 ;
        RECT 81.700 40.770 81.980 40.800 ;
        RECT 75.020 40.200 79.710 40.230 ;
        RECT 73.890 37.830 79.710 40.200 ;
        RECT 110.635 40.435 111.435 41.580 ;
        RECT 122.885 40.435 123.685 41.580 ;
        RECT 110.635 39.480 123.685 40.435 ;
        RECT 110.635 38.385 111.435 39.480 ;
        RECT 122.885 38.385 123.685 39.480 ;
        RECT 73.890 36.100 79.690 37.830 ;
        RECT 73.900 36.060 74.700 36.100 ;
        RECT 75.020 36.090 79.690 36.100 ;
        RECT 110.635 37.430 123.685 38.385 ;
        RECT 110.635 36.235 111.435 37.430 ;
        RECT 122.885 36.235 123.685 37.430 ;
        RECT 110.635 35.280 123.685 36.235 ;
        RECT 74.130 34.110 74.740 34.570 ;
        RECT 110.635 34.185 111.435 35.280 ;
        RECT 122.885 34.185 123.685 35.280 ;
        RECT 110.635 33.230 123.685 34.185 ;
        RECT 110.635 32.085 111.435 33.230 ;
        RECT 122.885 32.085 123.685 33.230 ;
        RECT 110.635 31.130 123.685 32.085 ;
        RECT 110.635 30.035 111.435 31.130 ;
        RECT 122.885 30.035 123.685 31.130 ;
        RECT 110.635 29.080 123.685 30.035 ;
        RECT 110.635 27.930 111.435 29.080 ;
        RECT 122.885 27.930 123.685 29.080 ;
        RECT 110.635 27.280 123.685 27.930 ;
        RECT 123.985 42.075 124.785 42.080 ;
        RECT 130.080 42.075 130.710 42.390 ;
        RECT 143.360 43.105 143.995 44.690 ;
        RECT 149.600 44.340 150.210 44.400 ;
        RECT 143.360 42.925 143.990 43.105 ;
        RECT 143.360 42.390 144.060 42.925 ;
        RECT 137.300 42.080 138.100 42.085 ;
        RECT 143.360 42.080 143.990 42.390 ;
        RECT 148.840 42.380 153.840 44.340 ;
        RECT 189.930 43.710 190.540 44.170 ;
        RECT 149.550 42.080 150.350 42.085 ;
        RECT 136.235 42.075 137.035 42.080 ;
        RECT 123.985 41.580 137.035 42.075 ;
        RECT 123.985 40.435 124.785 41.580 ;
        RECT 136.235 40.435 137.035 41.580 ;
        RECT 123.985 39.480 137.035 40.435 ;
        RECT 123.985 38.385 124.785 39.480 ;
        RECT 136.235 38.385 137.035 39.480 ;
        RECT 123.985 37.430 137.035 38.385 ;
        RECT 123.985 36.235 124.785 37.430 ;
        RECT 136.235 36.235 137.035 37.430 ;
        RECT 123.985 35.280 137.035 36.235 ;
        RECT 123.985 34.185 124.785 35.280 ;
        RECT 136.235 34.185 137.035 35.280 ;
        RECT 123.985 33.230 137.035 34.185 ;
        RECT 123.985 32.085 124.785 33.230 ;
        RECT 136.235 32.085 137.035 33.230 ;
        RECT 123.985 31.130 137.035 32.085 ;
        RECT 123.985 30.035 124.785 31.130 ;
        RECT 136.235 30.035 137.035 31.130 ;
        RECT 123.985 29.080 137.035 30.035 ;
        RECT 123.985 27.930 124.785 29.080 ;
        RECT 136.235 27.930 137.035 29.080 ;
        RECT 123.985 27.280 137.035 27.930 ;
        RECT 137.300 41.585 150.350 42.080 ;
        RECT 137.300 40.440 138.100 41.585 ;
        RECT 149.550 40.440 150.350 41.585 ;
        RECT 137.300 39.485 150.350 40.440 ;
        RECT 137.300 38.390 138.100 39.485 ;
        RECT 149.550 38.390 150.350 39.485 ;
        RECT 137.300 37.435 150.350 38.390 ;
        RECT 137.300 36.240 138.100 37.435 ;
        RECT 149.550 36.240 150.350 37.435 ;
        RECT 250.470 36.740 252.980 38.960 ;
        RECT 271.850 38.440 274.360 40.660 ;
        RECT 272.160 36.810 274.320 37.170 ;
        RECT 137.300 35.285 150.350 36.240 ;
        RECT 137.300 34.190 138.100 35.285 ;
        RECT 149.550 34.190 150.350 35.285 ;
        RECT 272.230 35.210 274.430 35.600 ;
        RECT 137.300 33.235 150.350 34.190 ;
        RECT 137.300 32.090 138.100 33.235 ;
        RECT 149.550 32.090 150.350 33.235 ;
        RECT 137.300 31.135 150.350 32.090 ;
        RECT 137.300 30.040 138.100 31.135 ;
        RECT 149.550 30.040 150.350 31.135 ;
        RECT 137.300 29.085 150.350 30.040 ;
        RECT 137.300 27.935 138.100 29.085 ;
        RECT 149.550 27.935 150.350 29.085 ;
        RECT 137.300 27.320 150.350 27.935 ;
        RECT 137.300 27.285 144.010 27.320 ;
        RECT 144.160 27.285 150.350 27.320 ;
        RECT 116.230 25.720 116.890 27.280 ;
        RECT 127.250 27.270 128.090 27.280 ;
        RECT 116.260 25.670 116.890 25.720 ;
        RECT 116.010 24.660 117.180 25.070 ;
        RECT 118.210 24.940 119.020 25.650 ;
        RECT 129.370 25.490 130.000 27.280 ;
        RECT 140.650 27.270 141.490 27.285 ;
        RECT 143.340 25.660 144.010 27.285 ;
        RECT 143.410 25.650 143.950 25.660 ;
        RECT 119.480 24.890 119.920 25.460 ;
        RECT 131.280 24.790 132.090 25.500 ;
        RECT 129.410 24.550 129.950 24.780 ;
        RECT 143.410 24.680 143.950 24.910 ;
        RECT 145.200 24.870 146.010 25.580 ;
        RECT 106.280 22.050 108.800 22.660 ;
        RECT 116.010 22.050 117.180 22.060 ;
        RECT 151.960 22.050 153.840 32.700 ;
        RECT 303.060 29.330 304.080 53.380 ;
        RECT 377.870 53.170 378.170 57.240 ;
        RECT 377.850 52.150 378.170 53.170 ;
        RECT 377.850 44.680 378.150 52.150 ;
        RECT 377.830 43.750 378.150 44.680 ;
        RECT 377.830 37.420 378.130 43.750 ;
        RECT 377.800 35.260 378.130 37.420 ;
        RECT 377.800 32.480 378.100 35.260 ;
        RECT 378.710 34.430 379.180 57.370 ;
        RECT 453.850 55.930 508.340 60.530 ;
        RECT 378.640 33.490 379.180 34.430 ;
        RECT 294.710 29.230 304.080 29.330 ;
        RECT 293.060 29.195 304.080 29.230 ;
        RECT 293.050 29.000 304.080 29.195 ;
        RECT 293.050 28.965 295.330 29.000 ;
        RECT 293.060 28.950 295.330 28.965 ;
        RECT 270.660 25.930 274.690 25.970 ;
        RECT 270.660 25.920 275.840 25.930 ;
        RECT 270.660 25.880 279.850 25.920 ;
        RECT 270.660 25.660 279.860 25.880 ;
        RECT 270.690 25.650 279.860 25.660 ;
        RECT 249.830 25.280 270.080 25.290 ;
        RECT 249.830 25.020 270.090 25.280 ;
        RECT 257.650 23.170 257.790 25.020 ;
        RECT 269.830 23.840 270.090 25.020 ;
        RECT 249.550 22.910 257.510 23.170 ;
        RECT 249.660 22.900 257.510 22.910 ;
        RECT 257.650 22.940 257.800 23.170 ;
        RECT 249.660 22.880 257.430 22.900 ;
        RECT 249.710 22.830 257.430 22.880 ;
        RECT 257.650 22.770 257.820 22.940 ;
        RECT 257.590 22.760 257.820 22.770 ;
        RECT 257.560 22.730 257.820 22.760 ;
        RECT 106.280 21.540 153.840 22.050 ;
        RECT 106.280 20.520 153.830 21.540 ;
        RECT 257.540 21.480 257.820 22.730 ;
        RECT 274.660 21.630 274.970 25.500 ;
        RECT 279.620 25.490 279.860 25.650 ;
        RECT 279.610 23.790 279.890 25.490 ;
        RECT 280.950 23.920 281.290 28.930 ;
        RECT 282.240 26.480 282.590 28.940 ;
        RECT 288.550 26.630 288.860 28.360 ;
        RECT 286.320 26.500 286.560 26.510 ;
        RECT 284.690 26.490 288.410 26.500 ;
        RECT 284.550 26.480 288.410 26.490 ;
        RECT 282.240 26.020 283.640 26.480 ;
        RECT 284.550 26.150 288.540 26.480 ;
        RECT 282.240 23.920 282.590 26.020 ;
        RECT 282.290 23.750 282.540 23.920 ;
        RECT 281.290 23.490 282.540 23.750 ;
        RECT 282.980 21.770 283.240 23.060 ;
        RECT 283.020 21.630 283.190 21.770 ;
        RECT 257.590 21.160 257.820 21.480 ;
        RECT 258.400 21.380 283.190 21.630 ;
        RECT 258.400 21.370 282.960 21.380 ;
        RECT 258.400 21.360 266.830 21.370 ;
        RECT 267.200 21.360 282.960 21.370 ;
        RECT 106.280 19.990 108.800 20.520 ;
        RECT 116.010 20.400 117.180 20.520 ;
        RECT 257.590 20.150 257.790 21.160 ;
        RECT 268.320 20.850 268.870 20.860 ;
        RECT 270.380 20.850 270.840 21.360 ;
        RECT 274.660 21.340 274.970 21.360 ;
        RECT 258.510 20.570 283.030 20.850 ;
        RECT 258.510 20.560 282.910 20.570 ;
        RECT 249.600 20.130 257.790 20.150 ;
        RECT 106.500 13.860 108.600 19.990 ;
        RECT 249.600 19.900 257.800 20.130 ;
        RECT 121.260 15.900 124.300 15.960 ;
        RECT 121.240 15.500 124.300 15.900 ;
        RECT 105.760 11.700 109.280 13.860 ;
        RECT 113.440 12.710 119.380 15.030 ;
        RECT 121.240 14.090 121.670 15.500 ;
        RECT 115.800 12.700 117.510 12.710 ;
        RECT 115.980 11.700 116.890 12.700 ;
        RECT 105.760 11.120 116.890 11.700 ;
        RECT 121.260 11.550 121.660 14.090 ;
        RECT 128.090 11.610 129.490 19.850 ;
        RECT 145.840 19.800 146.340 19.890 ;
        RECT 249.600 19.870 257.530 19.900 ;
        RECT 249.700 19.850 257.530 19.870 ;
        RECT 249.700 19.800 257.430 19.850 ;
        RECT 145.840 18.270 147.160 19.800 ;
        RECT 249.300 18.450 249.570 19.730 ;
        RECT 257.580 18.440 257.880 19.700 ;
        RECT 138.170 15.810 141.210 15.870 ;
        RECT 138.150 15.410 141.210 15.810 ;
        RECT 130.350 12.620 136.290 14.940 ;
        RECT 138.150 14.460 138.580 15.410 ;
        RECT 140.940 14.940 142.700 14.970 ;
        RECT 138.150 14.000 138.760 14.460 ;
        RECT 140.930 14.080 142.700 14.940 ;
        RECT 140.930 14.040 141.160 14.080 ;
        RECT 138.170 13.850 138.760 14.000 ;
        RECT 132.710 12.610 134.420 12.620 ;
        RECT 132.890 11.610 133.800 12.610 ;
        RECT 105.760 11.080 116.870 11.120 ;
        RECT 121.240 11.090 124.250 11.550 ;
        RECT 105.760 9.430 109.280 11.080 ;
        RECT 121.240 9.580 121.700 11.090 ;
        RECT 128.090 11.030 133.800 11.610 ;
        RECT 138.170 11.460 138.570 13.850 ;
        RECT 142.450 12.590 142.700 14.080 ;
        RECT 143.300 12.590 144.290 12.610 ;
        RECT 142.440 12.120 144.290 12.590 ;
        RECT 128.090 10.990 133.780 11.030 ;
        RECT 138.150 11.000 141.160 11.460 ;
        RECT 128.090 10.960 129.490 10.990 ;
        RECT 123.690 10.380 123.970 10.440 ;
        RECT 123.690 10.150 123.980 10.380 ;
        RECT 123.690 10.120 123.970 10.150 ;
        RECT 117.010 9.550 121.700 9.580 ;
        RECT 115.880 7.180 121.700 9.550 ;
        RECT 138.150 9.490 138.610 11.000 ;
        RECT 142.450 10.840 142.700 12.120 ;
        RECT 140.840 10.820 142.700 10.840 ;
        RECT 140.830 10.530 142.700 10.820 ;
        RECT 140.830 10.500 141.110 10.530 ;
        RECT 142.450 10.500 142.700 10.530 ;
        RECT 140.600 10.290 140.880 10.350 ;
        RECT 140.600 10.060 140.890 10.290 ;
        RECT 140.600 10.030 140.880 10.060 ;
        RECT 133.920 9.460 138.610 9.490 ;
        RECT 115.880 5.450 121.680 7.180 ;
        RECT 115.890 5.410 116.690 5.450 ;
        RECT 117.010 5.440 121.680 5.450 ;
        RECT 132.790 7.090 138.610 9.460 ;
        RECT 132.790 5.360 138.590 7.090 ;
        RECT 132.800 5.320 133.600 5.360 ;
        RECT 133.920 5.350 138.590 5.360 ;
        RECT 116.120 3.460 116.730 3.920 ;
        RECT 133.030 3.370 133.640 3.830 ;
        RECT 143.300 0.000 144.290 12.120 ;
        RECT 145.950 11.700 147.160 18.270 ;
        RECT 156.640 15.900 159.680 15.960 ;
        RECT 156.620 15.500 159.680 15.900 ;
        RECT 148.820 12.710 154.760 15.030 ;
        RECT 156.620 14.590 157.050 15.500 ;
        RECT 159.410 15.030 161.170 15.060 ;
        RECT 156.580 13.960 157.200 14.590 ;
        RECT 159.400 14.170 161.170 15.030 ;
        RECT 268.320 14.570 268.870 20.560 ;
        RECT 283.040 15.600 283.330 20.430 ;
        RECT 283.470 15.020 283.640 26.020 ;
        RECT 284.260 25.590 285.220 25.600 ;
        RECT 286.250 25.590 286.560 26.150 ;
        RECT 284.100 25.540 292.080 25.590 ;
        RECT 284.100 25.270 292.090 25.540 ;
        RECT 292.100 25.120 292.350 25.130 ;
        RECT 288.590 24.430 288.940 24.460 ;
        RECT 292.070 24.440 292.390 25.120 ;
        RECT 292.070 24.430 292.350 24.440 ;
        RECT 288.590 24.050 292.350 24.430 ;
        RECT 284.280 22.380 288.300 22.680 ;
        RECT 287.630 22.100 288.060 22.380 ;
        RECT 288.590 22.230 288.940 24.050 ;
        RECT 292.740 23.750 293.030 28.770 ;
        RECT 295.060 28.760 295.330 28.950 ;
        RECT 303.060 28.780 304.080 29.000 ;
        RECT 295.010 24.170 295.350 28.760 ;
        RECT 295.010 24.090 295.470 24.170 ;
        RECT 295.010 23.770 295.490 24.090 ;
        RECT 295.010 23.740 295.470 23.770 ;
        RECT 294.050 23.190 295.010 23.210 ;
        RECT 289.530 22.980 290.530 23.000 ;
        RECT 289.520 22.960 290.530 22.980 ;
        RECT 293.400 22.990 295.030 23.190 ;
        RECT 293.400 22.960 293.590 22.990 ;
        RECT 294.050 22.980 295.010 22.990 ;
        RECT 289.520 22.940 291.820 22.960 ;
        RECT 293.400 22.940 293.560 22.960 ;
        RECT 289.520 22.730 293.560 22.940 ;
        RECT 295.190 22.820 295.470 23.740 ;
        RECT 295.060 22.790 295.470 22.820 ;
        RECT 289.530 22.720 293.560 22.730 ;
        RECT 289.530 22.700 291.820 22.720 ;
        RECT 288.310 22.100 288.940 22.230 ;
        RECT 287.630 21.760 288.940 22.100 ;
        RECT 288.050 21.750 288.940 21.760 ;
        RECT 290.520 22.690 291.690 22.700 ;
        RECT 288.310 21.190 288.590 21.750 ;
        RECT 290.520 19.570 290.820 22.690 ;
        RECT 295.040 22.540 295.470 22.790 ;
        RECT 295.060 22.470 295.470 22.540 ;
        RECT 295.060 21.800 295.290 22.470 ;
        RECT 294.050 21.410 295.010 21.640 ;
        RECT 377.760 19.960 378.120 32.480 ;
        RECT 378.640 22.930 379.110 33.490 ;
        RECT 510.620 24.950 514.060 77.140 ;
        RECT 521.130 53.450 524.990 109.260 ;
        RECT 538.080 108.650 541.720 110.190 ;
        RECT 538.360 82.690 541.720 108.650 ;
        RECT 536.610 77.580 543.320 82.690 ;
        RECT 565.030 78.530 572.050 109.980 ;
        RECT 565.030 76.780 572.530 78.530 ;
        RECT 565.560 56.810 572.530 76.780 ;
        RECT 522.460 43.240 524.990 53.450 ;
        RECT 547.840 43.240 549.820 44.050 ;
        RECT 522.460 43.030 549.820 43.240 ;
        RECT 522.460 24.950 524.990 43.030 ;
        RECT 547.840 41.870 549.820 43.030 ;
        RECT 530.970 29.490 533.090 31.610 ;
        RECT 378.600 22.910 393.060 22.930 ;
        RECT 495.690 22.910 510.150 22.930 ;
        RECT 523.600 22.910 523.820 24.950 ;
        RECT 378.600 22.890 416.260 22.910 ;
        RECT 481.730 22.890 523.830 22.910 ;
        RECT 378.600 22.870 428.940 22.890 ;
        RECT 454.140 22.870 523.830 22.890 ;
        RECT 378.600 22.660 523.830 22.870 ;
        RECT 378.640 22.650 379.110 22.660 ;
        RECT 388.980 22.640 496.190 22.660 ;
        RECT 509.370 22.640 523.830 22.660 ;
        RECT 394.920 22.630 398.290 22.640 ;
        RECT 414.480 22.620 482.050 22.640 ;
        RECT 426.510 22.600 454.710 22.620 ;
        RECT 531.620 19.960 532.430 29.490 ;
        RECT 377.760 19.000 532.430 19.960 ;
        RECT 377.760 18.960 532.350 19.000 ;
        RECT 377.760 18.950 395.110 18.960 ;
        RECT 397.810 18.950 532.350 18.960 ;
        RECT 307.910 15.250 312.120 16.500 ;
        RECT 297.990 15.050 301.960 15.070 ;
        RECT 303.990 15.050 312.120 15.250 ;
        RECT 297.990 15.020 312.120 15.050 ;
        RECT 258.460 14.300 283.030 14.570 ;
        RECT 283.460 14.430 312.120 15.020 ;
        RECT 258.460 14.290 282.910 14.300 ;
        RECT 283.470 14.170 283.640 14.430 ;
        RECT 297.990 14.400 312.120 14.430 ;
        RECT 300.890 14.380 312.120 14.400 ;
        RECT 303.990 14.360 312.120 14.380 ;
        RECT 159.400 14.130 159.630 14.170 ;
        RECT 151.180 12.700 152.890 12.710 ;
        RECT 151.360 11.700 152.270 12.700 ;
        RECT 145.950 11.120 152.270 11.700 ;
        RECT 156.640 11.550 157.040 13.960 ;
        RECT 160.920 12.680 161.170 14.170 ;
        RECT 283.260 14.160 283.640 14.170 ;
        RECT 283.050 14.100 283.640 14.160 ;
        RECT 283.020 13.930 283.640 14.100 ;
        RECT 283.020 13.770 283.630 13.930 ;
        RECT 161.690 12.680 162.680 12.780 ;
        RECT 160.910 12.210 162.680 12.680 ;
        RECT 283.050 12.670 283.350 13.770 ;
        RECT 307.910 13.350 312.120 14.360 ;
        RECT 283.060 12.650 283.320 12.670 ;
        RECT 145.950 11.080 152.250 11.120 ;
        RECT 156.620 11.090 159.630 11.550 ;
        RECT 145.950 11.020 147.160 11.080 ;
        RECT 156.620 9.580 157.080 11.090 ;
        RECT 160.920 10.930 161.170 12.210 ;
        RECT 159.310 10.910 161.170 10.930 ;
        RECT 159.300 10.620 161.170 10.910 ;
        RECT 159.300 10.590 159.580 10.620 ;
        RECT 160.920 10.590 161.170 10.620 ;
        RECT 159.070 10.380 159.350 10.440 ;
        RECT 159.070 10.150 159.360 10.380 ;
        RECT 159.070 10.120 159.350 10.150 ;
        RECT 152.390 9.550 157.080 9.580 ;
        RECT 151.260 7.180 157.080 9.550 ;
        RECT 151.260 5.450 157.060 7.180 ;
        RECT 151.270 5.410 152.070 5.450 ;
        RECT 152.390 5.440 157.060 5.450 ;
        RECT 161.690 4.830 162.680 12.210 ;
        RECT 151.500 3.460 152.110 3.920 ;
        RECT 161.690 3.800 162.700 4.830 ;
        RECT 161.750 1.660 162.700 3.800 ;
        RECT 161.690 0.200 162.700 1.660 ;
        RECT 161.690 0.170 162.680 0.200 ;
      LAYER via ;
        RECT 448.360 205.400 449.360 206.950 ;
        RECT 475.580 195.160 477.420 196.550 ;
        RECT 169.010 159.160 169.270 159.420 ;
        RECT 171.100 159.140 171.360 159.400 ;
        RECT 168.930 157.660 169.190 157.920 ;
        RECT 168.730 156.250 169.010 156.730 ;
        RECT 170.820 156.300 171.080 156.730 ;
        RECT 174.440 160.440 174.810 160.800 ;
        RECT 173.090 155.590 173.460 155.920 ;
        RECT 354.940 155.100 355.360 155.540 ;
        RECT 373.240 152.030 373.970 152.650 ;
        RECT 378.490 152.100 378.940 152.520 ;
        RECT 134.970 133.570 135.900 134.530 ;
        RECT 114.940 109.070 115.290 109.330 ;
        RECT 118.390 108.660 118.730 109.320 ;
        RECT 122.970 108.650 123.310 109.310 ;
        RECT 155.730 133.310 156.470 133.800 ;
        RECT 177.050 133.080 177.650 133.580 ;
        RECT 475.230 148.110 476.050 150.870 ;
        RECT 530.520 150.500 531.070 152.430 ;
        RECT 588.580 204.410 590.500 206.180 ;
        RECT 558.090 148.240 558.490 150.490 ;
        RECT 311.590 131.750 311.850 132.010 ;
        RECT 318.370 131.890 318.655 132.150 ;
        RECT 325.250 131.770 325.530 132.030 ;
        RECT 341.430 132.270 342.140 132.910 ;
        RECT 332.060 131.020 332.390 131.370 ;
        RECT 337.440 131.360 338.320 132.030 ;
        RECT 343.910 127.230 345.170 128.260 ;
        RECT 321.550 125.710 321.870 126.110 ;
        RECT 323.390 125.650 323.650 125.920 ;
        RECT 330.150 125.790 330.410 126.060 ;
        RECT 339.520 125.380 340.160 126.230 ;
        RECT 330.050 122.420 330.630 122.930 ;
        RECT 122.920 100.510 123.230 100.850 ;
        RECT 234.280 107.470 236.440 107.820 ;
        RECT 255.690 107.470 257.850 107.820 ;
        RECT 281.670 107.480 283.810 107.830 ;
        RECT 234.280 105.880 236.440 106.230 ;
        RECT 255.690 105.880 257.850 106.230 ;
        RECT 281.680 105.880 283.820 106.230 ;
        RECT 255.690 104.290 257.850 104.640 ;
        RECT 260.250 104.300 262.420 104.670 ;
        RECT 281.680 104.300 283.820 104.650 ;
        RECT 106.560 93.650 107.790 94.740 ;
        RECT 135.540 100.440 135.950 100.810 ;
        RECT 145.700 100.580 146.140 100.890 ;
        RECT 152.970 100.660 153.780 101.540 ;
        RECT 255.690 102.700 257.850 103.060 ;
        RECT 255.690 101.110 257.850 101.470 ;
        RECT 234.280 99.520 236.440 99.870 ;
        RECT 260.260 102.710 262.420 103.060 ;
        RECT 281.670 102.710 283.830 103.060 ;
        RECT 260.260 101.120 262.420 101.470 ;
        RECT 281.670 101.120 283.830 101.470 ;
        RECT 255.690 99.510 257.850 99.880 ;
        RECT 281.670 99.530 283.830 99.880 ;
        RECT 234.280 97.930 236.410 98.290 ;
        RECT 152.970 96.030 153.780 96.910 ;
        RECT 260.250 97.930 262.440 98.300 ;
        RECT 234.280 96.340 236.410 96.700 ;
        RECT 260.250 96.360 262.430 96.710 ;
        RECT 117.170 83.230 117.490 83.610 ;
        RECT 131.860 83.350 132.120 83.610 ;
        RECT 144.420 83.260 144.700 83.610 ;
        RECT 24.900 74.300 25.570 74.990 ;
        RECT 20.220 71.400 20.930 72.030 ;
        RECT 18.830 70.390 19.580 71.060 ;
        RECT 22.510 69.060 23.030 69.660 ;
        RECT 24.790 66.450 25.310 67.050 ;
        RECT 27.100 64.060 27.430 64.430 ;
        RECT 255.700 94.750 257.840 95.110 ;
        RECT 260.250 94.760 262.430 95.110 ;
        RECT 227.100 89.750 227.700 90.140 ;
        RECT 244.060 88.900 244.750 89.530 ;
        RECT 245.590 88.650 245.850 89.150 ;
        RECT 246.490 88.710 246.750 89.130 ;
        RECT 250.110 88.750 250.500 89.240 ;
        RECT 259.000 88.720 259.440 89.380 ;
        RECT 247.030 87.450 247.910 87.710 ;
        RECT 271.330 87.650 271.740 88.080 ;
        RECT 278.530 87.720 278.830 87.990 ;
        RECT 281.410 88.000 281.720 88.300 ;
        RECT 244.720 86.800 245.260 87.230 ;
        RECT 261.920 85.430 262.200 85.690 ;
        RECT 275.540 85.200 275.800 85.540 ;
        RECT 212.380 81.200 212.680 81.520 ;
        RECT 214.370 81.110 214.690 81.430 ;
        RECT 214.900 81.640 215.290 81.990 ;
        RECT 215.520 80.610 215.880 80.940 ;
        RECT 216.620 81.680 216.980 82.010 ;
        RECT 212.780 78.450 213.070 78.740 ;
        RECT 216.660 78.440 216.950 78.730 ;
        RECT 238.310 81.290 238.610 81.610 ;
        RECT 240.300 81.200 240.620 81.520 ;
        RECT 240.830 81.730 241.220 82.080 ;
        RECT 241.450 80.700 241.810 81.030 ;
        RECT 242.550 81.770 242.910 82.100 ;
        RECT 264.190 81.350 264.490 81.670 ;
        RECT 238.710 78.540 239.000 78.830 ;
        RECT 242.590 78.530 242.880 78.820 ;
        RECT 247.190 79.160 247.720 79.430 ;
        RECT 266.180 81.260 266.500 81.580 ;
        RECT 266.710 81.790 267.100 82.140 ;
        RECT 267.330 80.760 267.690 81.090 ;
        RECT 268.430 81.830 268.790 82.160 ;
        RECT 264.590 78.600 264.880 78.890 ;
        RECT 152.970 76.620 153.780 77.500 ;
        RECT 134.440 75.840 134.970 76.220 ;
        RECT 145.600 75.760 146.200 76.460 ;
        RECT 218.490 76.180 218.870 76.520 ;
        RECT 260.010 77.830 261.020 78.440 ;
        RECT 268.470 78.590 268.760 78.880 ;
        RECT 260.260 76.580 260.860 76.860 ;
        RECT 44.530 71.730 44.900 72.180 ;
        RECT 47.210 71.340 47.620 71.750 ;
        RECT 43.690 69.990 44.320 70.000 ;
        RECT 43.690 69.730 44.360 69.990 ;
        RECT 43.690 69.720 44.320 69.730 ;
        RECT 119.740 74.760 120.090 75.110 ;
        RECT 106.700 71.630 107.510 72.510 ;
        RECT 152.970 71.990 153.780 72.870 ;
        RECT 47.110 68.260 47.520 68.670 ;
        RECT 84.260 68.680 84.640 68.960 ;
        RECT 43.770 66.670 44.400 66.940 ;
        RECT 47.140 65.370 47.550 65.780 ;
        RECT 47.170 62.490 47.580 62.900 ;
        RECT 25.940 61.510 26.460 62.110 ;
        RECT 21.090 59.960 21.400 60.320 ;
        RECT 43.800 60.910 44.420 61.190 ;
        RECT 47.150 59.620 47.560 60.030 ;
        RECT 21.160 59.020 21.420 59.350 ;
        RECT 21.200 58.090 21.460 58.370 ;
        RECT 39.820 57.630 40.760 58.580 ;
        RECT 106.700 67.000 107.510 67.880 ;
        RECT 25.770 56.160 26.290 56.760 ;
        RECT 47.160 56.710 47.570 57.120 ;
        RECT 39.460 54.680 40.080 55.510 ;
        RECT 84.440 54.420 85.310 55.190 ;
        RECT 27.080 53.850 27.450 54.230 ;
        RECT 47.260 53.800 47.670 54.210 ;
        RECT 25.000 51.270 25.520 51.850 ;
        RECT 39.540 51.760 40.190 52.750 ;
        RECT 47.240 50.920 47.650 51.330 ;
        RECT 84.390 50.780 85.000 51.370 ;
        RECT 26.150 48.690 26.670 49.270 ;
        RECT 24.930 46.010 25.490 46.630 ;
        RECT 43.440 48.420 43.750 48.740 ;
        RECT 43.770 46.480 44.400 46.760 ;
        RECT 236.990 71.450 237.660 71.780 ;
        RECT 261.130 75.700 261.750 75.960 ;
        RECT 261.080 69.800 261.670 70.110 ;
        RECT 295.240 82.970 295.710 83.340 ;
        RECT 290.760 82.160 291.170 82.660 ;
        RECT 292.470 80.310 292.770 80.630 ;
        RECT 294.460 80.220 294.780 80.540 ;
        RECT 294.990 80.750 295.380 81.100 ;
        RECT 295.610 79.720 295.970 80.050 ;
        RECT 296.710 80.790 297.070 81.120 ;
        RECT 292.870 77.560 293.160 77.850 ;
        RECT 296.750 77.550 297.040 77.840 ;
        RECT 304.770 76.450 305.230 76.730 ;
        RECT 271.820 74.190 272.760 74.650 ;
        RECT 268.980 67.600 269.700 68.260 ;
        RECT 117.070 54.550 117.380 55.080 ;
        RECT 396.260 120.040 397.200 120.920 ;
        RECT 407.750 121.180 408.750 122.350 ;
        RECT 456.470 108.840 457.010 109.160 ;
        RECT 380.660 91.950 381.590 92.690 ;
        RECT 380.250 73.430 380.870 74.310 ;
        RECT 483.700 109.330 484.240 109.650 ;
        RECT 512.980 108.720 515.070 109.610 ;
        RECT 522.500 109.900 523.820 110.380 ;
        RECT 482.150 77.180 486.990 81.210 ;
        RECT 131.380 54.280 131.690 54.810 ;
        RECT 143.510 54.360 143.820 54.890 ;
        RECT 179.800 54.220 181.190 55.060 ;
        RECT 294.820 54.110 295.940 55.980 ;
        RECT 203.510 52.510 203.970 52.830 ;
        RECT 106.700 46.720 107.510 47.600 ;
        RECT 119.090 46.050 119.580 46.820 ;
        RECT 132.890 46.490 133.190 47.010 ;
        RECT 145.420 46.180 145.980 46.860 ;
        RECT 85.230 42.890 85.750 43.240 ;
        RECT 106.700 42.480 107.510 43.360 ;
        RECT 152.170 42.610 153.430 44.090 ;
        RECT 272.230 36.840 274.240 37.130 ;
        RECT 272.330 35.250 274.340 35.540 ;
        RECT 152.360 31.470 153.480 32.640 ;
        RECT 118.350 25.070 118.900 25.530 ;
        RECT 131.380 24.860 131.930 25.320 ;
        RECT 145.280 24.990 145.830 25.450 ;
        RECT 455.580 57.880 456.910 58.810 ;
        RECT 538.660 109.070 540.750 109.960 ;
        RECT 567.340 108.590 569.630 109.230 ;
        RECT 511.730 43.190 513.050 44.530 ;
        RECT 270.730 25.680 274.630 25.940 ;
        RECT 249.610 22.910 257.450 23.170 ;
        RECT 106.780 20.740 108.250 22.050 ;
        RECT 279.620 23.830 279.880 25.460 ;
        RECT 280.990 23.990 281.270 28.870 ;
        RECT 288.560 26.690 288.830 28.310 ;
        RECT 258.450 21.360 266.320 21.620 ;
        RECT 128.340 18.620 129.420 19.750 ;
        RECT 145.880 18.570 147.130 19.470 ;
        RECT 249.300 18.480 249.560 19.690 ;
        RECT 257.600 18.510 257.860 19.670 ;
        RECT 283.050 15.660 283.320 20.380 ;
        RECT 284.150 25.290 292.000 25.580 ;
        RECT 292.100 24.640 292.360 25.070 ;
        RECT 292.750 23.820 293.010 28.710 ;
        RECT 289.610 22.700 290.450 22.980 ;
        RECT 548.260 42.320 549.410 43.530 ;
        RECT 531.330 29.900 532.760 31.250 ;
        RECT 309.610 13.960 310.860 15.590 ;
        RECT 143.460 3.440 144.060 4.160 ;
        RECT 162.050 2.200 162.500 2.720 ;
      LAYER met2 ;
        RECT 447.640 208.670 448.320 208.720 ;
        RECT 447.640 208.630 448.380 208.670 ;
        RECT 447.560 204.110 450.970 208.630 ;
        RECT 174.360 160.360 174.890 160.870 ;
        RECT 168.870 158.260 171.470 160.270 ;
        RECT 168.100 157.970 169.230 157.980 ;
        RECT 167.660 157.610 169.230 157.970 ;
        RECT 167.660 157.440 168.150 157.610 ;
        RECT 168.920 157.600 169.230 157.610 ;
        RECT 168.660 156.680 171.160 157.030 ;
        RECT 166.750 156.390 171.160 156.680 ;
        RECT 166.750 154.680 167.040 156.390 ;
        RECT 168.660 156.040 171.160 156.390 ;
        RECT 354.570 156.030 355.580 156.070 ;
        RECT 173.020 155.500 173.540 156.010 ;
        RECT 166.690 154.270 167.040 154.680 ;
        RECT 354.090 154.470 355.580 156.030 ;
        RECT 354.090 154.400 354.540 154.470 ;
        RECT 166.690 141.030 167.030 154.270 ;
        RECT 106.710 140.690 167.080 141.030 ;
        RECT 106.710 140.670 115.570 140.690 ;
        RECT 23.890 77.960 40.600 78.000 ;
        RECT 23.890 76.850 40.700 77.960 ;
        RECT 18.950 71.230 19.630 71.400 ;
        RECT 18.700 70.270 19.720 71.230 ;
        RECT 20.040 71.220 21.140 72.170 ;
        RECT 18.950 59.440 19.630 70.270 ;
        RECT 20.270 64.540 20.970 71.220 ;
        RECT 22.450 69.850 23.060 72.020 ;
        RECT 23.890 71.790 24.470 76.850 ;
        RECT 24.760 74.990 25.690 75.130 ;
        RECT 34.690 74.990 35.920 75.040 ;
        RECT 24.760 74.220 35.920 74.990 ;
        RECT 24.760 74.160 25.690 74.220 ;
        RECT 23.980 71.260 24.430 71.790 ;
        RECT 22.370 68.920 23.380 69.850 ;
        RECT 23.990 67.140 24.410 71.260 ;
        RECT 24.670 67.140 25.410 67.150 ;
        RECT 23.990 66.530 25.410 67.140 ;
        RECT 24.670 66.350 25.410 66.530 ;
        RECT 25.550 64.540 25.780 64.550 ;
        RECT 20.270 64.530 21.010 64.540 ;
        RECT 25.550 64.530 27.100 64.540 ;
        RECT 20.270 64.500 27.100 64.530 ;
        RECT 20.270 64.490 27.460 64.500 ;
        RECT 20.270 64.050 27.520 64.490 ;
        RECT 20.270 64.000 20.970 64.050 ;
        RECT 25.560 64.020 27.520 64.050 ;
        RECT 20.280 60.360 20.820 64.000 ;
        RECT 25.700 63.990 27.520 64.020 ;
        RECT 26.010 62.220 26.620 62.250 ;
        RECT 25.820 61.380 26.620 62.220 ;
        RECT 20.280 59.920 21.420 60.360 ;
        RECT 20.330 59.890 21.420 59.920 ;
        RECT 18.920 59.400 21.420 59.440 ;
        RECT 18.920 58.960 21.470 59.400 ;
        RECT 18.920 58.890 21.420 58.960 ;
        RECT 18.950 58.830 19.630 58.890 ;
        RECT 34.690 58.600 35.920 74.220 ;
        RECT 39.730 67.320 40.700 76.850 ;
        RECT 44.460 71.650 44.980 72.240 ;
        RECT 47.110 71.270 47.720 71.830 ;
        RECT 47.130 71.260 47.720 71.270 ;
        RECT 44.160 70.020 44.420 70.030 ;
        RECT 43.550 69.710 44.420 70.020 ;
        RECT 47.010 68.200 47.620 68.760 ;
        RECT 39.620 66.310 40.810 67.320 ;
        RECT 43.350 66.610 44.480 66.970 ;
        RECT 63.720 66.560 66.700 127.560 ;
        RECT 106.720 109.495 107.010 140.670 ;
        RECT 166.690 140.640 167.030 140.690 ;
        RECT 134.800 133.300 136.210 134.840 ;
        RECT 155.540 133.050 156.920 134.240 ;
        RECT 176.870 132.830 178.080 133.840 ;
        RECT 337.290 132.180 338.490 132.220 ;
        RECT 318.310 132.030 318.700 132.180 ;
        RECT 311.510 131.700 318.700 132.030 ;
        RECT 311.510 131.690 311.880 131.700 ;
        RECT 318.030 131.690 318.700 131.700 ;
        RECT 325.080 132.040 325.790 132.140 ;
        RECT 325.080 131.690 332.500 132.040 ;
        RECT 318.030 131.490 318.310 131.690 ;
        RECT 325.080 131.510 325.790 131.690 ;
        RECT 318.030 126.070 318.300 131.490 ;
        RECT 332.090 131.400 332.490 131.690 ;
        RECT 332.060 131.390 332.490 131.400 ;
        RECT 331.770 131.360 332.490 131.390 ;
        RECT 331.770 131.060 332.530 131.360 ;
        RECT 337.270 131.240 338.580 132.180 ;
        RECT 340.880 131.750 342.750 133.420 ;
        RECT 337.290 131.220 338.490 131.240 ;
        RECT 331.770 130.890 332.490 131.060 ;
        RECT 332.040 130.860 332.490 130.890 ;
        RECT 332.040 129.780 332.410 130.860 ;
        RECT 332.050 129.570 332.410 129.780 ;
        RECT 331.890 129.410 332.970 129.570 ;
        RECT 331.540 128.410 333.260 129.410 ;
        RECT 342.690 127.570 346.530 129.000 ;
        RECT 346.760 127.570 351.850 127.580 ;
        RECT 342.690 127.560 351.850 127.570 ;
        RECT 354.100 127.560 354.410 154.400 ;
        RECT 373.110 152.690 374.230 152.800 ;
        RECT 373.110 152.010 379.280 152.690 ;
        RECT 373.110 151.970 374.230 152.010 ;
        RECT 447.640 146.720 448.380 204.110 ;
        RECT 464.080 204.050 581.480 208.310 ;
        RECT 588.390 204.070 591.020 206.560 ;
        RECT 464.080 203.810 581.940 204.050 ;
        RECT 464.080 201.440 470.930 203.810 ;
        RECT 464.340 164.120 470.850 201.440 ;
        RECT 474.570 197.240 477.910 202.240 ;
        RECT 575.510 200.820 581.940 203.810 ;
        RECT 474.120 194.090 478.350 197.240 ;
        RECT 464.340 156.840 470.860 164.120 ;
        RECT 464.340 153.080 465.570 156.840 ;
        RECT 468.980 153.080 470.860 156.840 ;
        RECT 475.260 153.820 476.490 194.090 ;
        RECT 494.860 193.950 556.120 199.240 ;
        RECT 494.890 163.650 500.850 193.950 ;
        RECT 494.520 155.200 500.900 163.650 ;
        RECT 494.520 154.130 497.030 155.200 ;
        RECT 498.320 154.130 500.900 155.200 ;
        RECT 464.340 152.030 470.860 153.080 ;
        RECT 464.340 151.140 470.850 152.030 ;
        RECT 475.010 151.260 476.520 153.820 ;
        RECT 494.520 151.560 500.900 154.130 ;
        RECT 548.950 159.490 554.910 193.950 ;
        RECT 475.010 147.920 476.240 151.260 ;
        RECT 494.890 150.470 500.850 151.560 ;
        RECT 530.340 150.300 531.180 152.900 ;
        RECT 548.950 152.170 549.940 159.490 ;
        RECT 554.750 152.170 554.910 159.490 ;
        RECT 548.950 150.240 554.910 152.170 ;
        RECT 575.430 160.750 581.940 200.820 ;
        RECT 575.430 153.430 576.350 160.750 ;
        RECT 581.160 153.430 581.940 160.750 ;
        RECT 575.430 151.480 581.940 153.430 ;
        RECT 557.920 147.990 558.760 150.770 ;
        RECT 447.700 146.670 448.380 146.720 ;
        RECT 342.690 127.310 354.410 127.560 ;
        RECT 342.690 127.300 346.890 127.310 ;
        RECT 339.100 126.410 340.410 126.870 ;
        RECT 342.690 126.480 346.530 127.300 ;
        RECT 351.730 127.290 354.410 127.310 ;
        RECT 354.100 127.280 354.410 127.290 ;
        RECT 464.420 133.430 471.520 134.780 ;
        RECT 321.450 126.160 321.910 126.330 ;
        RECT 321.450 126.070 321.930 126.160 ;
        RECT 330.130 126.110 330.530 126.210 ;
        RECT 318.030 125.850 321.930 126.070 ;
        RECT 330.060 126.010 330.530 126.110 ;
        RECT 321.450 125.680 321.930 125.850 ;
        RECT 321.450 125.540 321.910 125.680 ;
        RECT 323.290 125.600 330.530 126.010 ;
        RECT 330.130 125.530 330.530 125.600 ;
        RECT 330.130 123.700 330.410 125.530 ;
        RECT 339.100 125.470 340.590 126.410 ;
        RECT 464.420 126.110 465.370 133.430 ;
        RECT 470.180 126.110 471.520 133.430 ;
        RECT 534.420 133.410 548.000 134.290 ;
        RECT 493.020 131.600 496.260 132.720 ;
        RECT 339.100 124.900 340.410 125.470 ;
        RECT 330.130 123.220 330.560 123.700 ;
        RECT 329.780 122.260 331.050 123.220 ;
        RECT 396.020 119.600 397.410 121.430 ;
        RECT 407.570 120.800 408.970 122.790 ;
        RECT 106.720 109.480 112.970 109.495 ;
        RECT 115.020 109.480 115.310 109.495 ;
        RECT 106.720 108.370 115.310 109.480 ;
        RECT 118.110 108.590 123.410 109.420 ;
        RECT 456.290 108.730 457.430 109.360 ;
        RECT 256.750 108.230 275.990 108.420 ;
        RECT 256.750 107.910 257.000 108.230 ;
        RECT 234.210 105.830 236.460 107.890 ;
        RECT 255.660 107.380 257.930 107.910 ;
        RECT 255.650 104.220 257.930 106.300 ;
        RECT 260.200 104.250 262.470 104.720 ;
        RECT 261.130 103.780 261.360 104.250 ;
        RECT 261.130 103.590 271.540 103.780 ;
        RECT 106.280 89.870 108.240 95.020 ;
        RECT 122.780 84.160 123.450 100.990 ;
        RECT 135.270 84.490 136.370 100.930 ;
        RECT 122.780 83.880 123.410 84.160 ;
        RECT 135.250 84.050 136.420 84.490 ;
        RECT 117.110 83.180 123.410 83.880 ;
        RECT 131.770 83.250 136.440 84.050 ;
        RECT 145.470 83.690 146.490 101.060 ;
        RECT 152.810 95.950 153.960 101.750 ;
        RECT 234.240 99.900 236.480 99.920 ;
        RECT 227.140 99.460 236.480 99.900 ;
        RECT 227.140 99.450 235.170 99.460 ;
        RECT 255.620 99.450 257.900 103.150 ;
        RECT 260.210 101.060 262.440 103.120 ;
        RECT 227.270 98.560 227.550 99.450 ;
        RECT 227.270 90.290 227.530 98.560 ;
        RECT 234.210 98.300 236.460 98.340 ;
        RECT 234.210 97.110 236.470 98.300 ;
        RECT 260.220 97.880 262.490 98.350 ;
        RECT 261.530 97.490 261.720 97.880 ;
        RECT 261.530 97.250 265.970 97.490 ;
        RECT 245.640 97.110 245.820 97.140 ;
        RECT 234.210 96.900 245.820 97.110 ;
        RECT 234.210 96.330 236.470 96.900 ;
        RECT 234.210 96.280 236.460 96.330 ;
        RECT 226.990 89.580 227.830 90.290 ;
        RECT 243.900 88.760 244.960 89.680 ;
        RECT 245.640 89.250 245.820 96.900 ;
        RECT 260.200 95.790 262.470 96.790 ;
        RECT 246.470 95.530 262.470 95.790 ;
        RECT 246.470 95.520 247.350 95.530 ;
        RECT 246.470 89.250 246.790 95.520 ;
        RECT 255.670 94.690 257.910 95.160 ;
        RECT 256.410 94.520 256.690 94.690 ;
        RECT 260.200 94.660 262.470 95.530 ;
        RECT 250.090 94.340 256.690 94.520 ;
        RECT 250.090 94.320 256.610 94.340 ;
        RECT 250.090 89.340 250.370 94.320 ;
        RECT 245.530 88.550 245.910 89.250 ;
        RECT 246.410 88.590 246.840 89.250 ;
        RECT 250.050 88.590 250.550 89.340 ;
        RECT 258.930 89.310 259.520 89.510 ;
        RECT 265.640 89.310 265.970 97.250 ;
        RECT 258.930 89.010 265.970 89.310 ;
        RECT 258.930 88.980 265.950 89.010 ;
        RECT 258.930 88.620 259.520 88.980 ;
        RECT 271.330 88.140 271.540 103.590 ;
        RECT 245.910 87.660 246.270 87.670 ;
        RECT 246.910 87.660 248.070 87.830 ;
        RECT 245.910 87.460 248.070 87.660 ;
        RECT 271.260 87.560 271.800 88.140 ;
        RECT 275.790 87.950 275.990 108.230 ;
        RECT 281.610 105.380 283.900 107.890 ;
        RECT 281.610 105.120 283.910 105.380 ;
        RECT 281.610 104.200 283.900 105.120 ;
        RECT 284.520 103.120 284.910 103.130 ;
        RECT 283.160 103.110 284.910 103.120 ;
        RECT 281.650 102.660 284.910 103.110 ;
        RECT 283.160 102.640 284.910 102.660 ;
        RECT 281.650 99.470 283.880 101.530 ;
        RECT 284.520 88.520 284.910 102.640 ;
        RECT 347.650 93.550 352.890 93.600 ;
        RECT 345.800 93.530 352.890 93.550 ;
        RECT 356.720 93.540 358.890 93.560 ;
        RECT 354.330 93.530 358.890 93.540 ;
        RECT 342.790 93.510 358.890 93.530 ;
        RECT 342.790 93.150 359.280 93.510 ;
        RECT 380.550 93.150 382.140 93.170 ;
        RECT 342.790 91.680 382.150 93.150 ;
        RECT 342.790 91.640 359.280 91.680 ;
        RECT 380.550 91.670 382.140 91.680 ;
        RECT 342.050 91.580 359.280 91.640 ;
        RECT 338.060 91.100 359.280 91.580 ;
        RECT 338.060 90.210 338.470 91.100 ;
        RECT 342.790 90.240 359.280 91.100 ;
        RECT 342.790 90.210 352.890 90.240 ;
        RECT 354.780 90.220 359.280 90.240 ;
        RECT 357.240 90.210 359.280 90.220 ;
        RECT 290.890 89.790 338.470 90.210 ;
        RECT 345.800 90.150 352.890 90.210 ;
        RECT 345.800 90.100 349.220 90.150 ;
        RECT 281.320 88.190 281.810 88.390 ;
        RECT 284.510 88.190 284.920 88.520 ;
        RECT 281.320 88.080 284.920 88.190 ;
        RECT 281.320 88.050 284.910 88.080 ;
        RECT 278.420 87.950 278.910 88.020 ;
        RECT 275.790 87.710 278.910 87.950 ;
        RECT 281.320 87.910 281.810 88.050 ;
        RECT 278.420 87.640 278.910 87.710 ;
        RECT 244.640 86.700 245.340 87.320 ;
        RECT 244.740 85.160 245.260 86.700 ;
        RECT 212.360 84.900 245.260 85.160 ;
        RECT 144.280 83.190 146.510 83.690 ;
        RECT 117.120 83.140 117.620 83.180 ;
        RECT 145.470 83.170 146.490 83.190 ;
        RECT 212.360 82.320 212.730 84.900 ;
        RECT 245.910 84.170 246.270 87.460 ;
        RECT 246.910 87.350 248.070 87.460 ;
        RECT 261.790 85.730 262.320 85.750 ;
        RECT 261.790 85.690 262.460 85.730 ;
        RECT 261.460 85.370 262.460 85.690 ;
        RECT 261.790 85.230 262.460 85.370 ;
        RECT 217.760 83.890 246.270 84.170 ;
        RECT 213.400 82.320 213.670 82.330 ;
        RECT 212.290 82.290 213.670 82.320 ;
        RECT 214.370 82.300 214.720 82.320 ;
        RECT 214.360 82.290 214.720 82.300 ;
        RECT 212.290 80.320 214.720 82.290 ;
        RECT 214.860 82.010 217.000 82.320 ;
        RECT 217.760 82.010 218.140 83.890 ;
        RECT 245.910 83.880 246.270 83.890 ;
        RECT 239.330 82.410 239.600 82.420 ;
        RECT 214.860 81.670 218.140 82.010 ;
        RECT 214.860 81.550 217.000 81.670 ;
        RECT 217.760 81.650 218.140 81.670 ;
        RECT 238.220 82.380 239.600 82.410 ;
        RECT 240.300 82.390 240.650 82.410 ;
        RECT 240.290 82.380 240.650 82.390 ;
        RECT 214.910 81.540 217.000 81.550 ;
        RECT 215.080 81.520 216.850 81.540 ;
        RECT 217.510 80.990 217.780 81.020 ;
        RECT 215.470 80.560 217.780 80.990 ;
        RECT 212.290 80.310 213.490 80.320 ;
        RECT 213.650 80.310 214.720 80.320 ;
        RECT 214.360 80.300 214.720 80.310 ;
        RECT 212.690 78.120 217.000 79.130 ;
        RECT 134.400 76.400 135.010 76.460 ;
        RECT 132.420 75.790 135.150 76.400 ;
        RECT 145.560 76.020 146.310 76.550 ;
        RECT 119.540 72.940 120.300 75.380 ;
        RECT 84.070 68.490 84.800 69.100 ;
        RECT 106.540 66.920 107.690 72.560 ;
        RECT 53.750 65.910 66.700 66.560 ;
        RECT 47.030 65.300 47.640 65.860 ;
        RECT 53.750 64.910 66.520 65.910 ;
        RECT 43.700 63.750 44.440 64.070 ;
        RECT 47.060 62.430 47.670 62.990 ;
        RECT 43.740 60.890 44.490 61.200 ;
        RECT 47.050 59.540 47.660 60.100 ;
        RECT 39.680 58.600 40.890 58.760 ;
        RECT 20.360 58.450 20.910 58.540 ;
        RECT 20.360 58.000 21.500 58.450 ;
        RECT 20.360 54.270 20.910 58.000 ;
        RECT 34.690 57.710 40.890 58.600 ;
        RECT 51.510 57.930 55.000 63.350 ;
        RECT 34.690 57.690 35.920 57.710 ;
        RECT 39.680 57.430 40.890 57.710 ;
        RECT 25.590 55.880 26.520 56.900 ;
        RECT 47.040 56.650 47.650 57.210 ;
        RECT 51.460 56.880 55.000 57.930 ;
        RECT 39.240 55.510 40.280 55.730 ;
        RECT 33.700 54.860 40.280 55.510 ;
        RECT 24.710 54.270 27.520 54.300 ;
        RECT 20.360 53.810 27.520 54.270 ;
        RECT 20.380 53.800 27.520 53.810 ;
        RECT 20.380 53.790 25.860 53.800 ;
        RECT 20.380 53.170 20.910 53.790 ;
        RECT 20.360 45.810 20.910 53.170 ;
        RECT 24.860 51.210 25.680 51.980 ;
        RECT 20.300 43.030 20.980 45.810 ;
        RECT 22.950 45.740 24.200 46.990 ;
        RECT 24.860 46.790 25.400 51.210 ;
        RECT 33.720 50.550 34.760 54.860 ;
        RECT 39.240 54.530 40.280 54.860 ;
        RECT 47.150 53.730 47.760 54.290 ;
        RECT 39.310 52.590 40.410 52.910 ;
        RECT 35.840 52.530 40.410 52.590 ;
        RECT 25.960 48.560 26.830 49.450 ;
        RECT 24.760 45.870 25.640 46.790 ;
        RECT 23.170 44.860 24.110 45.740 ;
        RECT 24.860 45.670 25.400 45.870 ;
        RECT 24.890 45.060 25.400 45.670 ;
        RECT 26.080 45.150 26.650 48.560 ;
        RECT 33.670 48.370 34.760 50.550 ;
        RECT 35.620 51.770 40.410 52.530 ;
        RECT 33.670 44.860 34.710 48.370 ;
        RECT 23.100 44.830 24.800 44.860 ;
        RECT 25.760 44.830 34.710 44.860 ;
        RECT 23.100 43.860 34.710 44.830 ;
        RECT 23.100 43.760 34.010 43.860 ;
        RECT 35.620 43.100 36.760 51.770 ;
        RECT 39.310 51.560 40.410 51.770 ;
        RECT 47.130 50.860 47.740 51.420 ;
        RECT 43.370 48.350 43.840 48.800 ;
        RECT 43.710 46.470 44.470 46.790 ;
        RECT 33.980 43.030 36.760 43.100 ;
        RECT 20.300 41.870 36.760 43.030 ;
        RECT 20.300 41.780 34.760 41.870 ;
        RECT 35.620 41.820 36.760 41.870 ;
        RECT 51.460 -2.890 54.840 56.880 ;
        RECT 63.320 53.710 64.650 59.540 ;
        RECT 83.970 55.140 118.640 55.430 ;
        RECT 119.530 55.140 120.300 72.940 ;
        RECT 83.970 54.510 120.300 55.140 ;
        RECT 134.400 55.340 135.010 75.790 ;
        RECT 145.540 75.480 146.310 76.020 ;
        RECT 134.400 54.980 135.140 55.340 ;
        RECT 145.540 55.300 146.240 75.480 ;
        RECT 152.810 71.910 153.960 77.710 ;
        RECT 217.510 76.450 217.780 80.560 ;
        RECT 238.220 80.410 240.650 82.380 ;
        RECT 240.790 81.640 242.930 82.410 ;
        RECT 240.840 81.630 242.930 81.640 ;
        RECT 241.010 81.610 242.780 81.630 ;
        RECT 241.400 80.980 243.700 81.080 ;
        RECT 245.940 80.980 246.170 81.000 ;
        RECT 241.400 80.780 246.170 80.980 ;
        RECT 241.400 80.650 243.700 80.780 ;
        RECT 238.220 80.400 239.420 80.410 ;
        RECT 239.580 80.400 240.650 80.410 ;
        RECT 240.290 80.390 240.650 80.400 ;
        RECT 245.940 79.390 246.170 80.780 ;
        RECT 261.810 79.510 262.460 85.230 ;
        RECT 265.210 82.470 265.480 82.480 ;
        RECT 264.100 82.440 265.480 82.470 ;
        RECT 266.180 82.450 266.530 82.470 ;
        RECT 266.170 82.440 266.530 82.450 ;
        RECT 264.100 80.470 266.530 82.440 ;
        RECT 266.670 81.700 268.810 82.470 ;
        RECT 266.720 81.690 268.810 81.700 ;
        RECT 266.890 81.670 268.660 81.690 ;
        RECT 269.310 81.140 269.600 81.150 ;
        RECT 267.280 80.710 269.600 81.140 ;
        RECT 264.100 80.460 265.300 80.470 ;
        RECT 265.460 80.460 266.530 80.470 ;
        RECT 266.170 80.450 266.530 80.460 ;
        RECT 247.060 79.390 247.850 79.490 ;
        RECT 245.940 79.220 247.850 79.390 ;
        RECT 238.620 78.210 242.930 79.220 ;
        RECT 245.950 79.190 247.850 79.220 ;
        RECT 247.060 79.090 247.850 79.190 ;
        RECT 261.810 79.090 262.480 79.510 ;
        RECT 259.880 77.660 261.230 78.600 ;
        RECT 261.830 77.130 262.480 79.090 ;
        RECT 264.500 78.270 268.810 79.280 ;
        RECT 269.310 77.340 269.600 80.710 ;
        RECT 275.350 78.940 276.000 85.640 ;
        RECT 295.140 82.880 295.820 83.420 ;
        RECT 290.630 82.010 291.320 82.790 ;
        RECT 333.320 82.690 337.100 83.580 ;
        RECT 293.490 81.430 293.760 81.440 ;
        RECT 292.380 81.400 293.760 81.430 ;
        RECT 294.460 81.410 294.810 81.430 ;
        RECT 294.450 81.400 294.810 81.410 ;
        RECT 292.380 79.430 294.810 81.400 ;
        RECT 294.950 80.660 297.090 81.430 ;
        RECT 295.000 80.650 297.090 80.660 ;
        RECT 295.170 80.630 296.940 80.650 ;
        RECT 295.560 79.670 297.860 80.100 ;
        RECT 292.380 79.420 293.580 79.430 ;
        RECT 293.740 79.420 294.810 79.430 ;
        RECT 294.450 79.410 294.810 79.420 ;
        RECT 275.350 78.170 276.020 78.940 ;
        RECT 264.190 77.130 265.030 77.180 ;
        RECT 218.390 76.450 218.990 76.630 ;
        RECT 260.100 76.500 260.990 76.930 ;
        RECT 261.830 76.590 265.030 77.130 ;
        RECT 217.510 76.240 218.990 76.450 ;
        RECT 217.520 76.200 218.990 76.240 ;
        RECT 218.390 76.050 218.990 76.200 ;
        RECT 261.000 75.610 261.880 76.050 ;
        RECT 235.190 71.140 238.170 72.160 ;
        RECT 261.010 69.740 261.740 70.160 ;
        RECT 264.190 66.780 265.030 76.590 ;
        RECT 269.320 74.500 269.580 77.340 ;
        RECT 271.690 74.500 272.980 74.700 ;
        RECT 269.310 74.230 272.980 74.500 ;
        RECT 275.370 74.340 276.020 78.170 ;
        RECT 292.780 77.230 297.090 78.240 ;
        RECT 288.580 75.950 289.680 76.330 ;
        RECT 297.590 75.950 297.850 79.670 ;
        RECT 304.700 76.400 305.300 76.780 ;
        RECT 288.580 75.610 297.860 75.950 ;
        RECT 344.430 75.720 353.200 75.780 ;
        RECT 288.580 75.400 289.680 75.610 ;
        RECT 342.210 74.850 353.730 75.720 ;
        RECT 355.190 74.850 381.510 74.870 ;
        RECT 269.320 68.470 269.580 74.230 ;
        RECT 271.690 74.130 272.980 74.230 ;
        RECT 275.260 73.580 276.670 74.340 ;
        RECT 275.950 69.150 276.560 73.580 ;
        RECT 289.860 73.250 290.450 73.410 ;
        RECT 342.210 73.280 381.510 74.850 ;
        RECT 331.260 73.250 381.510 73.280 ;
        RECT 289.860 73.070 381.510 73.250 ;
        RECT 289.860 73.050 359.670 73.070 ;
        RECT 289.860 73.030 355.610 73.050 ;
        RECT 289.860 72.930 353.730 73.030 ;
        RECT 289.860 72.900 331.620 72.930 ;
        RECT 289.860 72.780 290.450 72.900 ;
        RECT 342.210 72.150 353.730 72.930 ;
        RECT 344.430 72.130 353.200 72.150 ;
        RECT 344.550 72.070 347.660 72.130 ;
        RECT 464.420 70.510 471.520 126.110 ;
        RECT 495.550 124.280 496.260 131.600 ;
        RECT 493.020 119.180 496.260 124.280 ;
        RECT 534.420 132.060 552.270 133.410 ;
        RECT 576.300 132.980 581.250 134.320 ;
        RECT 534.420 124.740 548.000 132.060 ;
        RECT 551.670 124.740 552.270 132.060 ;
        RECT 579.780 125.660 581.250 132.980 ;
        RECT 534.420 120.580 552.270 124.740 ;
        RECT 483.520 109.220 484.660 109.850 ;
        RECT 481.720 81.590 487.350 81.740 ;
        RECT 481.120 78.020 488.170 81.590 ;
        RECT 481.060 75.690 488.170 78.020 ;
        RECT 490.190 76.480 496.260 119.180 ;
        RECT 522.260 109.760 524.140 110.600 ;
        RECT 512.280 108.560 515.690 109.690 ;
        RECT 538.080 108.910 541.370 110.040 ;
        RECT 546.200 76.480 552.270 120.580 ;
        RECT 576.300 119.020 581.250 125.660 ;
        RECT 567.120 108.480 569.800 109.350 ;
        RECT 481.060 72.120 488.110 75.690 ;
        RECT 268.800 67.440 269.940 68.470 ;
        RECT 264.190 66.430 269.070 66.780 ;
        RECT 145.540 55.270 180.230 55.300 ;
        RECT 83.970 54.480 120.150 54.510 ;
        RECT 83.970 54.180 118.640 54.480 ;
        RECT 131.300 54.250 135.190 54.980 ;
        RECT 145.540 54.910 181.280 55.270 ;
        RECT 143.480 54.320 181.280 54.910 ;
        RECT 131.300 54.170 132.020 54.250 ;
        RECT 134.450 51.600 135.140 54.250 ;
        RECT 145.540 54.110 181.280 54.320 ;
        RECT 145.560 54.050 181.280 54.110 ;
        RECT 179.400 54.000 181.280 54.050 ;
        RECT 84.050 50.610 135.440 51.600 ;
        RECT 85.100 42.660 85.880 43.760 ;
        RECT 106.550 42.400 107.690 47.810 ;
        RECT 118.880 45.880 119.860 46.980 ;
        RECT 57.710 2.800 59.620 36.160 ;
        RECT 119.100 25.970 119.830 45.880 ;
        RECT 119.100 25.810 119.820 25.970 ;
        RECT 132.660 25.890 133.860 47.230 ;
        RECT 136.850 25.890 138.480 25.980 ;
        RECT 122.660 25.810 124.380 25.850 ;
        RECT 119.060 25.680 124.380 25.810 ;
        RECT 118.210 24.940 124.380 25.680 ;
        RECT 132.660 25.550 138.480 25.890 ;
        RECT 119.060 24.850 124.380 24.940 ;
        RECT 106.280 19.940 108.840 22.640 ;
        RECT 122.660 19.910 124.380 24.850 ;
        RECT 131.250 24.760 138.480 25.550 ;
        RECT 131.250 24.700 133.860 24.760 ;
        RECT 122.660 18.440 129.630 19.910 ;
        RECT 136.850 19.660 138.480 24.760 ;
        RECT 145.170 24.730 146.370 47.260 ;
        RECT 151.960 31.310 153.840 44.340 ;
        RECT 203.190 41.510 204.300 53.240 ;
        RECT 268.310 51.620 269.030 66.430 ;
        RECT 275.870 57.010 276.610 69.150 ;
        RECT 464.400 67.890 471.520 70.510 ;
        RECT 464.400 62.810 471.410 67.890 ;
        RECT 490.080 67.550 552.730 76.480 ;
        RECT 574.150 69.940 581.250 119.020 ;
        RECT 574.150 67.430 581.410 69.940 ;
        RECT 574.400 62.810 581.410 67.430 ;
        RECT 455.030 57.630 457.310 59.250 ;
        RECT 275.870 56.980 286.910 57.010 ;
        RECT 293.970 56.980 296.640 57.220 ;
        RECT 275.870 56.230 296.640 56.980 ;
        RECT 463.370 56.250 582.220 62.810 ;
        RECT 286.430 56.090 296.640 56.230 ;
        RECT 293.970 53.110 296.640 56.090 ;
        RECT 574.400 55.910 581.410 56.250 ;
        RECT 268.260 49.000 269.170 51.620 ;
        RECT 268.350 47.260 269.120 49.000 ;
        RECT 282.510 47.430 307.090 47.480 ;
        RECT 310.250 47.430 311.420 47.570 ;
        RECT 282.510 47.260 311.420 47.430 ;
        RECT 268.350 46.600 311.420 47.260 ;
        RECT 282.510 46.560 311.420 46.600 ;
        RECT 306.710 46.490 311.420 46.560 ;
        RECT 141.740 19.660 147.220 19.740 ;
        RECT 136.850 18.280 147.220 19.660 ;
        RECT 141.740 18.250 147.220 18.280 ;
        RECT 143.110 3.210 144.570 4.490 ;
        RECT 123.320 2.920 162.740 3.000 ;
        RECT 85.410 2.800 162.740 2.920 ;
        RECT 57.540 1.940 162.740 2.800 ;
        RECT 57.540 1.900 162.720 1.940 ;
        RECT 57.540 1.820 124.810 1.900 ;
        RECT 57.540 1.700 94.250 1.820 ;
        RECT 57.710 1.530 59.620 1.700 ;
        RECT 203.120 -2.890 204.430 41.510 ;
        RECT 277.170 37.320 277.830 37.350 ;
        RECT 273.850 37.170 277.880 37.320 ;
        RECT 272.160 36.810 277.880 37.170 ;
        RECT 273.850 36.780 277.880 36.810 ;
        RECT 277.170 36.380 277.830 36.780 ;
        RECT 272.230 35.210 274.430 35.600 ;
        RECT 277.170 33.290 277.850 36.380 ;
        RECT 277.140 32.480 277.850 33.290 ;
        RECT 277.170 31.740 277.850 32.480 ;
        RECT 277.190 31.120 277.850 31.740 ;
        RECT 277.150 30.700 277.870 31.120 ;
        RECT 284.540 30.700 293.040 30.730 ;
        RECT 277.150 30.420 293.040 30.700 ;
        RECT 277.180 30.240 293.040 30.420 ;
        RECT 277.180 30.230 284.720 30.240 ;
        RECT 273.950 29.170 285.300 29.630 ;
        RECT 273.950 25.970 274.560 29.170 ;
        RECT 270.660 25.660 274.730 25.970 ;
        RECT 251.000 23.190 251.190 23.200 ;
        RECT 249.560 22.910 257.490 23.190 ;
        RECT 271.350 23.170 271.820 25.660 ;
        RECT 279.610 25.490 279.900 25.500 ;
        RECT 249.660 22.900 257.490 22.910 ;
        RECT 249.660 22.880 257.430 22.900 ;
        RECT 251.000 20.830 251.190 22.880 ;
        RECT 256.870 21.580 257.160 22.880 ;
        RECT 271.340 21.940 271.820 23.170 ;
        RECT 258.380 21.580 266.380 21.630 ;
        RECT 256.870 21.360 266.380 21.580 ;
        RECT 256.870 21.340 258.530 21.360 ;
        RECT 249.350 20.640 251.190 20.830 ;
        RECT 249.350 19.730 249.530 20.640 ;
        RECT 251.000 20.630 251.190 20.640 ;
        RECT 249.300 18.450 249.570 19.730 ;
        RECT 257.570 19.100 257.880 19.700 ;
        RECT 271.340 19.100 271.810 21.940 ;
        RECT 279.580 19.840 279.900 25.490 ;
        RECT 280.950 23.920 281.290 28.930 ;
        RECT 284.740 25.600 285.290 29.170 ;
        RECT 288.550 26.630 288.860 28.360 ;
        RECT 292.730 28.150 293.040 30.240 ;
        RECT 284.080 25.590 285.290 25.600 ;
        RECT 284.080 25.270 292.080 25.590 ;
        RECT 292.070 24.310 292.390 25.120 ;
        RECT 292.080 23.430 292.390 24.310 ;
        RECT 292.740 23.750 293.030 28.150 ;
        RECT 303.720 23.450 307.870 24.920 ;
        RECT 292.080 23.410 299.090 23.430 ;
        RECT 300.720 23.410 307.870 23.450 ;
        RECT 292.080 23.120 307.870 23.410 ;
        RECT 298.590 23.100 302.140 23.120 ;
        RECT 289.530 22.690 290.530 23.000 ;
        RECT 303.720 22.600 307.870 23.120 ;
        RECT 279.580 19.570 279.890 19.840 ;
        RECT 283.040 19.570 283.330 20.430 ;
        RECT 279.580 19.340 283.330 19.570 ;
        RECT 280.170 19.330 283.330 19.340 ;
        RECT 257.570 18.610 271.840 19.100 ;
        RECT 257.570 18.470 257.880 18.610 ;
        RECT 271.340 18.600 271.810 18.610 ;
        RECT 257.580 18.440 257.880 18.470 ;
        RECT 283.040 15.600 283.330 19.330 ;
        RECT 310.250 16.500 311.420 46.490 ;
        RECT 511.320 42.860 513.380 44.880 ;
        RECT 547.840 41.870 549.820 44.050 ;
        RECT 530.970 29.490 533.090 31.610 ;
        RECT 307.910 13.350 312.120 16.500 ;
        RECT 310.250 13.240 311.420 13.350 ;
        RECT 51.370 -9.180 204.540 -2.890 ;
        RECT 51.460 -9.350 54.840 -9.180 ;
      LAYER via2 ;
        RECT 174.440 160.440 174.810 160.800 ;
        RECT 167.740 157.520 168.040 157.830 ;
        RECT 173.090 155.590 173.460 155.920 ;
        RECT 64.720 124.870 66.220 125.800 ;
        RECT 22.460 69.010 23.090 69.780 ;
        RECT 25.940 61.510 26.460 62.110 ;
        RECT 44.530 71.730 44.900 72.180 ;
        RECT 47.210 71.340 47.620 71.750 ;
        RECT 43.690 69.720 44.300 70.000 ;
        RECT 47.110 68.260 47.520 68.670 ;
        RECT 39.750 66.500 40.560 67.150 ;
        RECT 43.510 66.660 44.250 66.940 ;
        RECT 134.970 133.570 135.900 134.530 ;
        RECT 155.730 133.310 156.470 133.800 ;
        RECT 177.050 133.080 177.650 133.580 ;
        RECT 341.430 132.270 342.140 132.910 ;
        RECT 337.440 131.360 338.320 132.030 ;
        RECT 331.950 128.730 332.910 129.100 ;
        RECT 344.300 127.590 345.010 128.230 ;
        RECT 588.580 204.410 590.500 206.180 ;
        RECT 475.330 200.940 476.700 201.600 ;
        RECT 549.240 194.610 554.820 198.570 ;
        RECT 467.580 163.660 468.390 164.020 ;
        RECT 576.600 195.800 580.890 199.740 ;
        RECT 497.060 163.850 497.870 164.210 ;
        RECT 551.520 163.890 552.330 164.250 ;
        RECT 447.780 146.900 448.290 148.500 ;
        RECT 475.230 148.110 476.050 150.870 ;
        RECT 530.520 150.500 531.070 152.430 ;
        RECT 577.870 163.510 578.680 163.870 ;
        RECT 558.090 148.240 558.490 150.490 ;
        RECT 396.260 120.040 397.200 120.920 ;
        RECT 407.750 121.180 408.750 122.350 ;
        RECT 468.180 109.840 468.990 110.200 ;
        RECT 492.810 110.190 493.620 110.550 ;
        RECT 456.470 108.840 457.010 109.160 ;
        RECT 106.730 90.060 107.970 91.180 ;
        RECT 244.060 88.900 244.750 89.530 ;
        RECT 290.930 89.850 291.640 90.130 ;
        RECT 84.260 68.680 84.640 68.960 ;
        RECT 47.140 65.370 47.550 65.780 ;
        RECT 54.140 65.220 54.560 66.100 ;
        RECT 47.170 62.490 47.580 62.900 ;
        RECT 53.660 62.370 54.430 63.170 ;
        RECT 43.800 60.910 44.420 61.190 ;
        RECT 47.150 59.620 47.560 60.030 ;
        RECT 25.770 56.160 26.290 56.760 ;
        RECT 47.160 56.710 47.570 57.120 ;
        RECT 63.800 58.690 64.310 59.300 ;
        RECT 47.260 53.800 47.670 54.210 ;
        RECT 26.120 48.680 26.730 49.280 ;
        RECT 23.170 45.890 24.000 46.790 ;
        RECT 47.240 50.920 47.650 51.330 ;
        RECT 43.440 48.420 43.750 48.740 ;
        RECT 43.770 46.480 44.400 46.760 ;
        RECT 63.480 54.040 64.330 54.930 ;
        RECT 260.010 77.830 261.020 78.440 ;
        RECT 295.240 82.970 295.710 83.340 ;
        RECT 333.580 82.890 333.860 83.410 ;
        RECT 336.570 82.950 336.850 83.470 ;
        RECT 290.760 82.160 291.170 82.660 ;
        RECT 260.260 76.580 260.860 76.860 ;
        RECT 261.130 75.700 261.750 75.980 ;
        RECT 236.990 71.450 237.660 71.780 ;
        RECT 261.080 69.800 261.670 70.110 ;
        RECT 288.720 75.550 289.510 76.140 ;
        RECT 304.770 76.450 305.230 76.730 ;
        RECT 289.950 72.920 290.340 73.310 ;
        RECT 483.700 109.330 484.240 109.650 ;
        RECT 522.500 109.900 523.820 110.380 ;
        RECT 512.980 108.720 515.070 109.610 ;
        RECT 538.660 109.070 540.750 109.960 ;
        RECT 549.160 109.450 549.970 109.810 ;
        RECT 576.780 109.890 577.590 110.250 ;
        RECT 567.340 108.590 569.630 109.230 ;
        RECT 482.590 73.030 485.100 74.800 ;
        RECT 85.230 42.890 85.750 43.240 ;
        RECT 58.170 34.870 58.940 35.460 ;
        RECT 106.780 20.740 108.250 22.050 ;
        RECT 465.740 64.820 469.280 69.480 ;
        RECT 545.280 68.790 551.090 74.370 ;
        RECT 455.580 57.880 456.910 58.810 ;
        RECT 143.460 3.440 144.060 4.160 ;
        RECT 162.050 2.200 162.500 2.720 ;
        RECT 272.330 35.250 274.350 35.540 ;
        RECT 280.990 23.990 281.270 28.870 ;
        RECT 288.560 26.690 288.840 28.310 ;
        RECT 289.610 22.700 290.450 22.980 ;
        RECT 304.730 22.890 306.530 23.850 ;
        RECT 511.730 43.190 513.050 44.530 ;
        RECT 548.260 42.320 549.410 43.530 ;
        RECT 531.330 29.900 532.760 31.250 ;
      LAYER met3 ;
        RECT 588.390 204.070 591.020 206.560 ;
        RECT 475.020 200.870 476.880 201.870 ;
        RECT 575.790 200.420 626.940 200.550 ;
        RECT 393.420 192.920 558.370 199.230 ;
        RECT 575.790 195.330 627.380 200.420 ;
        RECT 174.300 160.230 337.120 162.730 ;
        RECT 168.100 157.970 169.010 157.980 ;
        RECT 167.660 157.940 169.010 157.970 ;
        RECT 167.660 157.520 169.350 157.940 ;
        RECT 167.660 157.440 168.150 157.520 ;
        RECT 167.670 155.440 167.980 157.440 ;
        RECT 168.830 157.400 169.350 157.520 ;
        RECT 173.020 155.500 173.540 156.010 ;
        RECT 55.450 142.800 104.650 142.950 ;
        RECT 55.080 142.040 104.650 142.800 ;
        RECT 134.780 142.040 136.250 142.100 ;
        RECT 55.080 140.840 136.350 142.040 ;
        RECT 167.670 141.530 168.010 155.440 ;
        RECT 173.090 154.750 173.460 155.500 ;
        RECT 175.340 155.050 333.120 155.110 ;
        RECT 175.340 154.750 333.840 155.050 ;
        RECT 173.090 154.670 333.840 154.750 ;
        RECT 173.090 154.410 333.880 154.670 ;
        RECT 175.340 153.620 333.880 154.410 ;
        RECT 172.380 141.530 172.690 141.560 ;
        RECT 167.670 141.500 174.040 141.530 ;
        RECT 332.880 141.510 333.880 153.620 ;
        RECT 335.950 141.810 336.770 160.230 ;
        RECT 174.970 141.500 176.460 141.510 ;
        RECT 167.670 141.490 177.090 141.500 ;
        RECT 180.120 141.490 205.910 141.500 ;
        RECT 167.670 141.020 205.910 141.490 ;
        RECT 332.920 141.130 333.880 141.510 ;
        RECT 167.670 141.010 175.260 141.020 ;
        RECT 176.090 141.010 205.910 141.020 ;
        RECT 55.080 139.640 104.650 140.840 ;
        RECT 55.080 114.920 58.200 139.640 ;
        RECT 134.780 133.290 136.250 140.840 ;
        RECT 167.670 140.650 174.040 141.010 ;
        RECT 176.970 140.960 180.420 141.010 ;
        RECT 59.570 132.670 62.120 132.880 ;
        RECT 59.570 132.010 104.650 132.670 ;
        RECT 155.210 132.010 157.310 134.780 ;
        RECT 59.570 130.640 157.530 132.010 ;
        RECT 59.570 129.550 104.650 130.640 ;
        RECT 55.080 111.790 58.380 114.920 ;
        RECT 55.260 101.910 58.380 111.790 ;
        RECT 55.180 83.910 58.380 101.910 ;
        RECT 22.410 79.220 28.230 79.240 ;
        RECT 22.410 79.190 29.830 79.220 ;
        RECT 34.240 79.190 41.210 79.230 ;
        RECT 22.410 78.550 41.360 79.190 ;
        RECT 22.410 69.850 23.130 78.550 ;
        RECT 24.190 78.530 41.360 78.550 ;
        RECT 29.720 78.520 41.360 78.530 ;
        RECT 29.720 78.500 34.470 78.520 ;
        RECT 40.470 78.500 41.360 78.520 ;
        RECT 25.850 73.010 26.400 73.070 ;
        RECT 33.480 73.010 34.400 73.020 ;
        RECT 25.850 72.210 34.400 73.010 ;
        RECT 22.370 68.920 23.380 69.850 ;
        RECT 20.080 64.900 20.480 65.560 ;
        RECT 25.850 62.220 26.400 72.210 ;
        RECT 25.820 61.380 26.620 62.220 ;
        RECT 33.480 61.250 34.400 72.210 ;
        RECT 40.900 70.030 41.340 78.500 ;
        RECT 55.180 72.840 58.300 83.910 ;
        RECT 44.440 71.650 44.990 72.240 ;
        RECT 53.660 71.870 58.360 72.840 ;
        RECT 44.580 70.610 44.910 71.650 ;
        RECT 47.100 71.290 58.360 71.870 ;
        RECT 47.110 71.270 47.720 71.290 ;
        RECT 47.130 71.260 47.720 71.270 ;
        RECT 53.660 70.720 58.360 71.290 ;
        RECT 44.580 70.290 45.020 70.610 ;
        RECT 40.900 70.020 42.710 70.030 ;
        RECT 43.520 70.020 44.420 70.030 ;
        RECT 40.900 69.730 44.420 70.020 ;
        RECT 40.900 69.720 41.970 69.730 ;
        RECT 42.590 69.720 44.420 69.730 ;
        RECT 43.510 69.680 44.420 69.720 ;
        RECT 44.720 69.390 45.020 70.290 ;
        RECT 59.570 69.940 62.120 129.550 ;
        RECT 64.160 126.570 106.480 126.980 ;
        RECT 176.520 126.570 178.720 134.190 ;
        RECT 64.160 124.100 178.740 126.570 ;
        RECT 64.160 123.860 106.480 124.100 ;
        RECT 44.590 69.090 45.020 69.390 ;
        RECT 44.590 67.600 44.890 69.090 ;
        RECT 53.940 68.770 62.120 69.940 ;
        RECT 47.030 68.760 62.120 68.770 ;
        RECT 47.010 68.200 62.120 68.760 ;
        RECT 47.030 68.190 62.120 68.200 ;
        RECT 53.940 67.770 62.120 68.190 ;
        RECT 39.620 67.090 40.810 67.320 ;
        RECT 44.590 67.260 44.930 67.600 ;
        RECT 39.620 66.970 43.350 67.090 ;
        RECT 39.620 66.960 44.300 66.970 ;
        RECT 39.620 66.640 44.310 66.960 ;
        RECT 39.620 66.590 44.300 66.640 ;
        RECT 39.620 66.560 43.350 66.590 ;
        RECT 39.620 66.310 40.810 66.560 ;
        RECT 44.620 66.340 44.930 67.260 ;
        RECT 59.570 67.230 62.120 67.770 ;
        RECT 65.330 70.860 65.990 70.920 ;
        RECT 65.330 69.630 68.530 70.860 ;
        RECT 65.330 68.250 84.880 69.630 ;
        RECT 44.590 65.800 44.930 66.340 ;
        RECT 47.030 65.840 47.640 65.860 ;
        RECT 53.530 65.840 54.940 66.690 ;
        RECT 44.590 64.670 44.890 65.800 ;
        RECT 47.030 65.300 54.940 65.840 ;
        RECT 47.050 65.260 54.940 65.300 ;
        RECT 53.530 64.710 54.940 65.260 ;
        RECT 44.590 64.370 45.040 64.670 ;
        RECT 44.740 63.450 45.040 64.370 ;
        RECT 44.730 63.440 45.040 63.450 ;
        RECT 44.590 63.140 45.040 63.440 ;
        RECT 44.590 61.880 44.890 63.140 ;
        RECT 47.060 62.970 47.670 62.990 ;
        RECT 53.110 62.970 55.590 63.730 ;
        RECT 47.030 62.390 55.590 62.970 ;
        RECT 44.590 61.560 45.090 61.880 ;
        RECT 53.110 61.850 55.590 62.390 ;
        RECT 43.620 61.250 44.490 61.260 ;
        RECT 33.440 60.880 44.490 61.250 ;
        RECT 33.440 60.870 44.460 60.880 ;
        RECT 33.480 60.850 34.400 60.870 ;
        RECT 44.790 60.580 45.090 61.560 ;
        RECT 44.770 60.320 45.090 60.580 ;
        RECT 44.750 60.290 45.090 60.320 ;
        RECT 44.590 60.010 45.090 60.290 ;
        RECT 54.010 60.110 64.800 60.130 ;
        RECT 25.590 56.520 26.520 56.900 ;
        RECT 25.580 56.430 26.550 56.520 ;
        RECT 23.220 55.910 26.550 56.430 ;
        RECT 23.220 46.990 24.020 55.910 ;
        RECT 25.590 55.880 26.520 55.910 ;
        RECT 35.540 49.730 36.430 50.630 ;
        RECT 25.950 48.560 26.840 49.460 ;
        RECT 43.390 48.800 43.860 48.810 ;
        RECT 43.370 48.730 43.860 48.800 ;
        RECT 44.590 48.730 44.890 60.010 ;
        RECT 47.000 59.530 64.800 60.110 ;
        RECT 54.010 59.440 64.800 59.530 ;
        RECT 63.240 58.490 64.800 59.440 ;
        RECT 65.330 57.250 67.050 68.250 ;
        RECT 47.040 57.170 47.650 57.210 ;
        RECT 53.890 57.170 67.050 57.250 ;
        RECT 46.990 56.590 67.050 57.170 ;
        RECT 53.890 56.580 67.050 56.590 ;
        RECT 65.330 56.510 67.050 56.580 ;
        RECT 61.420 54.310 62.030 54.430 ;
        RECT 54.200 54.290 62.030 54.310 ;
        RECT 47.150 53.710 62.030 54.290 ;
        RECT 54.200 53.700 62.030 53.710 ;
        RECT 54.100 51.430 58.920 51.440 ;
        RECT 47.130 50.850 59.040 51.430 ;
        RECT 22.950 45.740 24.200 46.990 ;
        RECT 23.220 44.810 24.020 45.740 ;
        RECT 26.110 45.260 26.650 48.560 ;
        RECT 43.370 48.410 44.890 48.730 ;
        RECT 43.370 48.350 43.860 48.410 ;
        RECT 43.390 48.340 43.860 48.350 ;
        RECT 26.080 41.170 26.650 45.260 ;
        RECT 40.770 46.790 41.350 46.850 ;
        RECT 43.690 46.790 44.480 46.820 ;
        RECT 40.770 46.430 44.480 46.790 ;
        RECT 40.770 46.410 43.480 46.430 ;
        RECT 40.770 41.210 41.350 46.410 ;
        RECT 33.630 41.170 41.430 41.210 ;
        RECT 26.080 40.820 41.430 41.170 ;
        RECT 26.090 40.750 41.430 40.820 ;
        RECT 26.090 40.730 34.210 40.750 ;
        RECT 40.770 40.690 41.350 40.750 ;
        RECT 58.430 36.750 59.040 50.850 ;
        RECT 61.420 39.650 62.030 53.700 ;
        RECT 62.950 43.760 65.010 55.690 ;
        RECT 66.760 43.760 86.250 43.810 ;
        RECT 62.950 42.270 86.250 43.760 ;
        RECT 62.950 42.250 67.920 42.270 ;
        RECT 62.950 42.210 65.010 42.250 ;
        RECT 57.640 34.330 59.760 36.750 ;
        RECT 61.070 6.370 62.530 39.650 ;
        RECT 106.280 19.970 108.850 91.570 ;
        RECT 205.590 76.800 205.910 141.010 ;
        RECT 333.080 136.410 333.450 141.130 ;
        RECT 336.250 136.810 336.680 141.810 ;
        RECT 336.250 136.790 337.670 136.810 ;
        RECT 343.890 136.790 345.120 136.830 ;
        RECT 336.250 136.510 345.190 136.790 ;
        RECT 336.380 136.490 345.190 136.510 ;
        RECT 332.925 135.925 333.585 136.410 ;
        RECT 337.460 136.380 345.190 136.490 ;
        RECT 341.290 135.940 342.420 135.970 ;
        RECT 337.190 135.925 342.520 135.940 ;
        RECT 332.925 135.645 342.520 135.925 ;
        RECT 333.210 135.595 342.520 135.645 ;
        RECT 337.190 135.320 342.520 135.595 ;
        RECT 341.290 133.420 342.420 135.320 ;
        RECT 337.090 131.140 338.610 132.240 ;
        RECT 340.880 131.750 342.750 133.420 ;
        RECT 336.330 129.630 336.930 129.670 ;
        RECT 335.070 129.210 337.040 129.630 ;
        RECT 331.860 128.610 337.040 129.210 ;
        RECT 343.890 128.660 345.120 136.380 ;
        RECT 335.070 128.550 337.040 128.610 ;
        RECT 336.330 121.980 336.930 128.550 ;
        RECT 343.300 126.870 345.670 128.660 ;
        RECT 334.590 120.370 335.970 121.300 ;
        RECT 334.590 120.140 335.960 120.370 ;
        RECT 244.160 90.300 245.570 90.340 ;
        RECT 244.160 90.220 245.590 90.300 ;
        RECT 244.160 90.030 291.730 90.220 ;
        RECT 244.160 89.680 244.550 90.030 ;
        RECT 245.280 89.800 291.730 90.030 ;
        RECT 243.900 88.760 244.960 89.680 ;
        RECT 295.140 83.340 295.820 83.420 ;
        RECT 333.090 83.340 334.130 83.890 ;
        RECT 335.480 83.830 335.960 120.140 ;
        RECT 336.360 83.900 336.740 121.980 ;
        RECT 335.430 83.340 335.970 83.830 ;
        RECT 295.140 82.960 334.130 83.340 ;
        RECT 335.410 82.960 335.970 83.340 ;
        RECT 295.140 82.880 295.820 82.960 ;
        RECT 290.630 82.010 291.320 82.800 ;
        RECT 333.090 82.450 334.130 82.960 ;
        RECT 259.880 78.370 261.230 78.600 ;
        RECT 259.880 77.870 290.450 78.370 ;
        RECT 259.880 77.660 261.230 77.870 ;
        RECT 260.100 76.870 260.990 76.930 ;
        RECT 255.550 76.860 260.990 76.870 ;
        RECT 247.060 76.850 260.990 76.860 ;
        RECT 242.310 76.840 260.990 76.850 ;
        RECT 237.160 76.830 260.990 76.840 ;
        RECT 232.090 76.820 260.990 76.830 ;
        RECT 206.910 76.800 212.250 76.810 ;
        RECT 217.320 76.800 260.990 76.820 ;
        RECT 205.580 76.560 260.990 76.800 ;
        RECT 205.580 76.550 255.880 76.560 ;
        RECT 205.580 76.540 247.650 76.550 ;
        RECT 205.580 76.530 242.500 76.540 ;
        RECT 205.580 76.520 237.430 76.530 ;
        RECT 205.580 76.510 232.880 76.520 ;
        RECT 205.580 76.500 217.500 76.510 ;
        RECT 260.100 76.500 260.990 76.560 ;
        RECT 205.580 76.490 207.640 76.500 ;
        RECT 212.160 76.490 217.500 76.500 ;
        RECT 205.590 76.460 205.910 76.490 ;
        RECT 261.000 75.930 261.880 76.050 ;
        RECT 288.580 75.930 289.680 76.330 ;
        RECT 261.000 75.610 289.680 75.930 ;
        RECT 288.580 75.400 289.680 75.610 ;
        RECT 290.050 73.410 290.450 77.870 ;
        RECT 289.860 72.780 290.450 73.410 ;
        RECT 236.880 72.160 238.580 72.230 ;
        RECT 235.190 71.140 238.580 72.160 ;
        RECT 236.880 71.110 238.580 71.140 ;
        RECT 237.160 63.150 238.540 71.110 ;
        RECT 290.820 70.290 291.150 82.010 ;
        RECT 304.680 76.770 305.320 76.810 ;
        RECT 304.680 76.760 326.070 76.770 ;
        RECT 335.430 76.760 335.970 82.960 ;
        RECT 336.310 82.460 337.350 83.900 ;
        RECT 304.680 76.380 336.090 76.760 ;
        RECT 319.050 76.370 336.090 76.380 ;
        RECT 335.430 76.360 335.970 76.370 ;
        RECT 290.030 70.280 291.400 70.290 ;
        RECT 261.210 70.160 291.400 70.280 ;
        RECT 261.010 69.850 291.400 70.160 ;
        RECT 261.010 69.740 261.740 69.850 ;
        RECT 290.030 69.840 291.400 69.850 ;
        RECT 237.160 62.730 238.590 63.150 ;
        RECT 237.210 54.680 238.590 62.730 ;
        RECT 285.380 54.680 286.930 54.700 ;
        RECT 237.210 53.660 286.930 54.680 ;
        RECT 285.380 53.650 286.930 53.660 ;
        RECT 286.110 48.350 286.910 53.650 ;
        RECT 393.830 52.210 400.370 192.920 ;
        RECT 467.460 163.880 468.550 164.170 ;
        RECT 496.940 164.070 498.030 164.360 ;
        RECT 551.400 164.110 552.490 164.400 ;
        RECT 467.450 163.370 468.550 163.880 ;
        RECT 496.930 163.370 498.030 164.070 ;
        RECT 551.390 163.570 552.490 164.110 ;
        RECT 577.750 163.730 578.840 164.020 ;
        RECT 449.150 162.680 474.380 163.370 ;
        RECT 447.710 146.750 448.370 148.720 ;
        RECT 449.150 138.300 474.400 162.680 ;
        RECT 476.770 162.600 502.000 163.370 ;
        RECT 475.090 147.940 476.140 151.010 ;
        RECT 476.770 146.210 502.070 162.600 ;
        RECT 449.150 137.780 474.380 138.300 ;
        RECT 476.770 137.780 502.000 146.210 ;
        RECT 504.295 137.780 529.525 163.370 ;
        RECT 530.340 150.300 531.180 152.900 ;
        RECT 531.715 137.980 556.945 163.570 ;
        RECT 577.740 163.370 578.840 163.730 ;
        RECT 557.920 147.990 558.760 150.770 ;
        RECT 559.340 137.780 584.570 163.370 ;
        RECT 504.500 135.690 529.370 137.780 ;
        RECT 476.680 135.425 501.610 135.490 ;
        RECT 407.570 120.800 408.970 122.790 ;
        RECT 449.660 110.060 474.590 135.190 ;
        RECT 476.680 110.360 502.030 135.425 ;
        RECT 504.500 110.560 529.435 135.690 ;
        RECT 504.500 110.420 529.370 110.560 ;
        RECT 532.015 110.465 556.945 135.990 ;
        RECT 532.015 110.460 556.350 110.465 ;
        RECT 468.050 109.460 469.150 110.060 ;
        RECT 456.290 108.730 457.430 109.360 ;
        RECT 483.520 109.220 484.660 109.850 ;
        RECT 492.680 109.810 493.780 110.360 ;
        RECT 500.335 110.350 502.030 110.360 ;
        RECT 512.280 108.560 515.690 109.690 ;
        RECT 520.840 109.640 526.070 110.420 ;
        RECT 538.080 108.910 541.370 110.040 ;
        RECT 549.000 109.580 550.290 110.460 ;
        RECT 559.340 110.060 584.570 135.590 ;
        RECT 549.030 109.070 550.130 109.580 ;
        RECT 576.650 109.510 577.750 110.060 ;
        RECT 567.120 108.480 569.800 109.350 ;
        RECT 545.280 75.530 552.720 76.230 ;
        RECT 481.770 72.590 485.420 75.010 ;
        RECT 455.030 57.630 457.310 59.250 ;
        RECT 464.440 52.210 472.070 72.270 ;
        RECT 543.660 65.940 552.720 75.530 ;
        RECT 543.750 52.350 551.380 65.940 ;
        RECT 616.450 60.420 627.380 195.330 ;
        RECT 513.030 52.210 521.910 52.350 ;
        RECT 305.900 48.350 307.870 48.600 ;
        RECT 285.960 46.830 307.920 48.350 ;
        RECT 393.830 47.310 521.910 52.210 ;
        RECT 286.130 46.600 286.780 46.830 ;
        RECT 272.260 35.200 274.420 35.610 ;
        RECT 272.280 35.190 273.330 35.200 ;
        RECT 272.280 26.930 273.060 35.190 ;
        RECT 280.940 26.930 281.320 28.940 ;
        RECT 272.250 26.910 273.060 26.930 ;
        RECT 273.490 26.910 281.320 26.930 ;
        RECT 272.250 26.280 281.320 26.910 ;
        RECT 288.530 26.630 288.890 28.360 ;
        RECT 272.280 26.240 273.330 26.280 ;
        RECT 280.940 23.910 281.320 26.280 ;
        RECT 288.590 24.620 288.890 26.630 ;
        RECT 288.580 23.660 288.890 24.620 ;
        RECT 292.740 23.750 293.040 28.770 ;
        RECT 305.900 24.920 307.870 46.830 ;
        RECT 394.300 43.330 521.910 47.310 ;
        RECT 543.660 48.320 552.720 52.350 ;
        RECT 615.750 48.320 627.610 60.420 ;
        RECT 394.300 40.530 521.670 43.330 ;
        RECT 543.660 39.020 627.610 48.320 ;
        RECT 615.750 38.790 627.610 39.020 ;
        RECT 530.970 29.490 533.090 31.610 ;
        RECT 288.580 23.350 290.430 23.660 ;
        RECT 289.920 23.340 290.430 23.350 ;
        RECT 290.120 23.030 290.430 23.340 ;
        RECT 289.510 23.010 290.430 23.030 ;
        RECT 289.510 22.670 290.530 23.010 ;
        RECT 289.530 22.650 290.530 22.670 ;
        RECT 303.720 22.600 307.870 24.920 ;
        RECT 60.560 4.490 62.620 6.370 ;
        RECT 60.560 4.480 101.470 4.490 ;
        RECT 143.110 4.480 144.570 4.490 ;
        RECT 60.560 2.770 144.890 4.480 ;
        RECT 60.560 2.600 101.470 2.770 ;
        RECT 161.880 1.940 162.740 3.000 ;
      LAYER via3 ;
        RECT 588.580 204.410 590.500 206.180 ;
        RECT 475.330 200.940 476.700 201.600 ;
        RECT 337.400 131.320 338.370 132.040 ;
        RECT 335.100 120.560 335.550 120.910 ;
        RECT 447.830 146.930 448.250 148.480 ;
        RECT 475.230 148.110 476.050 150.870 ;
        RECT 530.520 150.500 531.070 152.430 ;
        RECT 558.090 148.240 558.490 150.490 ;
        RECT 407.750 121.180 408.750 122.350 ;
        RECT 483.700 109.330 484.240 109.650 ;
        RECT 456.470 108.840 457.010 109.160 ;
        RECT 512.980 108.720 515.070 109.610 ;
        RECT 538.660 109.070 540.750 109.960 ;
        RECT 567.340 108.590 569.630 109.230 ;
        RECT 482.590 73.030 485.100 74.800 ;
        RECT 455.580 57.880 456.910 58.810 ;
        RECT 531.330 29.900 532.760 31.250 ;
      LAYER met4 ;
        RECT 608.540 207.510 644.150 207.630 ;
        RECT 560.590 202.510 644.150 207.510 ;
        RECT 560.590 202.290 611.740 202.510 ;
        RECT 625.750 202.050 644.150 202.510 ;
        RECT 405.980 199.230 412.520 199.460 ;
        RECT 471.500 199.230 477.440 201.960 ;
        RECT 405.660 192.680 477.440 199.230 ;
        RECT 337.090 132.060 338.610 132.240 ;
        RECT 334.990 131.420 338.650 132.060 ;
        RECT 335.020 120.420 335.620 131.420 ;
        RECT 337.090 131.140 338.610 131.420 ;
        RECT 405.980 64.870 412.520 192.680 ;
        RECT 471.500 192.620 477.440 192.680 ;
        RECT 451.200 151.110 460.450 161.460 ;
        RECT 480.880 160.080 488.295 161.385 ;
        RECT 480.440 152.510 488.295 160.080 ;
        RECT 535.320 155.890 544.000 161.660 ;
        RECT 530.640 153.340 544.000 155.890 ;
        RECT 561.320 154.270 570.700 162.620 ;
        RECT 475.790 152.480 488.295 152.510 ;
        RECT 475.220 152.070 488.295 152.480 ;
        RECT 447.530 144.500 460.450 151.110 ;
        RECT 474.960 148.590 488.295 152.070 ;
        RECT 530.060 149.550 544.000 153.340 ;
        RECT 474.960 147.285 487.855 148.590 ;
        RECT 474.960 147.160 482.350 147.285 ;
        RECT 475.220 146.930 482.350 147.160 ;
        RECT 475.220 146.900 481.780 146.930 ;
        RECT 447.530 144.300 457.550 144.500 ;
        RECT 447.530 144.290 448.550 144.300 ;
        RECT 509.190 137.430 522.400 148.790 ;
        RECT 530.640 147.530 544.000 149.550 ;
        RECT 535.320 147.440 544.000 147.530 ;
        RECT 557.880 144.880 570.700 154.270 ;
        RECT 557.880 144.600 564.550 144.880 ;
        RECT 509.190 135.510 521.630 137.430 ;
        RECT 450.520 123.960 462.390 135.010 ;
        RECT 509.190 134.070 522.400 135.510 ;
        RECT 451.190 118.440 462.370 123.960 ;
        RECT 480.560 123.600 489.470 133.910 ;
        RECT 509.190 133.180 521.520 134.070 ;
        RECT 508.930 133.030 521.520 133.180 ;
        RECT 480.310 123.100 489.470 123.600 ;
        RECT 480.310 119.080 489.220 123.100 ;
        RECT 508.780 122.790 521.600 133.030 ;
        RECT 452.840 108.970 462.000 118.440 ;
        RECT 480.060 112.790 489.220 119.080 ;
        RECT 455.190 108.590 458.820 108.970 ;
        RECT 480.060 108.880 489.210 112.790 ;
        RECT 509.600 110.670 520.690 122.790 ;
        RECT 535.660 119.140 545.590 134.040 ;
        RECT 564.390 121.440 573.420 132.420 ;
        RECT 509.130 108.320 520.780 110.670 ;
        RECT 535.490 109.350 545.630 119.140 ;
        RECT 536.400 108.370 543.250 109.350 ;
        RECT 565.060 108.350 572.100 121.440 ;
        RECT 566.250 108.340 570.990 108.350 ;
        RECT 480.530 81.260 488.550 81.910 ;
        RECT 480.530 77.340 482.530 81.260 ;
        RECT 486.960 77.340 488.550 81.260 ;
        RECT 480.530 73.270 488.550 77.340 ;
        RECT 480.630 66.930 488.540 73.270 ;
        RECT 404.510 56.530 413.030 64.870 ;
        RECT 452.290 60.160 461.100 60.200 ;
        RECT 445.360 56.530 461.100 60.160 ;
        RECT 404.510 53.320 461.100 56.530 ;
        RECT 404.510 52.920 460.910 53.320 ;
        RECT 404.510 47.370 413.030 52.920 ;
        RECT 480.630 42.510 488.070 66.930 ;
        RECT 479.700 35.770 488.070 42.510 ;
        RECT 632.260 35.770 643.890 202.050 ;
        RECT 479.700 27.390 643.890 35.770 ;
        RECT 632.260 26.700 643.890 27.390 ;
  END
END analog_macro
END LIBRARY

