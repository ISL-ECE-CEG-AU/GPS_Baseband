magic
tech sky130A
magscale 1 2
timestamp 1637989401
<< locali >>
rect 544761 668423 544795 670361
rect 139811 643297 140237 643331
rect 183235 643297 183569 643331
rect 188353 638503 188387 645609
rect 188445 638367 188479 645881
rect 196357 642379 196391 645541
rect 196541 645167 196575 645881
rect 199853 640747 199887 645881
rect 475669 644895 475703 645813
rect 427035 643501 427461 643535
rect 429393 643399 429427 643977
rect 225797 643331 225831 643365
rect 433073 643331 433107 643977
rect 225797 643297 226441 643331
rect 233375 643297 233801 643331
rect 443653 643195 443687 644453
rect 476957 643331 476991 643841
rect 476957 643297 477509 643331
rect 189917 639557 190285 639591
rect 191055 639557 191297 639591
rect 189825 638979 189859 639489
rect 189917 639115 189951 639557
rect 190043 639489 190377 639523
rect 190963 639489 191389 639523
rect 190009 639421 190285 639455
rect 191055 639421 191297 639455
rect 190009 639047 190043 639421
rect 196357 635171 196391 635613
rect 58207 633369 58633 633403
rect 117823 632689 118433 632723
rect 198473 632519 198507 633981
rect 199577 632519 199611 633981
rect 201969 632247 202003 633709
rect 212457 631431 212491 631737
rect 139811 631397 140237 631431
rect 196115 631397 196357 631431
rect 214113 629323 214147 632757
rect 217793 629119 217827 635953
rect 441537 630819 441571 631737
rect 477049 630785 477509 630819
rect 477049 630683 477083 630785
rect 224911 630649 225153 630683
rect 228591 630649 228925 630683
rect 405691 630649 405783 630683
rect 462087 630649 462421 630683
rect 197369 628881 197478 628915
rect 197369 627963 197403 628881
rect 214113 628235 214147 629085
rect 405749 628983 405783 630649
rect 218897 620007 218931 627725
rect 545773 619871 545807 623033
rect 137109 618307 137143 618885
rect 138489 618579 138523 618953
rect 138489 618545 139041 618579
rect 137327 617049 137661 617083
rect 138523 617049 139041 617083
rect 146803 617049 147505 617083
rect 98653 577575 98687 577949
rect 145607 577473 146309 577507
rect 152047 577473 152749 577507
rect 158763 577473 159465 577507
rect 195621 313055 195655 313157
rect 39129 309927 39163 310165
rect 41337 309179 41371 310165
rect 46397 309247 46431 310165
rect 48789 309315 48823 310165
rect 55965 309383 55999 310233
rect 60657 309451 60691 310301
rect 63233 309519 63267 310301
rect 70317 309587 70351 310301
rect 269681 309859 269715 309961
rect 274649 309791 274683 309961
rect 296177 309723 296211 309961
rect 114845 31399 114879 31569
rect 94421 30991 94455 31161
rect 127449 30651 127483 31365
rect 179337 30515 179371 30753
rect 200589 30379 200623 30889
rect 238769 30583 238803 31433
rect 270141 30617 270601 30651
rect 269439 30549 269773 30583
rect 239505 30379 239539 30549
rect 270141 30515 270175 30617
rect 248245 30379 248279 30481
rect 283239 9333 283389 9367
rect 286885 9299 286919 9469
rect 286827 9265 286919 9299
rect 300627 8993 300961 9027
rect 218161 4199 218195 4505
rect 26249 3723 26283 3893
rect 103897 3859 103931 4165
rect 108221 3859 108255 4029
rect 111533 3995 111567 4165
rect 272349 4199 272383 4641
rect 272441 4403 272475 4709
rect 272533 4471 272567 4641
rect 272625 4267 272659 4437
rect 272567 4233 272659 4267
rect 272717 4267 272751 4573
rect 272809 4471 272843 4573
rect 272901 4471 272935 4981
rect 281917 4607 281951 5185
rect 282009 4607 282043 4913
rect 282193 4675 282227 4845
rect 282377 4539 282411 4981
rect 282469 4539 282503 5049
rect 282561 4607 282595 5117
rect 301421 5049 301639 5083
rect 301421 5015 301455 5049
rect 301513 4811 301547 4981
rect 301605 4811 301639 5049
rect 272349 4165 272809 4199
rect 368857 4165 369075 4199
rect 26433 3519 26467 3825
rect 108129 3825 108255 3859
rect 62129 3451 62163 3757
rect 71697 3383 71731 3825
rect 108129 3791 108163 3825
rect 88901 3689 89269 3723
rect 87521 3315 87555 3621
rect 88901 3519 88935 3689
rect 90465 3315 90499 3485
rect 104081 3383 104115 3757
rect 87521 3281 88073 3315
rect 90407 3281 90499 3315
rect 104541 2975 104575 3213
rect 108221 2975 108255 3757
rect 108313 3383 108347 3825
rect 111717 3791 111751 3961
rect 111809 3927 111843 4029
rect 111901 3859 111935 4029
rect 118065 3995 118099 4165
rect 368857 4131 368891 4165
rect 111993 3247 112027 3825
rect 117881 3315 117915 3893
rect 117973 3519 118007 3757
rect 104541 2941 105001 2975
rect 118065 3247 118099 3825
rect 121193 3519 121227 3961
rect 127541 3791 127575 3961
rect 127449 3451 127483 3757
rect 127725 3519 127759 4029
rect 132049 3519 132083 3689
rect 127817 3451 127851 3485
rect 127449 3417 127851 3451
rect 185685 3315 185719 3349
rect 185535 3281 185719 3315
rect 108313 2975 108347 3213
rect 178141 2839 178175 3213
rect 178233 2839 178267 3077
rect 194241 3043 194275 3281
rect 186271 2941 186513 2975
rect 194333 2907 194367 3009
rect 195161 2907 195195 3213
rect 195437 3179 195471 3213
rect 195287 3145 195471 3179
rect 196909 2907 196943 4097
rect 200129 3723 200163 3961
rect 200589 3383 200623 3621
rect 205005 3315 205039 3893
rect 320649 2771 320683 3077
rect 320741 2975 320775 3077
rect 320833 2839 320867 2941
rect 333161 2771 333195 3009
rect 344201 2839 344235 3145
rect 344661 2907 344695 3213
rect 349077 3043 349111 3281
rect 349813 3043 349847 3213
rect 349721 2975 349755 3009
rect 349905 2975 349939 3213
rect 349721 2941 349939 2975
rect 355885 2907 355919 3349
rect 368949 3247 368983 4097
rect 369041 3451 369075 4165
rect 382933 4165 383611 4199
rect 369041 3417 369351 3451
rect 369133 3043 369167 3145
rect 369225 3043 369259 3349
rect 369317 3247 369351 3417
rect 373089 3383 373123 4097
rect 382933 3995 382967 4165
rect 383577 4131 383611 4165
rect 383427 4029 383669 4063
rect 382875 3961 382967 3995
rect 369317 3213 369501 3247
rect 583401 3111 583435 6137
rect 344753 2839 344787 2873
rect 334023 2805 334173 2839
rect 344201 2805 344787 2839
rect 355735 2805 355977 2839
rect 358863 2805 359013 2839
<< viali >>
rect 544761 670361 544795 670395
rect 544761 668389 544795 668423
rect 226165 646017 226199 646051
rect 188445 645881 188479 645915
rect 188353 645609 188387 645643
rect 139777 643297 139811 643331
rect 140237 643297 140271 643331
rect 183201 643297 183235 643331
rect 183569 643297 183603 643331
rect 188353 638469 188387 638503
rect 196541 645881 196575 645915
rect 196357 645541 196391 645575
rect 196541 645133 196575 645167
rect 199853 645881 199887 645915
rect 196357 642345 196391 642379
rect 475669 645813 475703 645847
rect 475669 644861 475703 644895
rect 443653 644453 443687 644487
rect 429393 643977 429427 644011
rect 427001 643501 427035 643535
rect 427461 643501 427495 643535
rect 225797 643365 225831 643399
rect 429393 643365 429427 643399
rect 433073 643977 433107 644011
rect 226441 643297 226475 643331
rect 233341 643297 233375 643331
rect 233801 643297 233835 643331
rect 433073 643297 433107 643331
rect 476957 643841 476991 643875
rect 477509 643297 477543 643331
rect 443653 643161 443687 643195
rect 199853 640713 199887 640747
rect 190285 639557 190319 639591
rect 191021 639557 191055 639591
rect 191297 639557 191331 639591
rect 189825 639489 189859 639523
rect 190009 639489 190043 639523
rect 190377 639489 190411 639523
rect 190929 639489 190963 639523
rect 191389 639489 191423 639523
rect 189917 639081 189951 639115
rect 190285 639421 190319 639455
rect 191021 639421 191055 639455
rect 191297 639421 191331 639455
rect 190009 639013 190043 639047
rect 189825 638945 189859 638979
rect 188445 638333 188479 638367
rect 217793 635953 217827 635987
rect 196357 635613 196391 635647
rect 196357 635137 196391 635171
rect 198473 633981 198507 634015
rect 58173 633369 58207 633403
rect 58633 633369 58667 633403
rect 117789 632689 117823 632723
rect 118433 632689 118467 632723
rect 198473 632485 198507 632519
rect 199577 633981 199611 634015
rect 199577 632485 199611 632519
rect 201969 633709 202003 633743
rect 201969 632213 202003 632247
rect 214113 632757 214147 632791
rect 212457 631737 212491 631771
rect 139777 631397 139811 631431
rect 140237 631397 140271 631431
rect 196081 631397 196115 631431
rect 196357 631397 196391 631431
rect 212457 631397 212491 631431
rect 214113 629289 214147 629323
rect 441537 631737 441571 631771
rect 441537 630785 441571 630819
rect 477509 630785 477543 630819
rect 224877 630649 224911 630683
rect 225153 630649 225187 630683
rect 228557 630649 228591 630683
rect 228925 630649 228959 630683
rect 405657 630649 405691 630683
rect 462053 630649 462087 630683
rect 462421 630649 462455 630683
rect 477049 630649 477083 630683
rect 214113 629085 214147 629119
rect 217793 629085 217827 629119
rect 405749 628949 405783 628983
rect 214113 628201 214147 628235
rect 197369 627929 197403 627963
rect 218897 627725 218931 627759
rect 218897 619973 218931 620007
rect 545773 623033 545807 623067
rect 545773 619837 545807 619871
rect 138489 618953 138523 618987
rect 137109 618885 137143 618919
rect 139041 618545 139075 618579
rect 137109 618273 137143 618307
rect 137293 617049 137327 617083
rect 137661 617049 137695 617083
rect 138489 617049 138523 617083
rect 139041 617049 139075 617083
rect 146769 617049 146803 617083
rect 147505 617049 147539 617083
rect 98653 577949 98687 577983
rect 98653 577541 98687 577575
rect 145573 577473 145607 577507
rect 146309 577473 146343 577507
rect 152013 577473 152047 577507
rect 152749 577473 152783 577507
rect 158729 577473 158763 577507
rect 159465 577473 159499 577507
rect 195621 313157 195655 313191
rect 195621 313021 195655 313055
rect 60657 310301 60691 310335
rect 55965 310233 55999 310267
rect 39129 310165 39163 310199
rect 39129 309893 39163 309927
rect 41337 310165 41371 310199
rect 46397 310165 46431 310199
rect 48789 310165 48823 310199
rect 63233 310301 63267 310335
rect 70317 310301 70351 310335
rect 269681 309961 269715 309995
rect 269681 309825 269715 309859
rect 274649 309961 274683 309995
rect 274649 309757 274683 309791
rect 296177 309961 296211 309995
rect 296177 309689 296211 309723
rect 70317 309553 70351 309587
rect 63233 309485 63267 309519
rect 60657 309417 60691 309451
rect 55965 309349 55999 309383
rect 48789 309281 48823 309315
rect 46397 309213 46431 309247
rect 41337 309145 41371 309179
rect 114845 31569 114879 31603
rect 238769 31433 238803 31467
rect 114845 31365 114879 31399
rect 127449 31365 127483 31399
rect 94421 31161 94455 31195
rect 94421 30957 94455 30991
rect 200589 30889 200623 30923
rect 127449 30617 127483 30651
rect 179337 30753 179371 30787
rect 179337 30481 179371 30515
rect 270601 30617 270635 30651
rect 238769 30549 238803 30583
rect 239505 30549 239539 30583
rect 269405 30549 269439 30583
rect 269773 30549 269807 30583
rect 200589 30345 200623 30379
rect 239505 30345 239539 30379
rect 248245 30481 248279 30515
rect 270141 30481 270175 30515
rect 248245 30345 248279 30379
rect 286885 9469 286919 9503
rect 283205 9333 283239 9367
rect 283389 9333 283423 9367
rect 286793 9265 286827 9299
rect 300593 8993 300627 9027
rect 300961 8993 300995 9027
rect 583401 6137 583435 6171
rect 281917 5185 281951 5219
rect 272901 4981 272935 5015
rect 272441 4709 272475 4743
rect 272349 4641 272383 4675
rect 218161 4505 218195 4539
rect 103897 4165 103931 4199
rect 26249 3893 26283 3927
rect 111533 4165 111567 4199
rect 108221 4029 108255 4063
rect 118065 4165 118099 4199
rect 218161 4165 218195 4199
rect 272533 4641 272567 4675
rect 272717 4573 272751 4607
rect 272533 4437 272567 4471
rect 272625 4437 272659 4471
rect 272441 4369 272475 4403
rect 272533 4233 272567 4267
rect 272809 4573 272843 4607
rect 272809 4437 272843 4471
rect 282561 5117 282595 5151
rect 282469 5049 282503 5083
rect 282377 4981 282411 5015
rect 281917 4573 281951 4607
rect 282009 4913 282043 4947
rect 282193 4845 282227 4879
rect 282193 4641 282227 4675
rect 282009 4573 282043 4607
rect 282377 4505 282411 4539
rect 301421 4981 301455 5015
rect 301513 4981 301547 5015
rect 301513 4777 301547 4811
rect 301605 4777 301639 4811
rect 282561 4573 282595 4607
rect 282469 4505 282503 4539
rect 272901 4437 272935 4471
rect 272717 4233 272751 4267
rect 272809 4165 272843 4199
rect 111809 4029 111843 4063
rect 111533 3961 111567 3995
rect 111717 3961 111751 3995
rect 26249 3689 26283 3723
rect 26433 3825 26467 3859
rect 71697 3825 71731 3859
rect 103897 3825 103931 3859
rect 108313 3825 108347 3859
rect 26433 3485 26467 3519
rect 62129 3757 62163 3791
rect 62129 3417 62163 3451
rect 104081 3757 104115 3791
rect 108129 3757 108163 3791
rect 108221 3757 108255 3791
rect 89269 3689 89303 3723
rect 71697 3349 71731 3383
rect 87521 3621 87555 3655
rect 88901 3485 88935 3519
rect 90465 3485 90499 3519
rect 104081 3349 104115 3383
rect 88073 3281 88107 3315
rect 90373 3281 90407 3315
rect 104541 3213 104575 3247
rect 111809 3893 111843 3927
rect 111901 4029 111935 4063
rect 196909 4097 196943 4131
rect 368857 4097 368891 4131
rect 368949 4097 368983 4131
rect 127725 4029 127759 4063
rect 118065 3961 118099 3995
rect 121193 3961 121227 3995
rect 117881 3893 117915 3927
rect 111901 3825 111935 3859
rect 111993 3825 112027 3859
rect 111717 3757 111751 3791
rect 108313 3349 108347 3383
rect 118065 3825 118099 3859
rect 117973 3757 118007 3791
rect 117973 3485 118007 3519
rect 117881 3281 117915 3315
rect 105001 2941 105035 2975
rect 108221 2941 108255 2975
rect 108313 3213 108347 3247
rect 111993 3213 112027 3247
rect 127541 3961 127575 3995
rect 121193 3485 121227 3519
rect 127449 3757 127483 3791
rect 127541 3757 127575 3791
rect 132049 3689 132083 3723
rect 127725 3485 127759 3519
rect 127817 3485 127851 3519
rect 132049 3485 132083 3519
rect 185685 3349 185719 3383
rect 185501 3281 185535 3315
rect 194241 3281 194275 3315
rect 118065 3213 118099 3247
rect 178141 3213 178175 3247
rect 108313 2941 108347 2975
rect 178141 2805 178175 2839
rect 178233 3077 178267 3111
rect 195161 3213 195195 3247
rect 194241 3009 194275 3043
rect 194333 3009 194367 3043
rect 186237 2941 186271 2975
rect 186513 2941 186547 2975
rect 194333 2873 194367 2907
rect 195437 3213 195471 3247
rect 195253 3145 195287 3179
rect 195161 2873 195195 2907
rect 200129 3961 200163 3995
rect 200129 3689 200163 3723
rect 205005 3893 205039 3927
rect 200589 3621 200623 3655
rect 200589 3349 200623 3383
rect 355885 3349 355919 3383
rect 205005 3281 205039 3315
rect 349077 3281 349111 3315
rect 344661 3213 344695 3247
rect 344201 3145 344235 3179
rect 196909 2873 196943 2907
rect 320649 3077 320683 3111
rect 178233 2805 178267 2839
rect 320741 3077 320775 3111
rect 333161 3009 333195 3043
rect 320741 2941 320775 2975
rect 320833 2941 320867 2975
rect 320833 2805 320867 2839
rect 320649 2737 320683 2771
rect 349813 3213 349847 3247
rect 349077 3009 349111 3043
rect 349721 3009 349755 3043
rect 349813 3009 349847 3043
rect 349905 3213 349939 3247
rect 373089 4097 373123 4131
rect 368949 3213 368983 3247
rect 369225 3349 369259 3383
rect 369133 3145 369167 3179
rect 369133 3009 369167 3043
rect 383577 4097 383611 4131
rect 383393 4029 383427 4063
rect 383669 4029 383703 4063
rect 382841 3961 382875 3995
rect 373089 3349 373123 3383
rect 369501 3213 369535 3247
rect 583401 3077 583435 3111
rect 369225 3009 369259 3043
rect 344661 2873 344695 2907
rect 344753 2873 344787 2907
rect 355885 2873 355919 2907
rect 333989 2805 334023 2839
rect 334173 2805 334207 2839
rect 355701 2805 355735 2839
rect 355977 2805 356011 2839
rect 358829 2805 358863 2839
rect 359013 2805 359047 2839
rect 333161 2737 333195 2771
<< metal1 >>
rect 24302 700952 24308 701004
rect 24360 700992 24366 701004
rect 196342 700992 196348 701004
rect 24360 700964 196348 700992
rect 24360 700952 24366 700964
rect 196342 700952 196348 700964
rect 196400 700952 196406 701004
rect 8110 700884 8116 700936
rect 8168 700924 8174 700936
rect 188982 700924 188988 700936
rect 8168 700896 188988 700924
rect 8168 700884 8174 700896
rect 188982 700884 188988 700896
rect 189040 700884 189046 700936
rect 164142 700816 164148 700868
rect 164200 700856 164206 700868
rect 348786 700856 348792 700868
rect 164200 700828 348792 700856
rect 164200 700816 164206 700828
rect 348786 700816 348792 700828
rect 348844 700816 348850 700868
rect 40494 700748 40500 700800
rect 40552 700788 40558 700800
rect 227714 700788 227720 700800
rect 40552 700760 227720 700788
rect 40552 700748 40558 700760
rect 227714 700748 227720 700760
rect 227772 700748 227778 700800
rect 154482 700680 154488 700732
rect 154540 700720 154546 700732
rect 397454 700720 397460 700732
rect 154540 700692 397460 700720
rect 154540 700680 154546 700692
rect 397454 700680 397460 700692
rect 397512 700680 397518 700732
rect 157242 700612 157248 700664
rect 157300 700652 157306 700664
rect 413646 700652 413652 700664
rect 157300 700624 413652 700652
rect 157300 700612 157306 700624
rect 413646 700612 413652 700624
rect 413704 700612 413710 700664
rect 148318 700544 148324 700596
rect 148376 700584 148382 700596
rect 462314 700584 462320 700596
rect 148376 700556 462320 700584
rect 148376 700544 148382 700556
rect 462314 700544 462320 700556
rect 462372 700544 462378 700596
rect 150342 700476 150348 700528
rect 150400 700516 150406 700528
rect 478506 700516 478512 700528
rect 150400 700488 478512 700516
rect 150400 700476 150406 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 144822 700408 144828 700460
rect 144880 700448 144886 700460
rect 494790 700448 494796 700460
rect 144880 700420 494796 700448
rect 144880 700408 144886 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 140682 700340 140688 700392
rect 140740 700380 140746 700392
rect 527174 700380 527180 700392
rect 140740 700352 527180 700380
rect 140740 700340 140746 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 98638 700312 98644 700324
rect 89220 700284 98644 700312
rect 89220 700272 89226 700284
rect 98638 700272 98644 700284
rect 98696 700272 98702 700324
rect 137094 700272 137100 700324
rect 137152 700312 137158 700324
rect 559650 700312 559656 700324
rect 137152 700284 559656 700312
rect 137152 700272 137158 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 162762 700204 162768 700256
rect 162820 700244 162826 700256
rect 332502 700244 332508 700256
rect 162820 700216 332508 700244
rect 162820 700204 162826 700216
rect 332502 700204 332508 700216
rect 332560 700204 332566 700256
rect 72970 700136 72976 700188
rect 73028 700176 73034 700188
rect 188338 700176 188344 700188
rect 73028 700148 188344 700176
rect 73028 700136 73034 700148
rect 188338 700136 188344 700148
rect 188396 700136 188402 700188
rect 188430 700136 188436 700188
rect 188488 700176 188494 700188
rect 218974 700176 218980 700188
rect 188488 700148 218980 700176
rect 188488 700136 188494 700148
rect 218974 700136 218980 700148
rect 219032 700136 219038 700188
rect 172422 700068 172428 700120
rect 172480 700108 172486 700120
rect 283834 700108 283840 700120
rect 172480 700080 283840 700108
rect 172480 700068 172486 700080
rect 283834 700068 283840 700080
rect 283892 700068 283898 700120
rect 169662 700000 169668 700052
rect 169720 700040 169726 700052
rect 267642 700040 267648 700052
rect 169720 700012 267648 700040
rect 169720 700000 169726 700012
rect 267642 700000 267648 700012
rect 267700 700000 267706 700052
rect 105446 699932 105452 699984
rect 105504 699972 105510 699984
rect 187970 699972 187976 699984
rect 105504 699944 187976 699972
rect 105504 699932 105510 699944
rect 187970 699932 187976 699944
rect 188028 699932 188034 699984
rect 173802 699864 173808 699916
rect 173860 699904 173866 699916
rect 235166 699904 235172 699916
rect 173860 699876 235172 699904
rect 173860 699864 173866 699876
rect 235166 699864 235172 699876
rect 235224 699864 235230 699916
rect 175918 699796 175924 699848
rect 175976 699836 175982 699848
rect 202782 699836 202788 699848
rect 175976 699808 202788 699836
rect 175976 699796 175982 699808
rect 202782 699796 202788 699808
rect 202840 699796 202846 699848
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 251450 699660 251456 699712
rect 251508 699700 251514 699712
rect 252462 699700 252468 699712
rect 251508 699672 252468 699700
rect 251508 699660 251514 699672
rect 252462 699660 252468 699672
rect 252520 699660 252526 699712
rect 381170 699660 381176 699712
rect 381228 699700 381234 699712
rect 382182 699700 382188 699712
rect 381228 699672 382188 699700
rect 381228 699660 381234 699672
rect 382182 699660 382188 699672
rect 382240 699660 382246 699712
rect 133598 696940 133604 696992
rect 133656 696980 133662 696992
rect 580166 696980 580172 696992
rect 133656 696952 580172 696980
rect 133656 696940 133662 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 410610 692792 410616 692844
rect 410668 692832 410674 692844
rect 463326 692832 463332 692844
rect 410668 692804 463332 692832
rect 410668 692792 410674 692804
rect 463326 692792 463332 692804
rect 463384 692792 463390 692844
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 188522 670732 188528 670744
rect 3568 670704 188528 670732
rect 3568 670692 3574 670704
rect 188522 670692 188528 670704
rect 188580 670692 188586 670744
rect 542354 670352 542360 670404
rect 542412 670392 542418 670404
rect 544749 670395 544807 670401
rect 544749 670392 544761 670395
rect 542412 670364 544761 670392
rect 542412 670352 542418 670364
rect 544749 670361 544761 670364
rect 544795 670361 544807 670395
rect 544749 670355 544807 670361
rect 542354 668380 542360 668432
rect 542412 668420 542418 668432
rect 544749 668423 544807 668429
rect 544749 668420 544761 668423
rect 542412 668392 544761 668420
rect 542412 668380 542418 668392
rect 544749 668389 544761 668392
rect 544795 668389 544807 668423
rect 544749 668383 544807 668389
rect 2866 657500 2872 657552
rect 2924 657540 2930 657552
rect 197814 657540 197820 657552
rect 2924 657512 197820 657540
rect 2924 657500 2930 657512
rect 197814 657500 197820 657512
rect 197872 657500 197878 657552
rect 429194 648320 429200 648372
rect 429252 648320 429258 648372
rect 429212 648100 429240 648320
rect 429194 648048 429200 648100
rect 429252 648048 429258 648100
rect 227714 647136 227720 647148
rect 226168 647108 227720 647136
rect 226168 646400 226196 647108
rect 227714 647096 227720 647108
rect 227772 647096 227778 647148
rect 226150 646348 226156 646400
rect 226208 646348 226214 646400
rect 226150 646048 226156 646060
rect 225708 646020 226156 646048
rect 4798 645872 4804 645924
rect 4856 645912 4862 645924
rect 32030 645912 32036 645924
rect 4856 645884 32036 645912
rect 4856 645872 4862 645884
rect 32030 645872 32036 645884
rect 32088 645872 32094 645924
rect 188433 645915 188491 645921
rect 188433 645881 188445 645915
rect 188479 645912 188491 645915
rect 188522 645912 188528 645924
rect 188479 645884 188528 645912
rect 188479 645881 188491 645884
rect 188433 645875 188491 645881
rect 188522 645872 188528 645884
rect 188580 645872 188586 645924
rect 196529 645915 196587 645921
rect 196529 645881 196541 645915
rect 196575 645912 196587 645915
rect 198182 645912 198188 645924
rect 196575 645884 198188 645912
rect 196575 645881 196587 645884
rect 196529 645875 196587 645881
rect 198182 645872 198188 645884
rect 198240 645872 198246 645924
rect 199841 645915 199899 645921
rect 199841 645881 199853 645915
rect 199887 645912 199899 645915
rect 225708 645912 225736 646020
rect 226150 646008 226156 646020
rect 226208 646008 226214 646060
rect 199887 645884 225736 645912
rect 199887 645881 199899 645884
rect 199841 645875 199899 645881
rect 475657 645847 475715 645853
rect 475657 645813 475669 645847
rect 475703 645844 475715 645847
rect 580350 645844 580356 645856
rect 475703 645816 580356 645844
rect 475703 645813 475715 645816
rect 475657 645807 475715 645813
rect 580350 645804 580356 645816
rect 580408 645804 580414 645856
rect 188062 645600 188068 645652
rect 188120 645600 188126 645652
rect 188338 645640 188344 645652
rect 188299 645612 188344 645640
rect 188338 645600 188344 645612
rect 188396 645600 188402 645652
rect 188430 645600 188436 645652
rect 188488 645600 188494 645652
rect 187970 645328 187976 645380
rect 188028 645368 188034 645380
rect 188080 645368 188108 645600
rect 188448 645380 188476 645600
rect 196342 645572 196348 645584
rect 196303 645544 196348 645572
rect 196342 645532 196348 645544
rect 196400 645532 196406 645584
rect 188028 645340 188108 645368
rect 188028 645328 188034 645340
rect 188430 645328 188436 645380
rect 188488 645328 188494 645380
rect 196529 645167 196587 645173
rect 196529 645133 196541 645167
rect 196575 645164 196587 645167
rect 197906 645164 197912 645176
rect 196575 645136 197912 645164
rect 196575 645133 196587 645136
rect 196529 645127 196587 645133
rect 197906 645124 197912 645136
rect 197964 645124 197970 645176
rect 471882 644852 471888 644904
rect 471940 644892 471946 644904
rect 475657 644895 475715 644901
rect 475657 644892 475669 644895
rect 471940 644864 475669 644892
rect 471940 644852 471946 644864
rect 475657 644861 475669 644864
rect 475703 644861 475715 644895
rect 475657 644855 475715 644861
rect 443641 644487 443699 644493
rect 443641 644453 443653 644487
rect 443687 644484 443699 644487
rect 459554 644484 459560 644496
rect 443687 644456 459560 644484
rect 443687 644453 443699 644456
rect 443641 644447 443699 644453
rect 459554 644444 459560 644456
rect 459612 644444 459618 644496
rect 429381 644011 429439 644017
rect 429381 643977 429393 644011
rect 429427 644008 429439 644011
rect 433061 644011 433119 644017
rect 433061 644008 433073 644011
rect 429427 643980 433073 644008
rect 429427 643977 429439 643980
rect 429381 643971 429439 643977
rect 433061 643977 433073 643980
rect 433107 643977 433119 644011
rect 433061 643971 433119 643977
rect 476945 643875 477003 643881
rect 476945 643872 476957 643875
rect 451246 643844 476957 643872
rect 426989 643535 427047 643541
rect 426989 643532 427001 643535
rect 412606 643504 427001 643532
rect 225785 643399 225843 643405
rect 225785 643396 225797 643399
rect 219406 643368 225797 643396
rect 124766 643288 124772 643340
rect 124824 643328 124830 643340
rect 128906 643328 128912 643340
rect 124824 643300 128912 643328
rect 124824 643288 124830 643300
rect 128906 643288 128912 643300
rect 128964 643288 128970 643340
rect 129274 643288 129280 643340
rect 129332 643328 129338 643340
rect 132770 643328 132776 643340
rect 129332 643300 132776 643328
rect 129332 643288 129338 643300
rect 132770 643288 132776 643300
rect 132828 643288 132834 643340
rect 133138 643288 133144 643340
rect 133196 643328 133202 643340
rect 136634 643328 136640 643340
rect 133196 643300 136640 643328
rect 133196 643288 133202 643300
rect 136634 643288 136640 643300
rect 136692 643288 136698 643340
rect 137002 643288 137008 643340
rect 137060 643328 137066 643340
rect 139765 643331 139823 643337
rect 139765 643328 139777 643331
rect 137060 643300 139777 643328
rect 137060 643288 137066 643300
rect 139765 643297 139777 643300
rect 139811 643297 139823 643331
rect 139765 643291 139823 643297
rect 140225 643331 140283 643337
rect 140225 643297 140237 643331
rect 140271 643328 140283 643331
rect 183189 643331 183247 643337
rect 183189 643328 183201 643331
rect 140271 643300 183201 643328
rect 140271 643297 140283 643300
rect 140225 643291 140283 643297
rect 183189 643297 183201 643300
rect 183235 643297 183247 643331
rect 183189 643291 183247 643297
rect 183557 643331 183615 643337
rect 183557 643297 183569 643331
rect 183603 643328 183615 643331
rect 219406 643328 219434 643368
rect 225785 643365 225797 643368
rect 225831 643365 225843 643399
rect 225785 643359 225843 643365
rect 183603 643300 219434 643328
rect 226429 643331 226487 643337
rect 183603 643297 183615 643300
rect 183557 643291 183615 643297
rect 226429 643297 226441 643331
rect 226475 643328 226487 643331
rect 233329 643331 233387 643337
rect 233329 643328 233341 643331
rect 226475 643300 233341 643328
rect 226475 643297 226487 643300
rect 226429 643291 226487 643297
rect 233329 643297 233341 643300
rect 233375 643297 233387 643331
rect 233329 643291 233387 643297
rect 233789 643331 233847 643337
rect 233789 643297 233801 643331
rect 233835 643328 233847 643331
rect 412606 643328 412634 643504
rect 426989 643501 427001 643504
rect 427035 643501 427047 643535
rect 426989 643495 427047 643501
rect 427449 643535 427507 643541
rect 427449 643501 427461 643535
rect 427495 643501 427507 643535
rect 427449 643495 427507 643501
rect 427464 643464 427492 643495
rect 427464 643436 429424 643464
rect 429396 643405 429424 643436
rect 429381 643399 429439 643405
rect 429381 643365 429393 643399
rect 429427 643365 429439 643399
rect 429381 643359 429439 643365
rect 233835 643300 412634 643328
rect 433061 643331 433119 643337
rect 233835 643297 233847 643300
rect 233789 643291 233847 643297
rect 433061 643297 433073 643331
rect 433107 643328 433119 643331
rect 451246 643328 451274 643844
rect 476945 643841 476957 643844
rect 476991 643841 477003 643875
rect 476945 643835 477003 643841
rect 433107 643300 451274 643328
rect 477497 643331 477555 643337
rect 433107 643297 433119 643300
rect 433061 643291 433119 643297
rect 477497 643297 477509 643331
rect 477543 643328 477555 643331
rect 579614 643328 579620 643340
rect 477543 643300 579620 643328
rect 477543 643297 477555 643300
rect 477497 643291 477555 643297
rect 579614 643288 579620 643300
rect 579672 643288 579678 643340
rect 443638 643192 443644 643204
rect 443599 643164 443644 643192
rect 443638 643152 443644 643164
rect 443696 643152 443702 643204
rect 196345 642379 196403 642385
rect 196345 642345 196357 642379
rect 196391 642376 196403 642379
rect 196894 642376 196900 642388
rect 196391 642348 196900 642376
rect 196391 642345 196403 642348
rect 196345 642339 196403 642345
rect 196894 642336 196900 642348
rect 196952 642336 196958 642388
rect 199562 640976 199568 641028
rect 199620 641016 199626 641028
rect 205560 641016 205588 641206
rect 214558 641016 214564 641028
rect 199620 640988 214564 641016
rect 199620 640976 199626 640988
rect 214558 640976 214564 640988
rect 214616 640976 214622 641028
rect 196986 640704 196992 640756
rect 197044 640744 197050 640756
rect 199841 640747 199899 640753
rect 199841 640744 199853 640747
rect 197044 640716 199853 640744
rect 197044 640704 197050 640716
rect 199841 640713 199853 640716
rect 199887 640713 199899 640747
rect 199841 640707 199899 640713
rect 90818 639888 90824 639940
rect 90876 639928 90882 639940
rect 96338 639928 96344 639940
rect 90876 639900 96344 639928
rect 90876 639888 90882 639900
rect 96338 639888 96344 639900
rect 96396 639888 96402 639940
rect 190273 639591 190331 639597
rect 190273 639557 190285 639591
rect 190319 639588 190331 639591
rect 191009 639591 191067 639597
rect 191009 639588 191021 639591
rect 190319 639560 191021 639588
rect 190319 639557 190331 639560
rect 190273 639551 190331 639557
rect 191009 639557 191021 639560
rect 191055 639557 191067 639591
rect 191009 639551 191067 639557
rect 191285 639591 191343 639597
rect 191285 639557 191297 639591
rect 191331 639588 191343 639591
rect 197446 639588 197452 639600
rect 191331 639560 197452 639588
rect 191331 639557 191343 639560
rect 191285 639551 191343 639557
rect 197446 639548 197452 639560
rect 197504 639548 197510 639600
rect 233878 639548 233884 639600
rect 233936 639588 233942 639600
rect 415302 639588 415308 639600
rect 233936 639560 415308 639588
rect 233936 639548 233942 639560
rect 415302 639548 415308 639560
rect 415360 639548 415366 639600
rect 189813 639523 189871 639529
rect 189813 639489 189825 639523
rect 189859 639520 189871 639523
rect 189997 639523 190055 639529
rect 189997 639520 190009 639523
rect 189859 639492 190009 639520
rect 189859 639489 189871 639492
rect 189813 639483 189871 639489
rect 189997 639489 190009 639492
rect 190043 639489 190055 639523
rect 189997 639483 190055 639489
rect 190365 639523 190423 639529
rect 190365 639489 190377 639523
rect 190411 639520 190423 639523
rect 190917 639523 190975 639529
rect 190917 639520 190929 639523
rect 190411 639492 190929 639520
rect 190411 639489 190423 639492
rect 190365 639483 190423 639489
rect 190917 639489 190929 639492
rect 190963 639489 190975 639523
rect 190917 639483 190975 639489
rect 191377 639523 191435 639529
rect 191377 639489 191389 639523
rect 191423 639520 191435 639523
rect 194686 639520 194692 639532
rect 191423 639492 194692 639520
rect 191423 639489 191435 639492
rect 191377 639483 191435 639489
rect 194686 639480 194692 639492
rect 194744 639480 194750 639532
rect 190273 639455 190331 639461
rect 190273 639421 190285 639455
rect 190319 639452 190331 639455
rect 191009 639455 191067 639461
rect 191009 639452 191021 639455
rect 190319 639424 191021 639452
rect 190319 639421 190331 639424
rect 190273 639415 190331 639421
rect 191009 639421 191021 639424
rect 191055 639421 191067 639455
rect 191009 639415 191067 639421
rect 191285 639455 191343 639461
rect 191285 639421 191297 639455
rect 191331 639452 191343 639455
rect 194594 639452 194600 639464
rect 191331 639424 194600 639452
rect 191331 639421 191343 639424
rect 191285 639415 191343 639421
rect 194594 639412 194600 639424
rect 194652 639412 194658 639464
rect 182910 639072 182916 639124
rect 182968 639112 182974 639124
rect 189905 639115 189963 639121
rect 189905 639112 189917 639115
rect 182968 639084 189917 639112
rect 182968 639072 182974 639084
rect 189905 639081 189917 639084
rect 189951 639081 189963 639115
rect 189905 639075 189963 639081
rect 196342 639072 196348 639124
rect 196400 639112 196406 639124
rect 197078 639112 197084 639124
rect 196400 639084 197084 639112
rect 196400 639072 196406 639084
rect 197078 639072 197084 639084
rect 197136 639072 197142 639124
rect 184014 639004 184020 639056
rect 184072 639044 184078 639056
rect 189997 639047 190055 639053
rect 189997 639044 190009 639047
rect 184072 639016 190009 639044
rect 184072 639004 184078 639016
rect 189997 639013 190009 639016
rect 190043 639013 190055 639047
rect 189997 639007 190055 639013
rect 182542 638936 182548 638988
rect 182600 638976 182606 638988
rect 189813 638979 189871 638985
rect 189813 638976 189825 638979
rect 182600 638948 189825 638976
rect 182600 638936 182606 638948
rect 189813 638945 189825 638948
rect 189859 638945 189871 638979
rect 189813 638939 189871 638945
rect 187970 638800 187976 638852
rect 188028 638800 188034 638852
rect 188430 638800 188436 638852
rect 188488 638800 188494 638852
rect 188982 638800 188988 638852
rect 189040 638800 189046 638852
rect 187988 638512 188016 638800
rect 188448 638512 188476 638800
rect 189000 638580 189028 638800
rect 188982 638528 188988 638580
rect 189040 638528 189046 638580
rect 187970 638460 187976 638512
rect 188028 638460 188034 638512
rect 188338 638500 188344 638512
rect 188299 638472 188344 638500
rect 188338 638460 188344 638472
rect 188396 638460 188402 638512
rect 188430 638460 188436 638512
rect 188488 638460 188494 638512
rect 196250 638392 196256 638444
rect 196308 638432 196314 638444
rect 196986 638432 196992 638444
rect 196308 638404 196992 638432
rect 196308 638392 196314 638404
rect 196986 638392 196992 638404
rect 197044 638392 197050 638444
rect 188433 638367 188491 638373
rect 188433 638333 188445 638367
rect 188479 638364 188491 638367
rect 188522 638364 188528 638376
rect 188479 638336 188528 638364
rect 188479 638333 188491 638336
rect 188433 638327 188491 638333
rect 188522 638324 188528 638336
rect 188580 638324 188586 638376
rect 214558 637848 214564 637900
rect 214616 637848 214622 637900
rect 218882 637848 218888 637900
rect 218940 637848 218946 637900
rect 214576 637628 214604 637848
rect 218900 637628 218928 637848
rect 214558 637576 214564 637628
rect 214616 637576 214622 637628
rect 218882 637576 218888 637628
rect 218940 637576 218946 637628
rect 217781 635987 217839 635993
rect 217781 635953 217793 635987
rect 217827 635984 217839 635987
rect 218882 635984 218888 635996
rect 217827 635956 218888 635984
rect 217827 635953 217839 635956
rect 217781 635947 217839 635953
rect 218882 635944 218888 635956
rect 218940 635944 218946 635996
rect 196250 635604 196256 635656
rect 196308 635604 196314 635656
rect 196342 635604 196348 635656
rect 196400 635644 196406 635656
rect 196400 635616 196445 635644
rect 196400 635604 196406 635616
rect 196158 635332 196164 635384
rect 196216 635372 196222 635384
rect 196268 635372 196296 635604
rect 196216 635344 196296 635372
rect 196216 635332 196222 635344
rect 196342 635168 196348 635180
rect 196303 635140 196348 635168
rect 196342 635128 196348 635140
rect 196400 635128 196406 635180
rect 90818 634924 90824 634976
rect 90876 634964 90882 634976
rect 96982 634964 96988 634976
rect 90876 634936 96988 634964
rect 90876 634924 90882 634936
rect 96982 634924 96988 634936
rect 97040 634924 97046 634976
rect 120258 634856 120264 634908
rect 120316 634896 120322 634908
rect 126790 634896 126796 634908
rect 120316 634868 126796 634896
rect 120316 634856 120322 634868
rect 126790 634856 126796 634868
rect 126848 634856 126854 634908
rect 189258 634856 189264 634908
rect 189316 634896 189322 634908
rect 191558 634896 191564 634908
rect 189316 634868 191564 634896
rect 189316 634856 189322 634868
rect 191558 634856 191564 634868
rect 191616 634856 191622 634908
rect 198458 634012 198464 634024
rect 198419 633984 198464 634012
rect 198458 633972 198464 633984
rect 198516 633972 198522 634024
rect 199562 634012 199568 634024
rect 199523 633984 199568 634012
rect 199562 633972 199568 633984
rect 199620 633972 199626 634024
rect 201957 633743 202015 633749
rect 201957 633709 201969 633743
rect 202003 633740 202015 633743
rect 202201 633740 202207 633752
rect 202003 633712 202207 633740
rect 202003 633709 202015 633712
rect 201957 633703 202015 633709
rect 202201 633700 202207 633712
rect 202259 633700 202265 633752
rect 3234 633360 3240 633412
rect 3292 633400 3298 633412
rect 58161 633403 58219 633409
rect 58161 633400 58173 633403
rect 3292 633372 58173 633400
rect 3292 633360 3298 633372
rect 58161 633369 58173 633372
rect 58207 633369 58219 633403
rect 58161 633363 58219 633369
rect 58621 633403 58679 633409
rect 58621 633369 58633 633403
rect 58667 633400 58679 633403
rect 97902 633400 97908 633412
rect 58667 633372 97908 633400
rect 58667 633369 58679 633372
rect 58621 633363 58679 633369
rect 97902 633360 97908 633372
rect 97960 633360 97966 633412
rect 214101 632791 214159 632797
rect 214101 632757 214113 632791
rect 214147 632788 214159 632791
rect 214558 632788 214564 632800
rect 214147 632760 214564 632788
rect 214147 632757 214159 632760
rect 214101 632751 214159 632757
rect 214558 632748 214564 632760
rect 214616 632748 214622 632800
rect 99742 632680 99748 632732
rect 99800 632720 99806 632732
rect 117777 632723 117835 632729
rect 117777 632720 117789 632723
rect 99800 632692 117789 632720
rect 99800 632680 99806 632692
rect 117777 632689 117789 632692
rect 117823 632689 117835 632723
rect 117777 632683 117835 632689
rect 118421 632723 118479 632729
rect 118421 632689 118433 632723
rect 118467 632720 118479 632723
rect 126882 632720 126888 632732
rect 118467 632692 126888 632720
rect 118467 632689 118479 632692
rect 118421 632683 118479 632689
rect 126882 632680 126888 632692
rect 126940 632680 126946 632732
rect 198458 632516 198464 632528
rect 198419 632488 198464 632516
rect 198458 632476 198464 632488
rect 198516 632476 198522 632528
rect 199562 632516 199568 632528
rect 199523 632488 199568 632516
rect 199562 632476 199568 632488
rect 199620 632476 199626 632528
rect 189810 632408 189816 632460
rect 189868 632448 189874 632460
rect 191558 632448 191564 632460
rect 189868 632420 191564 632448
rect 189868 632408 189874 632420
rect 191558 632408 191564 632420
rect 191616 632408 191622 632460
rect 201954 632244 201960 632256
rect 201915 632216 201960 632244
rect 201954 632204 201960 632216
rect 202012 632204 202018 632256
rect 436738 631796 436744 631848
rect 436796 631836 436802 631848
rect 436796 631808 438900 631836
rect 436796 631796 436802 631808
rect 212445 631771 212503 631777
rect 212445 631737 212457 631771
rect 212491 631768 212503 631771
rect 215386 631768 215392 631780
rect 212491 631740 215392 631768
rect 212491 631737 212503 631740
rect 212445 631731 212503 631737
rect 215386 631728 215392 631740
rect 215444 631728 215450 631780
rect 438872 631768 438900 631808
rect 441525 631771 441583 631777
rect 441525 631768 441537 631771
rect 438872 631740 441537 631768
rect 441525 631737 441537 631740
rect 441571 631737 441583 631771
rect 441525 631731 441583 631737
rect 128262 631388 128268 631440
rect 128320 631428 128326 631440
rect 128906 631428 128912 631440
rect 128320 631400 128912 631428
rect 128320 631388 128326 631400
rect 128906 631388 128912 631400
rect 128964 631388 128970 631440
rect 129274 631388 129280 631440
rect 129332 631428 129338 631440
rect 132770 631428 132776 631440
rect 129332 631400 132776 631428
rect 129332 631388 129338 631400
rect 132770 631388 132776 631400
rect 132828 631388 132834 631440
rect 133138 631388 133144 631440
rect 133196 631428 133202 631440
rect 136634 631428 136640 631440
rect 133196 631400 136640 631428
rect 133196 631388 133202 631400
rect 136634 631388 136640 631400
rect 136692 631388 136698 631440
rect 137002 631388 137008 631440
rect 137060 631428 137066 631440
rect 139765 631431 139823 631437
rect 139765 631428 139777 631431
rect 137060 631400 139777 631428
rect 137060 631388 137066 631400
rect 139765 631397 139777 631400
rect 139811 631397 139823 631431
rect 139765 631391 139823 631397
rect 140225 631431 140283 631437
rect 140225 631397 140237 631431
rect 140271 631428 140283 631431
rect 191558 631428 191564 631440
rect 140271 631400 191564 631428
rect 140271 631397 140283 631400
rect 140225 631391 140283 631397
rect 191558 631388 191564 631400
rect 191616 631388 191622 631440
rect 196069 631431 196127 631437
rect 196069 631428 196081 631431
rect 194152 631400 196081 631428
rect 192938 631116 192944 631168
rect 192996 631156 193002 631168
rect 194152 631156 194180 631400
rect 196069 631397 196081 631400
rect 196115 631397 196127 631431
rect 196069 631391 196127 631397
rect 196345 631431 196403 631437
rect 196345 631397 196357 631431
rect 196391 631428 196403 631431
rect 212445 631431 212503 631437
rect 212445 631428 212457 631431
rect 196391 631400 212457 631428
rect 196391 631397 196403 631400
rect 196345 631391 196403 631397
rect 212445 631397 212457 631400
rect 212491 631397 212503 631431
rect 212445 631391 212503 631397
rect 579798 631360 579804 631372
rect 509206 631332 579804 631360
rect 506658 631184 506664 631236
rect 506716 631224 506722 631236
rect 509206 631224 509234 631332
rect 579798 631320 579804 631332
rect 579856 631320 579862 631372
rect 506716 631196 509234 631224
rect 506716 631184 506722 631196
rect 192996 631128 194180 631156
rect 192996 631116 193002 631128
rect 441525 630819 441583 630825
rect 441525 630785 441537 630819
rect 441571 630816 441583 630819
rect 477497 630819 477555 630825
rect 441571 630788 460244 630816
rect 441571 630785 441583 630788
rect 441525 630779 441583 630785
rect 221090 630640 221096 630692
rect 221148 630680 221154 630692
rect 224865 630683 224923 630689
rect 224865 630680 224877 630683
rect 221148 630652 224877 630680
rect 221148 630640 221154 630652
rect 224865 630649 224877 630652
rect 224911 630649 224923 630683
rect 224865 630643 224923 630649
rect 225141 630683 225199 630689
rect 225141 630649 225153 630683
rect 225187 630680 225199 630683
rect 228545 630683 228603 630689
rect 228545 630680 228557 630683
rect 225187 630652 228557 630680
rect 225187 630649 225199 630652
rect 225141 630643 225199 630649
rect 228545 630649 228557 630652
rect 228591 630649 228603 630683
rect 228545 630643 228603 630649
rect 228913 630683 228971 630689
rect 228913 630649 228925 630683
rect 228959 630680 228971 630683
rect 405645 630683 405703 630689
rect 405645 630680 405657 630683
rect 228959 630652 405657 630680
rect 228959 630649 228971 630652
rect 228913 630643 228971 630649
rect 405645 630649 405657 630652
rect 405691 630649 405703 630683
rect 405645 630643 405703 630649
rect 460216 630612 460244 630788
rect 477497 630785 477509 630819
rect 477543 630816 477555 630819
rect 496078 630816 496084 630828
rect 477543 630788 496084 630816
rect 477543 630785 477555 630788
rect 477497 630779 477555 630785
rect 496078 630776 496084 630788
rect 496136 630776 496142 630828
rect 462041 630683 462099 630689
rect 462041 630680 462053 630683
rect 460952 630652 462053 630680
rect 460952 630612 460980 630652
rect 462041 630649 462053 630652
rect 462087 630649 462099 630683
rect 462041 630643 462099 630649
rect 462409 630683 462467 630689
rect 462409 630649 462421 630683
rect 462455 630680 462467 630683
rect 477037 630683 477095 630689
rect 477037 630680 477049 630683
rect 462455 630652 477049 630680
rect 462455 630649 462467 630652
rect 462409 630643 462467 630649
rect 477037 630649 477049 630652
rect 477083 630649 477095 630683
rect 477037 630643 477095 630649
rect 460216 630584 460980 630612
rect 214101 629323 214159 629329
rect 214101 629289 214113 629323
rect 214147 629289 214159 629323
rect 214101 629283 214159 629289
rect 214116 629125 214144 629283
rect 214101 629119 214159 629125
rect 214101 629085 214113 629119
rect 214147 629085 214159 629119
rect 214101 629079 214159 629085
rect 217781 629119 217839 629125
rect 217781 629085 217793 629119
rect 217827 629116 217839 629119
rect 218882 629116 218888 629128
rect 217827 629088 218888 629116
rect 217827 629085 217839 629088
rect 217781 629079 217839 629085
rect 218882 629076 218888 629088
rect 218940 629076 218946 629128
rect 405737 628983 405795 628989
rect 405737 628949 405749 628983
rect 405783 628980 405795 628983
rect 414658 628980 414664 628992
rect 405783 628952 414664 628980
rect 405783 628949 405795 628952
rect 405737 628943 405795 628949
rect 414658 628940 414664 628952
rect 414716 628940 414722 628992
rect 198458 628300 198464 628312
rect 197832 628272 198464 628300
rect 197832 627972 197860 628272
rect 198458 628260 198464 628272
rect 198516 628260 198522 628312
rect 199562 628260 199568 628312
rect 199620 628260 199626 628312
rect 199580 627972 199608 628260
rect 201954 628192 201960 628244
rect 202012 628192 202018 628244
rect 210234 628192 210240 628244
rect 210292 628232 210298 628244
rect 214101 628235 214159 628241
rect 210292 628204 211016 628232
rect 210292 628192 210298 628204
rect 197354 627960 197360 627972
rect 197315 627932 197360 627960
rect 197354 627920 197360 627932
rect 197412 627920 197418 627972
rect 197814 627920 197820 627972
rect 197872 627920 197878 627972
rect 199562 627920 199568 627972
rect 199620 627920 199626 627972
rect 201972 627904 202000 628192
rect 210988 628040 211016 628204
rect 214101 628201 214113 628235
rect 214147 628232 214159 628235
rect 214558 628232 214564 628244
rect 214147 628204 214564 628232
rect 214147 628201 214159 628204
rect 214101 628195 214159 628201
rect 214558 628192 214564 628204
rect 214616 628192 214622 628244
rect 210970 627988 210976 628040
rect 211028 627988 211034 628040
rect 201954 627852 201960 627904
rect 202012 627852 202018 627904
rect 218882 627756 218888 627768
rect 218843 627728 218888 627756
rect 218882 627716 218888 627728
rect 218940 627716 218946 627768
rect 214558 626764 214564 626816
rect 214616 626764 214622 626816
rect 214576 626612 214604 626764
rect 214558 626560 214564 626612
rect 214616 626560 214622 626612
rect 187970 624656 187976 624708
rect 188028 624656 188034 624708
rect 188338 624656 188344 624708
rect 188396 624656 188402 624708
rect 188430 624656 188436 624708
rect 188488 624656 188494 624708
rect 188522 624656 188528 624708
rect 188580 624656 188586 624708
rect 188982 624656 188988 624708
rect 189040 624656 189046 624708
rect 187988 624368 188016 624656
rect 188356 624368 188384 624656
rect 188448 624368 188476 624656
rect 188540 624368 188568 624656
rect 189000 624368 189028 624656
rect 187970 624316 187976 624368
rect 188028 624316 188034 624368
rect 188338 624316 188344 624368
rect 188396 624316 188402 624368
rect 188430 624316 188436 624368
rect 188488 624316 188494 624368
rect 188522 624316 188528 624368
rect 188580 624316 188586 624368
rect 188982 624316 188988 624368
rect 189040 624316 189046 624368
rect 542354 623024 542360 623076
rect 542412 623064 542418 623076
rect 545761 623067 545819 623073
rect 545761 623064 545773 623067
rect 542412 623036 545773 623064
rect 542412 623024 542418 623036
rect 545761 623033 545773 623036
rect 545807 623033 545819 623067
rect 545761 623027 545819 623033
rect 128262 621868 128268 621920
rect 128320 621868 128326 621920
rect 128280 621376 128308 621868
rect 128262 621324 128268 621376
rect 128320 621324 128326 621376
rect 3602 620984 3608 621036
rect 3660 621024 3666 621036
rect 31754 621024 31760 621036
rect 3660 620996 31760 621024
rect 3660 620984 3666 620996
rect 31754 620984 31760 620996
rect 31812 620984 31818 621036
rect 218882 620004 218888 620016
rect 218843 619976 218888 620004
rect 218882 619964 218888 619976
rect 218940 619964 218946 620016
rect 542446 619828 542452 619880
rect 542504 619868 542510 619880
rect 545761 619871 545819 619877
rect 545761 619868 545773 619871
rect 542504 619840 545773 619868
rect 542504 619828 542510 619840
rect 545761 619837 545773 619840
rect 545807 619837 545819 619871
rect 545761 619831 545819 619837
rect 3510 619624 3516 619676
rect 3568 619664 3574 619676
rect 31754 619664 31760 619676
rect 3568 619636 31760 619664
rect 3568 619624 3574 619636
rect 31754 619624 31760 619636
rect 31812 619624 31818 619676
rect 382182 619624 382188 619676
rect 382240 619664 382246 619676
rect 382240 619636 452778 619664
rect 382240 619624 382246 619636
rect 142126 619024 151814 619052
rect 138477 618987 138535 618993
rect 138477 618984 138489 618987
rect 132466 618956 138489 618984
rect 3418 618536 3424 618588
rect 3476 618576 3482 618588
rect 79226 618576 79232 618588
rect 3476 618548 26234 618576
rect 3476 618536 3482 618548
rect 26206 618304 26234 618548
rect 45526 618548 79232 618576
rect 45526 618304 45554 618548
rect 79226 618536 79232 618548
rect 79284 618536 79290 618588
rect 79778 618536 79784 618588
rect 79836 618576 79842 618588
rect 132466 618576 132494 618956
rect 138477 618953 138489 618956
rect 138523 618953 138535 618987
rect 138477 618947 138535 618953
rect 137094 618916 137100 618928
rect 137055 618888 137100 618916
rect 137094 618876 137100 618888
rect 137152 618876 137158 618928
rect 79836 618548 132494 618576
rect 139029 618579 139087 618585
rect 79836 618536 79842 618548
rect 139029 618545 139041 618579
rect 139075 618576 139087 618579
rect 142126 618576 142154 619024
rect 139075 618548 142154 618576
rect 151786 618576 151814 619024
rect 199562 618576 199568 618588
rect 151786 618548 199568 618576
rect 139075 618545 139087 618548
rect 139029 618539 139087 618545
rect 199562 618536 199568 618548
rect 199620 618536 199626 618588
rect 137094 618304 137100 618316
rect 26206 618276 45554 618304
rect 137055 618276 137100 618304
rect 137094 618264 137100 618276
rect 137152 618264 137158 618316
rect 124122 617992 124128 618044
rect 124180 618032 124186 618044
rect 131482 618032 131488 618044
rect 124180 618004 131488 618032
rect 124180 617992 124186 618004
rect 131482 617992 131488 618004
rect 131540 617992 131546 618044
rect 132034 617040 132040 617092
rect 132092 617080 132098 617092
rect 137281 617083 137339 617089
rect 137281 617080 137293 617083
rect 132092 617052 137293 617080
rect 132092 617040 132098 617052
rect 137281 617049 137293 617052
rect 137327 617049 137339 617083
rect 137281 617043 137339 617049
rect 137649 617083 137707 617089
rect 137649 617049 137661 617083
rect 137695 617080 137707 617083
rect 138477 617083 138535 617089
rect 138477 617080 138489 617083
rect 137695 617052 138489 617080
rect 137695 617049 137707 617052
rect 137649 617043 137707 617049
rect 138477 617049 138489 617052
rect 138523 617049 138535 617083
rect 138477 617043 138535 617049
rect 139029 617083 139087 617089
rect 139029 617049 139041 617083
rect 139075 617080 139087 617083
rect 146757 617083 146815 617089
rect 146757 617080 146769 617083
rect 139075 617052 146769 617080
rect 139075 617049 139087 617052
rect 139029 617043 139087 617049
rect 146757 617049 146769 617052
rect 146803 617049 146815 617083
rect 146757 617043 146815 617049
rect 147493 617083 147551 617089
rect 147493 617049 147505 617083
rect 147539 617080 147551 617083
rect 580166 617080 580172 617092
rect 147539 617052 580172 617080
rect 147539 617049 147551 617052
rect 147493 617043 147551 617049
rect 580166 617040 580172 617052
rect 580224 617040 580230 617092
rect 160094 607112 160100 607164
rect 160152 607152 160158 607164
rect 160922 607152 160928 607164
rect 160152 607124 160928 607152
rect 160152 607112 160158 607124
rect 160922 607112 160928 607124
rect 160980 607112 160986 607164
rect 124122 601944 124128 601996
rect 124180 601944 124186 601996
rect 124766 601944 124772 601996
rect 124824 601944 124830 601996
rect 128262 601944 128268 601996
rect 128320 601944 128326 601996
rect 133598 601944 133604 601996
rect 133656 601944 133662 601996
rect 124140 601588 124168 601944
rect 124784 601588 124812 601944
rect 128280 601588 128308 601944
rect 133616 601588 133644 601944
rect 124122 601536 124128 601588
rect 124180 601536 124186 601588
rect 124766 601536 124772 601588
rect 124824 601536 124830 601588
rect 128262 601536 128268 601588
rect 128320 601536 128326 601588
rect 133598 601536 133604 601588
rect 133656 601536 133662 601588
rect 159542 591268 159548 591320
rect 159600 591308 159606 591320
rect 580166 591308 580172 591320
rect 159600 591280 580172 591308
rect 159600 591268 159606 591280
rect 580166 591268 580172 591280
rect 580224 591268 580230 591320
rect 3510 578212 3516 578264
rect 3568 578252 3574 578264
rect 31846 578252 31852 578264
rect 3568 578224 31852 578252
rect 3568 578212 3574 578224
rect 31846 578212 31852 578224
rect 31904 578212 31910 578264
rect 98638 577980 98644 577992
rect 98599 577952 98644 577980
rect 98638 577940 98644 577952
rect 98696 577940 98702 577992
rect 98638 577572 98644 577584
rect 98599 577544 98644 577572
rect 98638 577532 98644 577544
rect 98696 577532 98702 577584
rect 139486 577464 139492 577516
rect 139544 577504 139550 577516
rect 145561 577507 145619 577513
rect 145561 577504 145573 577507
rect 139544 577476 145573 577504
rect 139544 577464 139550 577476
rect 145561 577473 145573 577476
rect 145607 577473 145619 577507
rect 145561 577467 145619 577473
rect 146297 577507 146355 577513
rect 146297 577473 146309 577507
rect 146343 577504 146355 577507
rect 152001 577507 152059 577513
rect 152001 577504 152013 577507
rect 146343 577476 152013 577504
rect 146343 577473 146355 577476
rect 146297 577467 146355 577473
rect 152001 577473 152013 577476
rect 152047 577473 152059 577507
rect 152001 577467 152059 577473
rect 152737 577507 152795 577513
rect 152737 577473 152749 577507
rect 152783 577504 152795 577507
rect 158717 577507 158775 577513
rect 158717 577504 158729 577507
rect 152783 577476 158729 577504
rect 152783 577473 152795 577476
rect 152737 577467 152795 577473
rect 158717 577473 158729 577476
rect 158763 577473 158775 577507
rect 158717 577467 158775 577473
rect 159453 577507 159511 577513
rect 159453 577473 159465 577507
rect 159499 577504 159511 577507
rect 579982 577504 579988 577516
rect 159499 577476 579988 577504
rect 159499 577473 159511 577476
rect 159453 577467 159511 577473
rect 579982 577464 579988 577476
rect 580040 577464 580046 577516
rect 410334 569916 410340 569968
rect 410392 569956 410398 569968
rect 410610 569956 410616 569968
rect 410392 569928 410616 569956
rect 410392 569916 410398 569928
rect 410610 569916 410616 569928
rect 410668 569956 410674 569968
rect 579614 569956 579620 569968
rect 410668 569928 579620 569956
rect 410668 569916 410674 569928
rect 579614 569916 579620 569928
rect 579672 569916 579678 569968
rect 404262 566856 404268 566908
rect 404320 566856 404326 566908
rect 404280 566488 404308 566856
rect 427814 566488 427820 566500
rect 404280 566460 427820 566488
rect 427814 566448 427820 566460
rect 427872 566448 427878 566500
rect 92382 558900 92388 558952
rect 92440 558940 92446 558952
rect 391842 558940 391848 558952
rect 92440 558912 391848 558940
rect 92440 558900 92446 558912
rect 391842 558900 391848 558912
rect 391900 558900 391906 558952
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 211798 553432 211804 553444
rect 3384 553404 211804 553432
rect 3384 553392 3390 553404
rect 211798 553392 211804 553404
rect 211856 553392 211862 553444
rect 99282 542376 99288 542428
rect 99340 542416 99346 542428
rect 391382 542416 391388 542428
rect 99340 542388 391388 542416
rect 99340 542376 99346 542388
rect 391382 542376 391388 542388
rect 391440 542416 391446 542428
rect 391750 542416 391756 542428
rect 391440 542388 391756 542416
rect 391440 542376 391446 542388
rect 391750 542376 391756 542388
rect 391808 542376 391814 542428
rect 3326 540880 3332 540932
rect 3384 540920 3390 540932
rect 31754 540920 31760 540932
rect 3384 540892 31760 540920
rect 3384 540880 3390 540892
rect 31754 540880 31760 540892
rect 31812 540880 31818 540932
rect 111702 536800 111708 536852
rect 111760 536840 111766 536852
rect 580166 536840 580172 536852
rect 111760 536812 580172 536840
rect 111760 536800 111766 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 417694 534012 417700 534064
rect 417752 534052 417758 534064
rect 580350 534052 580356 534064
rect 417752 534024 580356 534052
rect 417752 534012 417758 534024
rect 580350 534012 580356 534024
rect 580408 534012 580414 534064
rect 401594 533944 401600 533996
rect 401652 533984 401658 533996
rect 402054 533984 402060 533996
rect 401652 533956 402060 533984
rect 401652 533944 401658 533956
rect 402054 533944 402060 533956
rect 402112 533984 402118 533996
rect 542354 533984 542360 533996
rect 402112 533956 542360 533984
rect 402112 533944 402118 533956
rect 542354 533944 542360 533956
rect 542412 533944 542418 533996
rect 143442 533400 143448 533452
rect 143500 533440 143506 533452
rect 401594 533440 401600 533452
rect 143500 533412 401600 533440
rect 143500 533400 143506 533412
rect 401594 533400 401600 533412
rect 401652 533400 401658 533452
rect 115842 533332 115848 533384
rect 115900 533372 115906 533384
rect 417694 533372 417700 533384
rect 115900 533344 417700 533372
rect 115900 533332 115906 533344
rect 417694 533332 417700 533344
rect 417752 533332 417758 533384
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 223574 527184 223580 527196
rect 3384 527156 223580 527184
rect 3384 527144 3390 527156
rect 223574 527144 223580 527156
rect 223632 527144 223638 527196
rect 114462 524424 114468 524476
rect 114520 524464 114526 524476
rect 580166 524464 580172 524476
rect 114520 524436 580172 524464
rect 114520 524424 114526 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 515380 3332 515432
rect 3384 515420 3390 515432
rect 197354 515420 197360 515432
rect 3384 515392 197360 515420
rect 3384 515380 3390 515392
rect 197354 515380 197360 515392
rect 197412 515380 197418 515432
rect 197354 514768 197360 514820
rect 197412 514808 197418 514820
rect 197998 514808 198004 514820
rect 197412 514780 198004 514808
rect 197412 514768 197418 514780
rect 197998 514768 198004 514780
rect 198056 514768 198062 514820
rect 108942 510620 108948 510672
rect 109000 510660 109006 510672
rect 580166 510660 580172 510672
rect 109000 510632 580172 510660
rect 109000 510620 109006 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 2866 500964 2872 501016
rect 2924 501004 2930 501016
rect 218698 501004 218704 501016
rect 2924 500976 218704 501004
rect 2924 500964 2930 500976
rect 218698 500964 218704 500976
rect 218756 500964 218762 501016
rect 104802 484372 104808 484424
rect 104860 484412 104866 484424
rect 579982 484412 579988 484424
rect 104860 484384 579988 484412
rect 104860 484372 104866 484384
rect 579982 484372 579988 484384
rect 580040 484372 580046 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 230474 474756 230480 474768
rect 3108 474728 230480 474756
rect 3108 474716 3114 474728
rect 230474 474716 230480 474728
rect 230532 474716 230538 474768
rect 106182 470568 106188 470620
rect 106240 470608 106246 470620
rect 580166 470608 580172 470620
rect 106240 470580 580172 470608
rect 106240 470568 106246 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 200758 462380 200764 462392
rect 3384 462352 200764 462380
rect 3384 462340 3390 462352
rect 200758 462340 200764 462352
rect 200816 462340 200822 462392
rect 100754 457444 100760 457496
rect 100812 457484 100818 457496
rect 579614 457484 579620 457496
rect 100812 457456 579620 457484
rect 100812 457444 100818 457456
rect 579614 457444 579620 457456
rect 579672 457444 579678 457496
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 226978 448576 226984 448588
rect 3384 448548 226984 448576
rect 3384 448536 3390 448548
rect 226978 448536 226984 448548
rect 227036 448536 227042 448588
rect 96522 430584 96528 430636
rect 96580 430624 96586 430636
rect 579890 430624 579896 430636
rect 96580 430596 579896 430624
rect 96580 430584 96586 430596
rect 579890 430584 579896 430596
rect 579948 430584 579954 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 237374 422328 237380 422340
rect 3568 422300 237380 422328
rect 3568 422288 3574 422300
rect 237374 422288 237380 422300
rect 237432 422288 237438 422340
rect 391750 419432 391756 419484
rect 391808 419472 391814 419484
rect 580166 419472 580172 419484
rect 391808 419444 580172 419472
rect 391808 419432 391814 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 221458 409884 221464 409896
rect 2924 409856 221464 409884
rect 2924 409844 2930 409856
rect 221458 409844 221464 409856
rect 221516 409844 221522 409896
rect 95142 404336 95148 404388
rect 95200 404376 95206 404388
rect 580166 404376 580172 404388
rect 95200 404348 580172 404376
rect 95200 404336 95206 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 233878 397508 233884 397520
rect 3568 397480 233884 397508
rect 3568 397468 3574 397480
rect 233878 397468 233884 397480
rect 233936 397468 233942 397520
rect 89622 378156 89628 378208
rect 89680 378196 89686 378208
rect 580166 378196 580172 378208
rect 89680 378168 580172 378196
rect 89680 378156 89686 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3510 371220 3516 371272
rect 3568 371260 3574 371272
rect 245654 371260 245660 371272
rect 3568 371232 245660 371260
rect 3568 371220 3574 371232
rect 245654 371220 245660 371232
rect 245712 371220 245718 371272
rect 391842 365644 391848 365696
rect 391900 365684 391906 365696
rect 580166 365684 580172 365696
rect 391900 365656 580172 365684
rect 391900 365644 391906 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 88242 351908 88248 351960
rect 88300 351948 88306 351960
rect 580166 351948 580172 351960
rect 88300 351920 580172 351948
rect 88300 351908 88306 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 82538 324300 82544 324352
rect 82596 324340 82602 324352
rect 580166 324340 580172 324352
rect 82596 324312 580172 324340
rect 82596 324300 82602 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 252738 318832 252744 318844
rect 3384 318804 252744 318832
rect 3384 318792 3390 318804
rect 252738 318792 252744 318804
rect 252796 318792 252802 318844
rect 171042 314236 171048 314288
rect 171100 314276 171106 314288
rect 180886 314276 180892 314288
rect 171100 314248 180892 314276
rect 171100 314236 171106 314248
rect 180886 314236 180892 314248
rect 180944 314236 180950 314288
rect 98638 314168 98644 314220
rect 98696 314208 98702 314220
rect 192570 314208 192576 314220
rect 98696 314180 192576 314208
rect 98696 314168 98702 314180
rect 192570 314168 192576 314180
rect 192628 314168 192634 314220
rect 197998 314168 198004 314220
rect 198056 314208 198062 314220
rect 228726 314208 228732 314220
rect 198056 314180 228732 314208
rect 198056 314168 198062 314180
rect 228726 314168 228732 314180
rect 228784 314168 228790 314220
rect 166810 314100 166816 314152
rect 166868 314140 166874 314152
rect 299474 314140 299480 314152
rect 166868 314112 299480 314140
rect 166868 314100 166874 314112
rect 299474 314100 299480 314112
rect 299532 314100 299538 314152
rect 3418 314032 3424 314084
rect 3476 314072 3482 314084
rect 216674 314072 216680 314084
rect 3476 314044 216680 314072
rect 3476 314032 3482 314044
rect 216674 314032 216680 314044
rect 216732 314032 216738 314084
rect 135070 313964 135076 314016
rect 135128 314004 135134 314016
rect 443638 314004 443644 314016
rect 135128 313976 443644 314004
rect 135128 313964 135134 313976
rect 443638 313964 443644 313976
rect 443696 313964 443702 314016
rect 130654 313896 130660 313948
rect 130712 313936 130718 313948
rect 580258 313936 580264 313948
rect 130712 313908 580264 313936
rect 130712 313896 130718 313908
rect 580258 313896 580264 313908
rect 580316 313896 580322 313948
rect 188338 313216 188344 313268
rect 188396 313256 188402 313268
rect 190454 313256 190460 313268
rect 188396 313228 190460 313256
rect 188396 313216 188402 313228
rect 190454 313216 190460 313228
rect 190512 313216 190518 313268
rect 196342 313216 196348 313268
rect 196400 313256 196406 313268
rect 200114 313256 200120 313268
rect 196400 313228 200120 313256
rect 196400 313216 196406 313228
rect 200114 313216 200120 313228
rect 200172 313216 200178 313268
rect 204898 313216 204904 313268
rect 204956 313256 204962 313268
rect 211890 313256 211896 313268
rect 204956 313228 211896 313256
rect 204956 313216 204962 313228
rect 211890 313216 211896 313228
rect 211948 313216 211954 313268
rect 218882 313216 218888 313268
rect 218940 313256 218946 313268
rect 221550 313256 221556 313268
rect 218940 313228 221556 313256
rect 218940 313216 218946 313228
rect 221550 313216 221556 313228
rect 221608 313216 221614 313268
rect 233878 313216 233884 313268
rect 233936 313256 233942 313268
rect 240778 313256 240784 313268
rect 233936 313228 240784 313256
rect 233936 313216 233942 313228
rect 240778 313216 240784 313228
rect 240836 313216 240842 313268
rect 154390 313148 154396 313200
rect 154448 313188 154454 313200
rect 154448 313160 161474 313188
rect 154448 313148 154454 313160
rect 142706 313080 142712 313132
rect 142764 313120 142770 313132
rect 143442 313120 143448 313132
rect 142764 313092 143448 313120
rect 142764 313080 142770 313092
rect 143442 313080 143448 313092
rect 143500 313080 143506 313132
rect 147490 313080 147496 313132
rect 147548 313120 147554 313132
rect 148318 313120 148324 313132
rect 147548 313092 148324 313120
rect 147548 313080 147554 313092
rect 148318 313080 148324 313092
rect 148376 313080 148382 313132
rect 149882 313080 149888 313132
rect 149940 313120 149946 313132
rect 150342 313120 150348 313132
rect 149940 313092 150348 313120
rect 149940 313080 149946 313092
rect 150342 313080 150348 313092
rect 150400 313080 150406 313132
rect 152274 313080 152280 313132
rect 152332 313120 152338 313132
rect 153102 313120 153108 313132
rect 152332 313092 153108 313120
rect 152332 313080 152338 313092
rect 153102 313080 153108 313092
rect 153160 313080 153166 313132
rect 159542 313080 159548 313132
rect 159600 313120 159606 313132
rect 160002 313120 160008 313132
rect 159600 313092 160008 313120
rect 159600 313080 159606 313092
rect 160002 313080 160008 313092
rect 160060 313080 160066 313132
rect 161446 313120 161474 313160
rect 161934 313148 161940 313200
rect 161992 313188 161998 313200
rect 162762 313188 162768 313200
rect 161992 313160 162768 313188
rect 161992 313148 161998 313160
rect 162762 313148 162768 313160
rect 162820 313148 162826 313200
rect 169202 313148 169208 313200
rect 169260 313188 169266 313200
rect 169662 313188 169668 313200
rect 169260 313160 169668 313188
rect 169260 313148 169266 313160
rect 169662 313148 169668 313160
rect 169720 313148 169726 313200
rect 171594 313148 171600 313200
rect 171652 313188 171658 313200
rect 172422 313188 172428 313200
rect 171652 313160 172428 313188
rect 171652 313148 171658 313160
rect 172422 313148 172428 313160
rect 172480 313148 172486 313200
rect 178770 313148 178776 313200
rect 178828 313188 178834 313200
rect 188430 313188 188436 313200
rect 178828 313160 188436 313188
rect 178828 313148 178834 313160
rect 188430 313148 188436 313160
rect 188488 313148 188494 313200
rect 195609 313191 195667 313197
rect 195609 313157 195621 313191
rect 195655 313188 195667 313191
rect 197446 313188 197452 313200
rect 195655 313160 197452 313188
rect 195655 313157 195667 313160
rect 195609 313151 195667 313157
rect 197446 313148 197452 313160
rect 197504 313148 197510 313200
rect 197814 313148 197820 313200
rect 197872 313188 197878 313200
rect 204622 313188 204628 313200
rect 197872 313160 204628 313188
rect 197872 313148 197878 313160
rect 204622 313148 204628 313160
rect 204680 313148 204686 313200
rect 218698 313148 218704 313200
rect 218756 313188 218762 313200
rect 226334 313188 226340 313200
rect 218756 313160 226340 313188
rect 218756 313148 218762 313160
rect 226334 313148 226340 313160
rect 226392 313148 226398 313200
rect 226978 313148 226984 313200
rect 227036 313188 227042 313200
rect 233510 313188 233516 313200
rect 227036 313160 233516 313188
rect 227036 313148 227042 313160
rect 233510 313148 233516 313160
rect 233568 313148 233574 313200
rect 185394 313120 185400 313132
rect 161446 313092 185400 313120
rect 185394 313080 185400 313092
rect 185452 313080 185458 313132
rect 188522 313080 188528 313132
rect 188580 313120 188586 313132
rect 207014 313120 207020 313132
rect 188580 313092 207020 313120
rect 188580 313080 188586 313092
rect 207014 313080 207020 313092
rect 207072 313080 207078 313132
rect 211798 313080 211804 313132
rect 211856 313120 211862 313132
rect 219066 313120 219072 313132
rect 211856 313092 219072 313120
rect 211856 313080 211862 313092
rect 219066 313080 219072 313092
rect 219124 313080 219130 313132
rect 221458 313080 221464 313132
rect 221516 313120 221522 313132
rect 243170 313120 243176 313132
rect 221516 313092 243176 313120
rect 221516 313080 221522 313092
rect 243170 313080 243176 313092
rect 243228 313080 243234 313132
rect 87322 313012 87328 313064
rect 87380 313052 87386 313064
rect 88242 313052 88248 313064
rect 87380 313024 88248 313052
rect 87380 313012 87386 313024
rect 88242 313012 88248 313024
rect 88300 313012 88306 313064
rect 94498 313012 94504 313064
rect 94556 313052 94562 313064
rect 95142 313052 95148 313064
rect 94556 313024 95148 313052
rect 94556 313012 94562 313024
rect 95142 313012 95148 313024
rect 95200 313012 95206 313064
rect 104158 313012 104164 313064
rect 104216 313052 104222 313064
rect 104802 313052 104808 313064
rect 104216 313024 104808 313052
rect 104216 313012 104222 313024
rect 104802 313012 104808 313024
rect 104860 313012 104866 313064
rect 113818 313012 113824 313064
rect 113876 313052 113882 313064
rect 114462 313052 114468 313064
rect 113876 313024 114468 313052
rect 113876 313012 113882 313024
rect 114462 313012 114468 313024
rect 114520 313012 114526 313064
rect 123386 313012 123392 313064
rect 123444 313052 123450 313064
rect 124122 313052 124128 313064
rect 123444 313024 124128 313052
rect 123444 313012 123450 313024
rect 124122 313012 124128 313024
rect 124180 313012 124186 313064
rect 124766 313012 124772 313064
rect 124824 313052 124830 313064
rect 125226 313052 125232 313064
rect 124824 313024 125232 313052
rect 124824 313012 124830 313024
rect 125226 313012 125232 313024
rect 125284 313012 125290 313064
rect 133046 313012 133052 313064
rect 133104 313052 133110 313064
rect 133598 313052 133604 313064
rect 133104 313024 133604 313052
rect 133104 313012 133110 313024
rect 133598 313012 133604 313024
rect 133656 313012 133662 313064
rect 137922 313012 137928 313064
rect 137980 313052 137986 313064
rect 183002 313052 183008 313064
rect 137980 313024 183008 313052
rect 137980 313012 137986 313024
rect 183002 313012 183008 313024
rect 183060 313012 183066 313064
rect 188982 313012 188988 313064
rect 189040 313052 189046 313064
rect 195609 313055 195667 313061
rect 195609 313052 195621 313055
rect 189040 313024 195621 313052
rect 189040 313012 189046 313024
rect 195609 313021 195621 313024
rect 195655 313021 195667 313055
rect 195609 313015 195667 313021
rect 195698 313012 195704 313064
rect 195756 313052 195762 313064
rect 196250 313052 196256 313064
rect 195756 313024 196256 313052
rect 195756 313012 195762 313024
rect 196250 313012 196256 313024
rect 196308 313012 196314 313064
rect 200758 313012 200764 313064
rect 200816 313052 200822 313064
rect 235994 313052 236000 313064
rect 200816 313024 236000 313052
rect 200816 313012 200822 313024
rect 235994 313012 236000 313024
rect 236052 313012 236058 313064
rect 77662 312944 77668 312996
rect 77720 312984 77726 312996
rect 303430 312984 303436 312996
rect 77720 312956 303436 312984
rect 77720 312944 77726 312956
rect 303430 312944 303436 312956
rect 303488 312944 303494 312996
rect 75270 312876 75276 312928
rect 75328 312916 75334 312928
rect 303522 312916 303528 312928
rect 75328 312888 303528 312916
rect 75328 312876 75334 312888
rect 303522 312876 303528 312888
rect 303580 312876 303586 312928
rect 3970 312808 3976 312860
rect 4028 312848 4034 312860
rect 247954 312848 247960 312860
rect 4028 312820 247960 312848
rect 4028 312808 4034 312820
rect 247954 312808 247960 312820
rect 248012 312808 248018 312860
rect 3602 312740 3608 312792
rect 3660 312780 3666 312792
rect 250438 312780 250444 312792
rect 3660 312752 250444 312780
rect 3660 312740 3666 312752
rect 250438 312740 250444 312752
rect 250496 312740 250502 312792
rect 6362 312672 6368 312724
rect 6420 312712 6426 312724
rect 257614 312712 257620 312724
rect 6420 312684 257620 312712
rect 6420 312672 6426 312684
rect 257614 312672 257620 312684
rect 257672 312672 257678 312724
rect 5350 312604 5356 312656
rect 5408 312644 5414 312656
rect 262490 312644 262496 312656
rect 5408 312616 262496 312644
rect 5408 312604 5414 312616
rect 262490 312604 262496 312616
rect 262548 312604 262554 312656
rect 6270 312536 6276 312588
rect 6328 312576 6334 312588
rect 264974 312576 264980 312588
rect 6328 312548 264980 312576
rect 6328 312536 6334 312548
rect 264974 312536 264980 312548
rect 265032 312536 265038 312588
rect 3326 312468 3332 312520
rect 3384 312508 3390 312520
rect 272058 312508 272064 312520
rect 3384 312480 272064 312508
rect 3384 312468 3390 312480
rect 272058 312468 272064 312480
rect 272116 312468 272122 312520
rect 3878 312400 3884 312452
rect 3936 312440 3942 312452
rect 276934 312440 276940 312452
rect 3936 312412 276940 312440
rect 3936 312400 3942 312412
rect 276934 312400 276940 312412
rect 276992 312400 276998 312452
rect 6178 312332 6184 312384
rect 6236 312372 6242 312384
rect 279326 312372 279332 312384
rect 6236 312344 279332 312372
rect 6236 312332 6242 312344
rect 279326 312332 279332 312344
rect 279384 312332 279390 312384
rect 5166 312264 5172 312316
rect 5224 312304 5230 312316
rect 281718 312304 281724 312316
rect 5224 312276 281724 312304
rect 5224 312264 5230 312276
rect 281718 312264 281724 312276
rect 281776 312264 281782 312316
rect 5074 312196 5080 312248
rect 5132 312236 5138 312248
rect 284294 312236 284300 312248
rect 5132 312208 284300 312236
rect 5132 312196 5138 312208
rect 284294 312196 284300 312208
rect 284352 312196 284358 312248
rect 3786 312128 3792 312180
rect 3844 312168 3850 312180
rect 286502 312168 286508 312180
rect 3844 312140 286508 312168
rect 3844 312128 3850 312140
rect 286502 312128 286508 312140
rect 286560 312128 286566 312180
rect 4982 312060 4988 312112
rect 5040 312100 5046 312112
rect 288894 312100 288900 312112
rect 5040 312072 288900 312100
rect 5040 312060 5046 312072
rect 288894 312060 288900 312072
rect 288952 312060 288958 312112
rect 4890 311992 4896 312044
rect 4948 312032 4954 312044
rect 291378 312032 291384 312044
rect 4948 312004 291384 312032
rect 4948 311992 4954 312004
rect 291378 311992 291384 312004
rect 291436 311992 291442 312044
rect 3694 311924 3700 311976
rect 3752 311964 3758 311976
rect 293954 311964 293960 311976
rect 3752 311936 293960 311964
rect 3752 311924 3758 311936
rect 293954 311924 293960 311936
rect 294012 311924 294018 311976
rect 84930 311856 84936 311908
rect 84988 311896 84994 311908
rect 580166 311896 580172 311908
rect 84988 311868 580172 311896
rect 84988 311856 84994 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 31754 310496 31760 310548
rect 31812 310536 31818 310548
rect 302878 310536 302884 310548
rect 31812 310508 302884 310536
rect 31812 310496 31818 310508
rect 302878 310496 302884 310508
rect 302936 310496 302942 310548
rect 79962 310428 79968 310480
rect 80020 310468 80026 310480
rect 304626 310468 304632 310480
rect 80020 310440 304632 310468
rect 80020 310428 80026 310440
rect 304626 310428 304632 310440
rect 304684 310428 304690 310480
rect 65610 310360 65616 310412
rect 65668 310400 65674 310412
rect 65668 310372 70440 310400
rect 65668 310360 65674 310372
rect 60642 310332 60648 310344
rect 60603 310304 60648 310332
rect 60642 310292 60648 310304
rect 60700 310292 60706 310344
rect 63218 310332 63224 310344
rect 63179 310304 63224 310332
rect 63218 310292 63224 310304
rect 63276 310292 63282 310344
rect 70302 310332 70308 310344
rect 70263 310304 70308 310332
rect 70302 310292 70308 310304
rect 70360 310292 70366 310344
rect 70412 310332 70440 310372
rect 72878 310360 72884 310412
rect 72936 310400 72942 310412
rect 304534 310400 304540 310412
rect 72936 310372 304540 310400
rect 72936 310360 72942 310372
rect 304534 310360 304540 310372
rect 304592 310360 304598 310412
rect 303338 310332 303344 310344
rect 70412 310304 303344 310332
rect 303338 310292 303344 310304
rect 303396 310292 303402 310344
rect 55950 310264 55956 310276
rect 55911 310236 55956 310264
rect 55950 310224 55956 310236
rect 56008 310224 56014 310276
rect 58434 310224 58440 310276
rect 58492 310264 58498 310276
rect 303154 310264 303160 310276
rect 58492 310236 303160 310264
rect 58492 310224 58498 310236
rect 303154 310224 303160 310236
rect 303212 310224 303218 310276
rect 39114 310196 39120 310208
rect 39075 310168 39120 310196
rect 39114 310156 39120 310168
rect 39172 310156 39178 310208
rect 41322 310196 41328 310208
rect 41283 310168 41328 310196
rect 41322 310156 41328 310168
rect 41380 310156 41386 310208
rect 46382 310196 46388 310208
rect 46343 310168 46388 310196
rect 46382 310156 46388 310168
rect 46440 310156 46446 310208
rect 48774 310196 48780 310208
rect 48735 310168 48780 310196
rect 48774 310156 48780 310168
rect 48832 310156 48838 310208
rect 53558 310156 53564 310208
rect 53616 310196 53622 310208
rect 304350 310196 304356 310208
rect 53616 310168 304356 310196
rect 53616 310156 53622 310168
rect 304350 310156 304356 310168
rect 304408 310156 304414 310208
rect 4706 310088 4712 310140
rect 4764 310128 4770 310140
rect 255314 310128 255320 310140
rect 4764 310100 255320 310128
rect 4764 310088 4770 310100
rect 255314 310088 255320 310100
rect 255372 310088 255378 310140
rect 5442 310020 5448 310072
rect 5500 310060 5506 310072
rect 260006 310060 260012 310072
rect 5500 310032 260012 310060
rect 5500 310020 5506 310032
rect 260006 310020 260012 310032
rect 260064 310020 260070 310072
rect 304258 310060 304264 310072
rect 296686 310032 304264 310060
rect 5258 309952 5264 310004
rect 5316 309992 5322 310004
rect 267274 309992 267280 310004
rect 5316 309964 267280 309992
rect 5316 309952 5322 309964
rect 267274 309952 267280 309964
rect 267332 309952 267338 310004
rect 269666 309992 269672 310004
rect 269627 309964 269672 309992
rect 269666 309952 269672 309964
rect 269724 309952 269730 310004
rect 274634 309992 274640 310004
rect 274595 309964 274640 309992
rect 274634 309952 274640 309964
rect 274692 309952 274698 310004
rect 296162 309992 296168 310004
rect 296123 309964 296168 309992
rect 296162 309952 296168 309964
rect 296220 309952 296226 310004
rect 39117 309927 39175 309933
rect 39117 309893 39129 309927
rect 39163 309924 39175 309927
rect 296686 309924 296714 310032
rect 304258 310020 304264 310032
rect 304316 310020 304322 310072
rect 298554 309952 298560 310004
rect 298612 309952 298618 310004
rect 39163 309896 296714 309924
rect 39163 309893 39175 309896
rect 39117 309887 39175 309893
rect 4062 309816 4068 309868
rect 4120 309856 4126 309868
rect 269669 309859 269727 309865
rect 269669 309856 269681 309859
rect 4120 309828 269681 309856
rect 4120 309816 4126 309828
rect 269669 309825 269681 309828
rect 269715 309825 269727 309859
rect 269669 309819 269727 309825
rect 3970 309748 3976 309800
rect 4028 309788 4034 309800
rect 274637 309791 274695 309797
rect 274637 309788 274649 309791
rect 4028 309760 274649 309788
rect 4028 309748 4034 309760
rect 274637 309757 274649 309760
rect 274683 309757 274695 309791
rect 274637 309751 274695 309757
rect 3602 309680 3608 309732
rect 3660 309720 3666 309732
rect 296165 309723 296223 309729
rect 296165 309720 296177 309723
rect 3660 309692 296177 309720
rect 3660 309680 3666 309692
rect 296165 309689 296177 309692
rect 296211 309689 296223 309723
rect 296165 309683 296223 309689
rect 3418 309612 3424 309664
rect 3476 309652 3482 309664
rect 298572 309652 298600 309952
rect 3476 309624 298600 309652
rect 3476 309612 3482 309624
rect 70305 309587 70363 309593
rect 70305 309553 70317 309587
rect 70351 309584 70363 309587
rect 580902 309584 580908 309596
rect 70351 309556 580908 309584
rect 70351 309553 70363 309556
rect 70305 309547 70363 309553
rect 580902 309544 580908 309556
rect 580960 309544 580966 309596
rect 63221 309519 63279 309525
rect 63221 309485 63233 309519
rect 63267 309516 63279 309519
rect 580718 309516 580724 309528
rect 63267 309488 580724 309516
rect 63267 309485 63279 309488
rect 63221 309479 63279 309485
rect 580718 309476 580724 309488
rect 580776 309476 580782 309528
rect 60645 309451 60703 309457
rect 60645 309417 60657 309451
rect 60691 309448 60703 309451
rect 580810 309448 580816 309460
rect 60691 309420 580816 309448
rect 60691 309417 60703 309420
rect 60645 309411 60703 309417
rect 580810 309408 580816 309420
rect 580868 309408 580874 309460
rect 55953 309383 56011 309389
rect 55953 309349 55965 309383
rect 55999 309380 56011 309383
rect 580626 309380 580632 309392
rect 55999 309352 580632 309380
rect 55999 309349 56011 309352
rect 55953 309343 56011 309349
rect 580626 309340 580632 309352
rect 580684 309340 580690 309392
rect 48777 309315 48835 309321
rect 48777 309281 48789 309315
rect 48823 309312 48835 309315
rect 580442 309312 580448 309324
rect 48823 309284 580448 309312
rect 48823 309281 48835 309284
rect 48777 309275 48835 309281
rect 580442 309272 580448 309284
rect 580500 309272 580506 309324
rect 46385 309247 46443 309253
rect 46385 309213 46397 309247
rect 46431 309244 46443 309247
rect 580534 309244 580540 309256
rect 46431 309216 580540 309244
rect 46431 309213 46443 309216
rect 46385 309207 46443 309213
rect 580534 309204 580540 309216
rect 580592 309204 580598 309256
rect 41325 309179 41383 309185
rect 41325 309145 41337 309179
rect 41371 309176 41383 309179
rect 580350 309176 580356 309188
rect 41371 309148 580356 309176
rect 41371 309145 41383 309148
rect 41325 309139 41383 309145
rect 580350 309136 580356 309148
rect 580408 309136 580414 309188
rect 2958 306212 2964 306264
rect 3016 306252 3022 306264
rect 6362 306252 6368 306264
rect 3016 306224 6368 306252
rect 3016 306212 3022 306224
rect 6362 306212 6368 306224
rect 6420 306212 6426 306264
rect 304626 299412 304632 299464
rect 304684 299452 304690 299464
rect 580166 299452 580172 299464
rect 304684 299424 580172 299452
rect 304684 299412 304690 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 2774 293224 2780 293276
rect 2832 293264 2838 293276
rect 4706 293264 4712 293276
rect 2832 293236 4712 293264
rect 2832 293224 2838 293236
rect 4706 293224 4712 293236
rect 4764 293224 4770 293276
rect 303522 273164 303528 273216
rect 303580 273204 303586 273216
rect 579982 273204 579988 273216
rect 303580 273176 579988 273204
rect 303580 273164 303586 273176
rect 579982 273164 579988 273176
rect 580040 273164 580046 273216
rect 2774 267180 2780 267232
rect 2832 267220 2838 267232
rect 5442 267220 5448 267232
rect 2832 267192 5448 267220
rect 2832 267180 2838 267192
rect 5442 267180 5448 267192
rect 5500 267180 5506 267232
rect 303430 259360 303436 259412
rect 303488 259400 303494 259412
rect 580166 259400 580172 259412
rect 303488 259372 580172 259400
rect 303488 259360 303494 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3142 255144 3148 255196
rect 3200 255184 3206 255196
rect 6270 255184 6276 255196
rect 3200 255156 6276 255184
rect 3200 255144 3206 255156
rect 6270 255144 6276 255156
rect 6328 255144 6334 255196
rect 304534 245556 304540 245608
rect 304592 245596 304598 245608
rect 580166 245596 580172 245608
rect 304592 245568 580172 245596
rect 304592 245556 304598 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 2774 241068 2780 241120
rect 2832 241108 2838 241120
rect 5350 241108 5356 241120
rect 2832 241080 5356 241108
rect 2832 241068 2838 241080
rect 5350 241068 5356 241080
rect 5408 241068 5414 241120
rect 304442 233180 304448 233232
rect 304500 233220 304506 233232
rect 579982 233220 579988 233232
rect 304500 233192 579988 233220
rect 304500 233180 304506 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 2774 214956 2780 215008
rect 2832 214996 2838 215008
rect 5258 214996 5264 215008
rect 2832 214968 5264 214996
rect 2832 214956 2838 214968
rect 5258 214956 5264 214968
rect 5316 214956 5322 215008
rect 303338 206932 303344 206984
rect 303396 206972 303402 206984
rect 580166 206972 580172 206984
rect 303396 206944 580172 206972
rect 303396 206932 303402 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 303154 166948 303160 167000
rect 303212 166988 303218 167000
rect 579614 166988 579620 167000
rect 303212 166960 579620 166988
rect 303212 166948 303218 166960
rect 579614 166948 579620 166960
rect 579672 166948 579678 167000
rect 304350 153144 304356 153196
rect 304408 153184 304414 153196
rect 579798 153184 579804 153196
rect 304408 153156 579804 153184
rect 304408 153144 304414 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 3142 150220 3148 150272
rect 3200 150260 3206 150272
rect 6178 150260 6184 150272
rect 3200 150232 6184 150260
rect 3200 150220 3206 150232
rect 6178 150220 6184 150232
rect 6236 150220 6242 150272
rect 303246 126896 303252 126948
rect 303304 126936 303310 126948
rect 579706 126936 579712 126948
rect 303304 126908 579712 126936
rect 303304 126896 303310 126908
rect 579706 126896 579712 126908
rect 579764 126896 579770 126948
rect 2774 123836 2780 123888
rect 2832 123876 2838 123888
rect 4798 123876 4804 123888
rect 2832 123848 4804 123876
rect 2832 123836 2838 123848
rect 4798 123836 4804 123848
rect 4856 123836 4862 123888
rect 2774 111460 2780 111512
rect 2832 111500 2838 111512
rect 5166 111500 5172 111512
rect 2832 111472 5172 111500
rect 2832 111460 2838 111472
rect 5166 111460 5172 111472
rect 5224 111460 5230 111512
rect 303062 86912 303068 86964
rect 303120 86952 303126 86964
rect 579614 86952 579620 86964
rect 303120 86924 579620 86952
rect 303120 86912 303126 86924
rect 579614 86912 579620 86924
rect 579672 86912 579678 86964
rect 2774 85144 2780 85196
rect 2832 85184 2838 85196
rect 5074 85184 5080 85196
rect 2832 85156 5080 85184
rect 2832 85144 2838 85156
rect 5074 85144 5080 85156
rect 5132 85144 5138 85196
rect 304258 73108 304264 73160
rect 304316 73148 304322 73160
rect 580166 73148 580172 73160
rect 304316 73120 580172 73148
rect 304316 73108 304322 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 2774 71612 2780 71664
rect 2832 71652 2838 71664
rect 4982 71652 4988 71664
rect 2832 71624 4988 71652
rect 2832 71612 2838 71624
rect 4982 71612 4988 71624
rect 5040 71612 5046 71664
rect 302970 46860 302976 46912
rect 303028 46900 303034 46912
rect 580166 46900 580172 46912
rect 303028 46872 580172 46900
rect 303028 46860 303034 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 2774 45500 2780 45552
rect 2832 45540 2838 45552
rect 4890 45540 4896 45552
rect 2832 45512 4896 45540
rect 2832 45500 2838 45512
rect 4890 45500 4896 45512
rect 4948 45500 4954 45552
rect 302878 33056 302884 33108
rect 302936 33096 302942 33108
rect 580166 33096 580172 33108
rect 302936 33068 580172 33096
rect 302936 33056 302942 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 250806 31764 250812 31816
rect 250864 31804 250870 31816
rect 251082 31804 251088 31816
rect 250864 31776 251088 31804
rect 250864 31764 250870 31776
rect 251082 31764 251088 31776
rect 251140 31764 251146 31816
rect 261938 31764 261944 31816
rect 261996 31804 262002 31816
rect 262122 31804 262128 31816
rect 261996 31776 262128 31804
rect 261996 31764 262002 31776
rect 262122 31764 262128 31776
rect 262180 31764 262186 31816
rect 264698 31764 264704 31816
rect 264756 31804 264762 31816
rect 264882 31804 264888 31816
rect 264756 31776 264888 31804
rect 264756 31764 264762 31776
rect 264882 31764 264888 31776
rect 264940 31764 264946 31816
rect 20530 31696 20536 31748
rect 20588 31736 20594 31748
rect 37366 31736 37372 31748
rect 20588 31708 37372 31736
rect 20588 31696 20594 31708
rect 37366 31696 37372 31708
rect 37424 31696 37430 31748
rect 41322 31696 41328 31748
rect 41380 31736 41386 31748
rect 46934 31736 46940 31748
rect 41380 31708 46940 31736
rect 41380 31696 41386 31708
rect 46934 31696 46940 31708
rect 46992 31696 46998 31748
rect 88150 31696 88156 31748
rect 88208 31736 88214 31748
rect 127158 31736 127164 31748
rect 88208 31708 127164 31736
rect 88208 31696 88214 31708
rect 127158 31696 127164 31708
rect 127216 31696 127222 31748
rect 200758 31736 200764 31748
rect 186286 31708 200764 31736
rect 19242 31628 19248 31680
rect 19300 31668 19306 31680
rect 36262 31668 36268 31680
rect 19300 31640 36268 31668
rect 19300 31628 19306 31640
rect 36262 31628 36268 31640
rect 36320 31628 36326 31680
rect 44082 31628 44088 31680
rect 44140 31668 44146 31680
rect 47946 31668 47952 31680
rect 44140 31640 47952 31668
rect 44140 31628 44146 31640
rect 47946 31628 47952 31640
rect 48004 31628 48010 31680
rect 68830 31628 68836 31680
rect 68888 31668 68894 31680
rect 68888 31640 75040 31668
rect 68888 31628 68894 31640
rect 16482 31560 16488 31612
rect 16540 31600 16546 31612
rect 35158 31600 35164 31612
rect 16540 31572 35164 31600
rect 16540 31560 16546 31572
rect 35158 31560 35164 31572
rect 35216 31560 35222 31612
rect 42702 31560 42708 31612
rect 42760 31600 42766 31612
rect 47394 31600 47400 31612
rect 42760 31572 47400 31600
rect 42760 31560 42766 31572
rect 47394 31560 47400 31572
rect 47452 31560 47458 31612
rect 75012 31600 75040 31640
rect 83182 31628 83188 31680
rect 83240 31668 83246 31680
rect 90266 31668 90272 31680
rect 83240 31640 90272 31668
rect 83240 31628 83246 31640
rect 90266 31628 90272 31640
rect 90324 31628 90330 31680
rect 90358 31628 90364 31680
rect 90416 31668 90422 31680
rect 94498 31668 94504 31680
rect 90416 31640 94504 31668
rect 90416 31628 90422 31640
rect 94498 31628 94504 31640
rect 94556 31628 94562 31680
rect 108942 31628 108948 31680
rect 109000 31668 109006 31680
rect 159358 31668 159364 31680
rect 109000 31640 159364 31668
rect 109000 31628 109006 31640
rect 159358 31628 159364 31640
rect 159416 31628 159422 31680
rect 162210 31628 162216 31680
rect 162268 31668 162274 31680
rect 186286 31668 186314 31708
rect 200758 31696 200764 31708
rect 200816 31696 200822 31748
rect 215662 31696 215668 31748
rect 215720 31736 215726 31748
rect 358078 31736 358084 31748
rect 215720 31708 358084 31736
rect 215720 31696 215726 31708
rect 358078 31696 358084 31708
rect 358136 31696 358142 31748
rect 162268 31640 186314 31668
rect 162268 31628 162274 31640
rect 202322 31628 202328 31680
rect 202380 31668 202386 31680
rect 344278 31668 344284 31680
rect 202380 31640 344284 31668
rect 202380 31628 202386 31640
rect 344278 31628 344284 31640
rect 344336 31628 344342 31680
rect 85758 31600 85764 31612
rect 75012 31572 85764 31600
rect 85758 31560 85764 31572
rect 85816 31560 85822 31612
rect 93670 31560 93676 31612
rect 93728 31600 93734 31612
rect 95878 31600 95884 31612
rect 93728 31572 95884 31600
rect 93728 31560 93734 31572
rect 95878 31560 95884 31572
rect 95936 31560 95942 31612
rect 114833 31603 114891 31609
rect 114833 31569 114845 31603
rect 114879 31600 114891 31603
rect 157978 31600 157984 31612
rect 114879 31572 157984 31600
rect 114879 31569 114891 31572
rect 114833 31563 114891 31569
rect 157978 31560 157984 31572
rect 158036 31560 158042 31612
rect 188982 31560 188988 31612
rect 189040 31600 189046 31612
rect 330478 31600 330484 31612
rect 189040 31572 330484 31600
rect 189040 31560 189046 31572
rect 330478 31560 330484 31572
rect 330536 31560 330542 31612
rect 13722 31492 13728 31544
rect 13780 31532 13786 31544
rect 34054 31532 34060 31544
rect 13780 31504 34060 31532
rect 13780 31492 13786 31504
rect 34054 31492 34060 31504
rect 34112 31492 34118 31544
rect 72602 31492 72608 31544
rect 72660 31532 72666 31544
rect 87506 31532 87512 31544
rect 72660 31504 87512 31532
rect 72660 31492 72666 31504
rect 87506 31492 87512 31504
rect 87564 31492 87570 31544
rect 104342 31492 104348 31544
rect 104400 31532 104406 31544
rect 155218 31532 155224 31544
rect 104400 31504 155224 31532
rect 104400 31492 104406 31504
rect 155218 31492 155224 31504
rect 155276 31492 155282 31544
rect 166902 31492 166908 31544
rect 166960 31532 166966 31544
rect 208946 31532 208952 31544
rect 166960 31504 208952 31532
rect 166960 31492 166966 31504
rect 208946 31492 208952 31504
rect 209004 31492 209010 31544
rect 362218 31532 362224 31544
rect 219406 31504 362224 31532
rect 15102 31424 15108 31476
rect 15160 31464 15166 31476
rect 34606 31464 34612 31476
rect 15160 31436 34612 31464
rect 15160 31424 15166 31436
rect 34606 31424 34612 31436
rect 34664 31424 34670 31476
rect 38562 31424 38568 31476
rect 38620 31464 38626 31476
rect 45738 31464 45744 31476
rect 38620 31436 45744 31464
rect 38620 31424 38626 31436
rect 45738 31424 45744 31436
rect 45796 31424 45802 31476
rect 86494 31424 86500 31476
rect 86552 31464 86558 31476
rect 101398 31464 101404 31476
rect 86552 31436 101404 31464
rect 86552 31424 86558 31436
rect 101398 31424 101404 31436
rect 101456 31424 101462 31476
rect 105998 31424 106004 31476
rect 106056 31464 106062 31476
rect 156598 31464 156604 31476
rect 106056 31436 156604 31464
rect 106056 31424 106062 31436
rect 156598 31424 156604 31436
rect 156656 31424 156662 31476
rect 168926 31424 168932 31476
rect 168984 31464 168990 31476
rect 213178 31464 213184 31476
rect 168984 31436 213184 31464
rect 168984 31424 168990 31436
rect 213178 31424 213184 31436
rect 213236 31424 213242 31476
rect 219066 31424 219072 31476
rect 219124 31464 219130 31476
rect 219406 31464 219434 31504
rect 362218 31492 362224 31504
rect 362276 31492 362282 31544
rect 219124 31436 219434 31464
rect 219124 31424 219130 31436
rect 237926 31424 237932 31476
rect 237984 31464 237990 31476
rect 238662 31464 238668 31476
rect 237984 31436 238668 31464
rect 237984 31424 237990 31436
rect 238662 31424 238668 31436
rect 238720 31424 238726 31476
rect 238757 31467 238815 31473
rect 238757 31433 238769 31467
rect 238803 31464 238815 31467
rect 376018 31464 376024 31476
rect 238803 31436 376024 31464
rect 238803 31433 238815 31436
rect 238757 31427 238815 31433
rect 376018 31424 376024 31436
rect 376076 31424 376082 31476
rect 10962 31356 10968 31408
rect 11020 31396 11026 31408
rect 32398 31396 32404 31408
rect 11020 31368 32404 31396
rect 11020 31356 11026 31368
rect 32398 31356 32404 31368
rect 32456 31356 32462 31408
rect 70946 31356 70952 31408
rect 71004 31396 71010 31408
rect 88978 31396 88984 31408
rect 71004 31368 88984 31396
rect 71004 31356 71010 31368
rect 88978 31356 88984 31368
rect 89036 31356 89042 31408
rect 107562 31356 107568 31408
rect 107620 31396 107626 31408
rect 114833 31399 114891 31405
rect 114833 31396 114845 31399
rect 107620 31368 114845 31396
rect 107620 31356 107626 31368
rect 114833 31365 114845 31368
rect 114879 31365 114891 31399
rect 114833 31359 114891 31365
rect 127437 31399 127495 31405
rect 127437 31365 127449 31399
rect 127483 31396 127495 31399
rect 170398 31396 170404 31408
rect 127483 31368 170404 31396
rect 127483 31365 127495 31368
rect 127437 31359 127495 31365
rect 170398 31356 170404 31368
rect 170456 31356 170462 31408
rect 225690 31356 225696 31408
rect 225748 31396 225754 31408
rect 369118 31396 369124 31408
rect 225748 31368 369124 31396
rect 225748 31356 225754 31368
rect 369118 31356 369124 31368
rect 369176 31356 369182 31408
rect 12342 31288 12348 31340
rect 12400 31328 12406 31340
rect 33134 31328 33140 31340
rect 12400 31300 33140 31328
rect 12400 31288 12406 31300
rect 33134 31288 33140 31300
rect 33192 31288 33198 31340
rect 34422 31288 34428 31340
rect 34480 31328 34486 31340
rect 43530 31328 43536 31340
rect 34480 31300 43536 31328
rect 34480 31288 34486 31300
rect 43530 31288 43536 31300
rect 43588 31288 43594 31340
rect 84838 31288 84844 31340
rect 84896 31328 84902 31340
rect 105538 31328 105544 31340
rect 84896 31300 105544 31328
rect 84896 31288 84902 31300
rect 105538 31288 105544 31300
rect 105596 31288 105602 31340
rect 119338 31288 119344 31340
rect 119396 31328 119402 31340
rect 173158 31328 173164 31340
rect 119396 31300 173164 31328
rect 119396 31288 119402 31300
rect 173158 31288 173164 31300
rect 173216 31288 173222 31340
rect 212350 31288 212356 31340
rect 212408 31328 212414 31340
rect 355318 31328 355324 31340
rect 212408 31300 355324 31328
rect 212408 31288 212414 31300
rect 355318 31288 355324 31300
rect 355376 31288 355382 31340
rect 9582 31220 9588 31272
rect 9640 31260 9646 31272
rect 31846 31260 31852 31272
rect 9640 31232 31852 31260
rect 9640 31220 9646 31232
rect 31846 31220 31852 31232
rect 31904 31220 31910 31272
rect 35802 31220 35808 31272
rect 35860 31260 35866 31272
rect 44174 31260 44180 31272
rect 35860 31232 44180 31260
rect 35860 31220 35866 31232
rect 44174 31220 44180 31232
rect 44232 31220 44238 31272
rect 45462 31220 45468 31272
rect 45520 31260 45526 31272
rect 48498 31260 48504 31272
rect 45520 31232 48504 31260
rect 45520 31220 45526 31232
rect 48498 31220 48504 31232
rect 48556 31220 48562 31272
rect 77018 31220 77024 31272
rect 77076 31260 77082 31272
rect 102318 31260 102324 31272
rect 77076 31232 102324 31260
rect 77076 31220 77082 31232
rect 102318 31220 102324 31232
rect 102376 31220 102382 31272
rect 114370 31220 114376 31272
rect 114428 31260 114434 31272
rect 167638 31260 167644 31272
rect 114428 31232 167644 31260
rect 114428 31220 114434 31232
rect 167638 31220 167644 31232
rect 167696 31220 167702 31272
rect 205542 31220 205548 31272
rect 205600 31260 205606 31272
rect 348418 31260 348424 31272
rect 205600 31232 348424 31260
rect 205600 31220 205606 31232
rect 348418 31220 348424 31232
rect 348476 31220 348482 31272
rect 6822 31152 6828 31204
rect 6880 31192 6886 31204
rect 30742 31192 30748 31204
rect 6880 31164 30748 31192
rect 6880 31152 6886 31164
rect 30742 31152 30748 31164
rect 30800 31152 30806 31204
rect 33042 31152 33048 31204
rect 33100 31192 33106 31204
rect 42978 31192 42984 31204
rect 33100 31164 42984 31192
rect 33100 31152 33106 31164
rect 42978 31152 42984 31164
rect 43036 31152 43042 31204
rect 78582 31152 78588 31204
rect 78640 31192 78646 31204
rect 94409 31195 94467 31201
rect 94409 31192 94421 31195
rect 78640 31164 94421 31192
rect 78640 31152 78646 31164
rect 94409 31161 94421 31164
rect 94455 31161 94467 31195
rect 94409 31155 94467 31161
rect 112622 31152 112628 31204
rect 112680 31192 112686 31204
rect 166258 31192 166264 31204
rect 112680 31164 166264 31192
rect 112680 31152 112686 31164
rect 166258 31152 166264 31164
rect 166316 31152 166322 31204
rect 198642 31152 198648 31204
rect 198700 31192 198706 31204
rect 341518 31192 341524 31204
rect 198700 31164 341524 31192
rect 198700 31152 198706 31164
rect 341518 31152 341524 31164
rect 341576 31152 341582 31204
rect 4062 31084 4068 31136
rect 4120 31124 4126 31136
rect 29638 31124 29644 31136
rect 4120 31096 29644 31124
rect 4120 31084 4126 31096
rect 29638 31084 29644 31096
rect 29696 31084 29702 31136
rect 30282 31084 30288 31136
rect 30340 31124 30346 31136
rect 41874 31124 41880 31136
rect 30340 31096 41880 31124
rect 30340 31084 30346 31096
rect 41874 31084 41880 31096
rect 41932 31084 41938 31136
rect 45370 31084 45376 31136
rect 45428 31124 45434 31136
rect 49142 31124 49148 31136
rect 45428 31096 49148 31124
rect 45428 31084 45434 31096
rect 49142 31084 49148 31096
rect 49200 31084 49206 31136
rect 82078 31084 82084 31136
rect 82136 31124 82142 31136
rect 108298 31124 108304 31136
rect 82136 31096 108304 31124
rect 82136 31084 82142 31096
rect 108298 31084 108304 31096
rect 108356 31084 108362 31136
rect 115842 31084 115848 31136
rect 115900 31124 115906 31136
rect 169018 31124 169024 31136
rect 115900 31096 169024 31124
rect 115900 31084 115906 31096
rect 169018 31084 169024 31096
rect 169076 31084 169082 31136
rect 222010 31084 222016 31136
rect 222068 31124 222074 31136
rect 366358 31124 366364 31136
rect 222068 31096 366364 31124
rect 222068 31084 222074 31096
rect 366358 31084 366364 31096
rect 366416 31084 366422 31136
rect 5442 31016 5448 31068
rect 5500 31056 5506 31068
rect 30374 31056 30380 31068
rect 5500 31028 30380 31056
rect 5500 31016 5506 31028
rect 30374 31016 30380 31028
rect 30432 31016 30438 31068
rect 31662 31016 31668 31068
rect 31720 31056 31726 31068
rect 42426 31056 42432 31068
rect 31720 31028 42432 31056
rect 31720 31016 31726 31028
rect 42426 31016 42432 31028
rect 42484 31016 42490 31068
rect 67542 31016 67548 31068
rect 67600 31056 67606 31068
rect 82998 31056 83004 31068
rect 67600 31028 83004 31056
rect 67600 31016 67606 31028
rect 82998 31016 83004 31028
rect 83056 31016 83062 31068
rect 85390 31016 85396 31068
rect 85448 31056 85454 31068
rect 119338 31056 119344 31068
rect 85448 31028 119344 31056
rect 85448 31016 85454 31028
rect 119338 31016 119344 31028
rect 119396 31016 119402 31068
rect 120994 31016 121000 31068
rect 121052 31056 121058 31068
rect 175918 31056 175924 31068
rect 121052 31028 175924 31056
rect 121052 31016 121058 31028
rect 175918 31016 175924 31028
rect 175976 31016 175982 31068
rect 180518 31016 180524 31068
rect 180576 31056 180582 31068
rect 185486 31056 185492 31068
rect 180576 31028 185492 31056
rect 180576 31016 180582 31028
rect 185486 31016 185492 31028
rect 185544 31016 185550 31068
rect 228910 31016 228916 31068
rect 228968 31056 228974 31068
rect 373258 31056 373264 31068
rect 228968 31028 373264 31056
rect 228968 31016 228974 31028
rect 373258 31016 373264 31028
rect 373316 31016 373322 31068
rect 23382 30948 23388 31000
rect 23440 30988 23446 31000
rect 38654 30988 38660 31000
rect 23440 30960 38660 30988
rect 23440 30948 23446 30960
rect 38654 30948 38660 30960
rect 38712 30948 38718 31000
rect 39942 30948 39948 31000
rect 40000 30988 40006 31000
rect 46290 30988 46296 31000
rect 40000 30960 46296 30988
rect 40000 30948 40006 30960
rect 46290 30948 46296 30960
rect 46348 30948 46354 31000
rect 94409 30991 94467 30997
rect 94409 30957 94421 30991
rect 94455 30988 94467 30991
rect 104158 30988 104164 31000
rect 94455 30960 104164 30988
rect 94455 30957 94467 30960
rect 94409 30951 94467 30957
rect 104158 30948 104164 30960
rect 104216 30948 104222 31000
rect 110966 30948 110972 31000
rect 111024 30988 111030 31000
rect 160738 30988 160744 31000
rect 111024 30960 160744 30988
rect 111024 30948 111030 30960
rect 160738 30948 160744 30960
rect 160796 30948 160802 31000
rect 195606 30948 195612 31000
rect 195664 30988 195670 31000
rect 337378 30988 337384 31000
rect 195664 30960 337384 30988
rect 195664 30948 195670 30960
rect 337378 30948 337384 30960
rect 337436 30948 337442 31000
rect 20622 30880 20628 30932
rect 20680 30920 20686 30932
rect 36814 30920 36820 30932
rect 20680 30892 36820 30920
rect 20680 30880 20686 30892
rect 36814 30880 36820 30892
rect 36872 30880 36878 30932
rect 92290 30880 92296 30932
rect 92348 30920 92354 30932
rect 135438 30920 135444 30932
rect 92348 30892 135444 30920
rect 92348 30880 92354 30892
rect 135438 30880 135444 30892
rect 135496 30880 135502 30932
rect 179966 30920 179972 30932
rect 142126 30892 179972 30920
rect 22002 30812 22008 30864
rect 22060 30852 22066 30864
rect 37918 30852 37924 30864
rect 22060 30824 37924 30852
rect 22060 30812 22066 30824
rect 37918 30812 37924 30824
rect 37976 30812 37982 30864
rect 90910 30812 90916 30864
rect 90968 30852 90974 30864
rect 132494 30852 132500 30864
rect 90968 30824 132500 30852
rect 90968 30812 90974 30824
rect 132494 30812 132500 30824
rect 132552 30812 132558 30864
rect 137922 30812 137928 30864
rect 137980 30852 137986 30864
rect 142126 30852 142154 30892
rect 179966 30880 179972 30892
rect 180024 30880 180030 30932
rect 192294 30880 192300 30932
rect 192352 30920 192358 30932
rect 200577 30923 200635 30929
rect 192352 30892 195974 30920
rect 192352 30880 192358 30892
rect 177390 30852 177396 30864
rect 137980 30824 142154 30852
rect 151786 30824 177396 30852
rect 137980 30812 137986 30824
rect 24762 30744 24768 30796
rect 24820 30784 24826 30796
rect 39114 30784 39120 30796
rect 24820 30756 39120 30784
rect 24820 30744 24826 30756
rect 39114 30744 39120 30756
rect 39172 30744 39178 30796
rect 102042 30744 102048 30796
rect 102100 30784 102106 30796
rect 142798 30784 142804 30796
rect 102100 30756 142804 30784
rect 102100 30744 102106 30756
rect 142798 30744 142804 30756
rect 142856 30744 142862 30796
rect 28902 30676 28908 30728
rect 28960 30716 28966 30728
rect 41414 30716 41420 30728
rect 28960 30688 41420 30716
rect 28960 30676 28966 30688
rect 41414 30676 41420 30688
rect 41472 30676 41478 30728
rect 89622 30676 89628 30728
rect 89680 30716 89686 30728
rect 129734 30716 129740 30728
rect 89680 30688 129740 30716
rect 89680 30676 89686 30688
rect 129734 30676 129740 30688
rect 129792 30676 129798 30728
rect 136542 30676 136548 30728
rect 136600 30716 136606 30728
rect 151786 30716 151814 30824
rect 177390 30812 177396 30824
rect 177448 30812 177454 30864
rect 185578 30812 185584 30864
rect 185636 30852 185642 30864
rect 185636 30824 186314 30852
rect 185636 30812 185642 30824
rect 172238 30744 172244 30796
rect 172296 30784 172302 30796
rect 179325 30787 179383 30793
rect 179325 30784 179337 30787
rect 172296 30756 179337 30784
rect 172296 30744 172302 30756
rect 179325 30753 179337 30756
rect 179371 30753 179383 30787
rect 179325 30747 179383 30753
rect 180058 30744 180064 30796
rect 180116 30784 180122 30796
rect 180702 30784 180708 30796
rect 180116 30756 180708 30784
rect 180116 30744 180122 30756
rect 180702 30744 180708 30756
rect 180760 30744 180766 30796
rect 181162 30744 181168 30796
rect 181220 30784 181226 30796
rect 182082 30784 182088 30796
rect 181220 30756 182088 30784
rect 181220 30744 181226 30756
rect 182082 30744 182088 30756
rect 182140 30744 182146 30796
rect 183922 30744 183928 30796
rect 183980 30784 183986 30796
rect 184842 30784 184848 30796
rect 183980 30756 184848 30784
rect 183980 30744 183986 30756
rect 184842 30744 184848 30756
rect 184900 30744 184906 30796
rect 186286 30784 186314 30824
rect 187326 30812 187332 30864
rect 187384 30852 187390 30864
rect 187602 30852 187608 30864
rect 187384 30824 187608 30852
rect 187384 30812 187390 30824
rect 187602 30812 187608 30824
rect 187660 30812 187666 30864
rect 189534 30812 189540 30864
rect 189592 30852 189598 30864
rect 190270 30852 190276 30864
rect 189592 30824 190276 30852
rect 189592 30812 189598 30824
rect 190270 30812 190276 30824
rect 190328 30812 190334 30864
rect 191190 30812 191196 30864
rect 191248 30852 191254 30864
rect 191742 30852 191748 30864
rect 191248 30824 191748 30852
rect 191248 30812 191254 30824
rect 191742 30812 191748 30824
rect 191800 30812 191806 30864
rect 193950 30812 193956 30864
rect 194008 30852 194014 30864
rect 194502 30852 194508 30864
rect 194008 30824 194508 30852
rect 194008 30812 194014 30824
rect 194502 30812 194508 30824
rect 194560 30812 194566 30864
rect 195946 30852 195974 30892
rect 200577 30889 200589 30923
rect 200623 30920 200635 30923
rect 204898 30920 204904 30932
rect 200623 30892 204904 30920
rect 200623 30889 200635 30892
rect 200577 30883 200635 30889
rect 204898 30880 204904 30892
rect 204956 30880 204962 30932
rect 209038 30880 209044 30932
rect 209096 30920 209102 30932
rect 351178 30920 351184 30932
rect 209096 30892 351184 30920
rect 209096 30880 209102 30892
rect 351178 30880 351184 30892
rect 351236 30880 351242 30932
rect 333238 30852 333244 30864
rect 195946 30824 333244 30852
rect 333238 30812 333244 30824
rect 333296 30812 333302 30864
rect 323670 30784 323676 30796
rect 186286 30756 323676 30784
rect 323670 30744 323676 30756
rect 323728 30744 323734 30796
rect 136600 30688 151814 30716
rect 136600 30676 136606 30688
rect 175182 30676 175188 30728
rect 175240 30716 175246 30728
rect 301498 30716 301504 30728
rect 175240 30688 301504 30716
rect 175240 30676 175246 30688
rect 301498 30676 301504 30688
rect 301556 30676 301562 30728
rect 27522 30608 27528 30660
rect 27580 30648 27586 30660
rect 40218 30648 40224 30660
rect 27580 30620 40224 30648
rect 27580 30608 27586 30620
rect 40218 30608 40224 30620
rect 40276 30608 40282 30660
rect 117682 30608 117688 30660
rect 117740 30648 117746 30660
rect 127437 30651 127495 30657
rect 127437 30648 127449 30651
rect 117740 30620 127449 30648
rect 117740 30608 117746 30620
rect 127437 30617 127449 30620
rect 127483 30617 127495 30651
rect 127437 30611 127495 30617
rect 128262 30608 128268 30660
rect 128320 30648 128326 30660
rect 177206 30648 177212 30660
rect 128320 30620 177212 30648
rect 128320 30608 128326 30620
rect 177206 30608 177212 30620
rect 177264 30608 177270 30660
rect 178954 30608 178960 30660
rect 179012 30648 179018 30660
rect 179012 30620 269620 30648
rect 179012 30608 179018 30620
rect 26142 30540 26148 30592
rect 26200 30580 26206 30592
rect 39666 30580 39672 30592
rect 26200 30552 39672 30580
rect 26200 30540 26206 30552
rect 39666 30540 39672 30552
rect 39724 30540 39730 30592
rect 139946 30540 139952 30592
rect 140004 30580 140010 30592
rect 181438 30580 181444 30592
rect 140004 30552 181444 30580
rect 140004 30540 140010 30552
rect 181438 30540 181444 30552
rect 181496 30540 181502 30592
rect 182818 30540 182824 30592
rect 182876 30580 182882 30592
rect 183462 30580 183468 30592
rect 182876 30552 183468 30580
rect 182876 30540 182882 30552
rect 183462 30540 183468 30552
rect 183520 30540 183526 30592
rect 184474 30540 184480 30592
rect 184532 30580 184538 30592
rect 184750 30580 184756 30592
rect 184532 30552 184756 30580
rect 184532 30540 184538 30552
rect 184750 30540 184756 30552
rect 184808 30540 184814 30592
rect 186682 30540 186688 30592
rect 186740 30580 186746 30592
rect 187418 30580 187424 30592
rect 186740 30552 187424 30580
rect 186740 30540 186746 30552
rect 187418 30540 187424 30552
rect 187476 30540 187482 30592
rect 188430 30540 188436 30592
rect 188488 30580 188494 30592
rect 188982 30580 188988 30592
rect 188488 30552 188988 30580
rect 188488 30540 188494 30552
rect 188982 30540 188988 30552
rect 189040 30540 189046 30592
rect 192846 30540 192852 30592
rect 192904 30580 192910 30592
rect 193122 30580 193128 30592
rect 192904 30552 193128 30580
rect 192904 30540 192910 30552
rect 193122 30540 193128 30552
rect 193180 30540 193186 30592
rect 195054 30540 195060 30592
rect 195112 30580 195118 30592
rect 195790 30580 195796 30592
rect 195112 30552 195796 30580
rect 195112 30540 195118 30552
rect 195790 30540 195796 30552
rect 195848 30540 195854 30592
rect 196710 30540 196716 30592
rect 196768 30580 196774 30592
rect 197170 30580 197176 30592
rect 196768 30552 197176 30580
rect 196768 30540 196774 30552
rect 197170 30540 197176 30552
rect 197228 30540 197234 30592
rect 197906 30540 197912 30592
rect 197964 30580 197970 30592
rect 198642 30580 198648 30592
rect 197964 30552 198648 30580
rect 197964 30540 197970 30552
rect 198642 30540 198648 30552
rect 198700 30540 198706 30592
rect 199562 30540 199568 30592
rect 199620 30580 199626 30592
rect 200022 30580 200028 30592
rect 199620 30552 200028 30580
rect 199620 30540 199626 30552
rect 200022 30540 200028 30552
rect 200080 30540 200086 30592
rect 203426 30540 203432 30592
rect 203484 30580 203490 30592
rect 204070 30580 204076 30592
rect 203484 30552 204076 30580
rect 203484 30540 203490 30552
rect 204070 30540 204076 30552
rect 204128 30540 204134 30592
rect 210694 30540 210700 30592
rect 210752 30580 210758 30592
rect 211062 30580 211068 30592
rect 210752 30552 211068 30580
rect 210752 30540 210758 30552
rect 211062 30540 211068 30552
rect 211120 30540 211126 30592
rect 224034 30540 224040 30592
rect 224092 30580 224098 30592
rect 224862 30580 224868 30592
rect 224092 30552 224868 30580
rect 224092 30540 224098 30552
rect 224862 30540 224868 30552
rect 224920 30540 224926 30592
rect 227346 30540 227352 30592
rect 227404 30580 227410 30592
rect 227622 30580 227628 30592
rect 227404 30552 227628 30580
rect 227404 30540 227410 30552
rect 227622 30540 227628 30552
rect 227680 30540 227686 30592
rect 232406 30540 232412 30592
rect 232464 30580 232470 30592
rect 238757 30583 238815 30589
rect 238757 30580 238769 30583
rect 232464 30552 238769 30580
rect 232464 30540 232470 30552
rect 238757 30549 238769 30552
rect 238803 30549 238815 30583
rect 238757 30543 238815 30549
rect 239493 30583 239551 30589
rect 239493 30549 239505 30583
rect 239539 30580 239551 30583
rect 269393 30583 269451 30589
rect 269393 30580 269405 30583
rect 239539 30552 269405 30580
rect 239539 30549 239551 30552
rect 239493 30543 239551 30549
rect 269393 30549 269405 30552
rect 269439 30549 269451 30583
rect 269393 30543 269451 30549
rect 28810 30472 28816 30524
rect 28868 30512 28874 30524
rect 40770 30512 40776 30524
rect 28868 30484 40776 30512
rect 28868 30472 28874 30484
rect 40770 30472 40776 30484
rect 40828 30472 40834 30524
rect 49602 30472 49608 30524
rect 49660 30512 49666 30524
rect 51074 30512 51080 30524
rect 49660 30484 51080 30512
rect 49660 30472 49666 30484
rect 51074 30472 51080 30484
rect 51132 30472 51138 30524
rect 171686 30472 171692 30524
rect 171744 30512 171750 30524
rect 172422 30512 172428 30524
rect 171744 30484 172428 30512
rect 171744 30472 171750 30484
rect 172422 30472 172428 30484
rect 172480 30472 172486 30524
rect 173342 30472 173348 30524
rect 173400 30512 173406 30524
rect 173802 30512 173808 30524
rect 173400 30484 173808 30512
rect 173400 30472 173406 30484
rect 173802 30472 173808 30484
rect 173860 30472 173866 30524
rect 174446 30472 174452 30524
rect 174504 30512 174510 30524
rect 174998 30512 175004 30524
rect 174504 30484 175004 30512
rect 174504 30472 174510 30484
rect 174998 30472 175004 30484
rect 175056 30472 175062 30524
rect 177298 30472 177304 30524
rect 177356 30512 177362 30524
rect 177850 30512 177856 30524
rect 177356 30484 177856 30512
rect 177356 30472 177362 30484
rect 177850 30472 177856 30484
rect 177908 30472 177914 30524
rect 178402 30472 178408 30524
rect 178460 30512 178466 30524
rect 179230 30512 179236 30524
rect 178460 30484 179236 30512
rect 178460 30472 178466 30484
rect 179230 30472 179236 30484
rect 179288 30472 179294 30524
rect 179325 30515 179383 30521
rect 179325 30481 179337 30515
rect 179371 30512 179383 30515
rect 244918 30512 244924 30524
rect 179371 30484 244924 30512
rect 179371 30481 179383 30484
rect 179325 30475 179383 30481
rect 244918 30472 244924 30484
rect 244976 30472 244982 30524
rect 248233 30515 248291 30521
rect 248233 30512 248245 30515
rect 245396 30484 248245 30512
rect 37090 30404 37096 30456
rect 37148 30444 37154 30456
rect 45186 30444 45192 30456
rect 37148 30416 45192 30444
rect 37148 30404 37154 30416
rect 45186 30404 45192 30416
rect 45244 30404 45250 30456
rect 46842 30404 46848 30456
rect 46900 30444 46906 30456
rect 49694 30444 49700 30456
rect 46900 30416 49700 30444
rect 46900 30404 46906 30416
rect 49694 30404 49700 30416
rect 49752 30404 49758 30456
rect 56962 30404 56968 30456
rect 57020 30444 57026 30456
rect 57882 30444 57888 30456
rect 57020 30416 57888 30444
rect 57020 30404 57026 30416
rect 57882 30404 57888 30416
rect 57940 30404 57946 30456
rect 59722 30404 59728 30456
rect 59780 30444 59786 30456
rect 60642 30444 60648 30456
rect 59780 30416 60648 30444
rect 59780 30404 59786 30416
rect 60642 30404 60648 30416
rect 60700 30404 60706 30456
rect 79226 30404 79232 30456
rect 79284 30444 79290 30456
rect 79870 30444 79876 30456
rect 79284 30416 79876 30444
rect 79284 30404 79290 30416
rect 79870 30404 79876 30416
rect 79928 30404 79934 30456
rect 88702 30404 88708 30456
rect 88760 30444 88766 30456
rect 93118 30444 93124 30456
rect 88760 30416 93124 30444
rect 88760 30404 88766 30416
rect 93118 30404 93124 30416
rect 93176 30404 93182 30456
rect 97074 30404 97080 30456
rect 97132 30444 97138 30456
rect 97902 30444 97908 30456
rect 97132 30416 97908 30444
rect 97132 30404 97138 30416
rect 97902 30404 97908 30416
rect 97960 30404 97966 30456
rect 100294 30404 100300 30456
rect 100352 30444 100358 30456
rect 100662 30444 100668 30456
rect 100352 30416 100668 30444
rect 100352 30404 100358 30416
rect 100662 30404 100668 30416
rect 100720 30404 100726 30456
rect 123846 30404 123852 30456
rect 123904 30444 123910 30456
rect 124122 30444 124128 30456
rect 123904 30416 124128 30444
rect 123904 30404 123910 30416
rect 124122 30404 124128 30416
rect 124180 30404 124186 30456
rect 128814 30404 128820 30456
rect 128872 30444 128878 30456
rect 129642 30444 129648 30456
rect 128872 30416 129648 30444
rect 128872 30404 128878 30416
rect 129642 30404 129648 30416
rect 129700 30404 129706 30456
rect 132126 30404 132132 30456
rect 132184 30444 132190 30456
rect 132402 30444 132408 30456
rect 132184 30416 132408 30444
rect 132184 30404 132190 30416
rect 132402 30404 132408 30416
rect 132460 30404 132466 30456
rect 149422 30404 149428 30456
rect 149480 30444 149486 30456
rect 150342 30444 150348 30456
rect 149480 30416 150348 30444
rect 149480 30404 149486 30416
rect 150342 30404 150348 30416
rect 150400 30404 150406 30456
rect 152734 30404 152740 30456
rect 152792 30444 152798 30456
rect 153102 30444 153108 30456
rect 152792 30416 153108 30444
rect 152792 30404 152798 30416
rect 153102 30404 153108 30416
rect 153160 30404 153166 30456
rect 158346 30404 158352 30456
rect 158404 30444 158410 30456
rect 158622 30444 158628 30456
rect 158404 30416 158628 30444
rect 158404 30404 158410 30416
rect 158622 30404 158628 30416
rect 158680 30404 158686 30456
rect 161106 30404 161112 30456
rect 161164 30444 161170 30456
rect 161382 30444 161388 30456
rect 161164 30416 161388 30444
rect 161164 30404 161170 30416
rect 161382 30404 161388 30416
rect 161440 30404 161446 30456
rect 163314 30404 163320 30456
rect 163372 30444 163378 30456
rect 164142 30444 164148 30456
rect 163372 30416 164148 30444
rect 163372 30404 163378 30416
rect 164142 30404 164148 30416
rect 164200 30404 164206 30456
rect 165430 30404 165436 30456
rect 165488 30444 165494 30456
rect 165488 30416 168236 30444
rect 165488 30404 165494 30416
rect 37182 30336 37188 30388
rect 37240 30376 37246 30388
rect 44634 30376 44640 30388
rect 37240 30348 44640 30376
rect 37240 30336 37246 30348
rect 44634 30336 44640 30348
rect 44692 30336 44698 30388
rect 48222 30336 48228 30388
rect 48280 30376 48286 30388
rect 50246 30376 50252 30388
rect 48280 30348 50252 30376
rect 48280 30336 48286 30348
rect 50246 30336 50252 30348
rect 50304 30336 50310 30388
rect 52454 30336 52460 30388
rect 52512 30376 52518 30388
rect 53006 30376 53012 30388
rect 52512 30348 53012 30376
rect 52512 30336 52518 30348
rect 53006 30336 53012 30348
rect 53064 30336 53070 30388
rect 55858 30336 55864 30388
rect 55916 30376 55922 30388
rect 56502 30376 56508 30388
rect 55916 30348 56508 30376
rect 55916 30336 55922 30348
rect 56502 30336 56508 30348
rect 56560 30336 56566 30388
rect 57514 30336 57520 30388
rect 57572 30376 57578 30388
rect 57790 30376 57796 30388
rect 57572 30348 57796 30376
rect 57572 30336 57578 30348
rect 57790 30336 57796 30348
rect 57848 30336 57854 30388
rect 58618 30336 58624 30388
rect 58676 30376 58682 30388
rect 59262 30376 59268 30388
rect 58676 30348 59268 30376
rect 58676 30336 58682 30348
rect 59262 30336 59268 30348
rect 59320 30336 59326 30388
rect 60366 30336 60372 30388
rect 60424 30376 60430 30388
rect 60550 30376 60556 30388
rect 60424 30348 60556 30376
rect 60424 30336 60430 30348
rect 60550 30336 60556 30348
rect 60608 30336 60614 30388
rect 61470 30336 61476 30388
rect 61528 30376 61534 30388
rect 61930 30376 61936 30388
rect 61528 30348 61936 30376
rect 61528 30336 61534 30348
rect 61930 30336 61936 30348
rect 61988 30336 61994 30388
rect 62574 30336 62580 30388
rect 62632 30376 62638 30388
rect 63402 30376 63408 30388
rect 62632 30348 63408 30376
rect 62632 30336 62638 30348
rect 63402 30336 63408 30348
rect 63460 30336 63466 30388
rect 64230 30336 64236 30388
rect 64288 30376 64294 30388
rect 64690 30376 64696 30388
rect 64288 30348 64696 30376
rect 64288 30336 64294 30348
rect 64690 30336 64696 30348
rect 64748 30336 64754 30388
rect 65334 30336 65340 30388
rect 65392 30376 65398 30388
rect 65886 30376 65892 30388
rect 65392 30348 65892 30376
rect 65392 30336 65398 30348
rect 65886 30336 65892 30348
rect 65944 30336 65950 30388
rect 66990 30336 66996 30388
rect 67048 30376 67054 30388
rect 67542 30376 67548 30388
rect 67048 30348 67548 30376
rect 67048 30336 67054 30348
rect 67542 30336 67548 30348
rect 67600 30336 67606 30388
rect 68094 30336 68100 30388
rect 68152 30376 68158 30388
rect 68922 30376 68928 30388
rect 68152 30348 68928 30376
rect 68152 30336 68158 30348
rect 68922 30336 68928 30348
rect 68980 30336 68986 30388
rect 69750 30336 69756 30388
rect 69808 30376 69814 30388
rect 70302 30376 70308 30388
rect 69808 30348 70308 30376
rect 69808 30336 69814 30348
rect 70302 30336 70308 30348
rect 70360 30336 70366 30388
rect 73706 30336 73712 30388
rect 73764 30376 73770 30388
rect 74442 30376 74448 30388
rect 73764 30348 74448 30376
rect 73764 30336 73770 30348
rect 74442 30336 74448 30348
rect 74500 30336 74506 30388
rect 75362 30336 75368 30388
rect 75420 30376 75426 30388
rect 75822 30376 75828 30388
rect 75420 30348 75828 30376
rect 75420 30336 75426 30348
rect 75822 30336 75828 30348
rect 75880 30336 75886 30388
rect 76466 30336 76472 30388
rect 76524 30376 76530 30388
rect 77202 30376 77208 30388
rect 76524 30348 77208 30376
rect 76524 30336 76530 30348
rect 77202 30336 77208 30348
rect 77260 30336 77266 30388
rect 78122 30336 78128 30388
rect 78180 30376 78186 30388
rect 78582 30376 78588 30388
rect 78180 30348 78588 30376
rect 78180 30336 78186 30348
rect 78582 30336 78588 30348
rect 78640 30336 78646 30388
rect 79686 30336 79692 30388
rect 79744 30376 79750 30388
rect 79962 30376 79968 30388
rect 79744 30348 79968 30376
rect 79744 30336 79750 30348
rect 79962 30336 79968 30348
rect 80020 30336 80026 30388
rect 85942 30336 85948 30388
rect 86000 30376 86006 30388
rect 86770 30376 86776 30388
rect 86000 30348 86776 30376
rect 86000 30336 86006 30348
rect 86770 30336 86776 30348
rect 86828 30336 86834 30388
rect 87598 30336 87604 30388
rect 87656 30376 87662 30388
rect 88242 30376 88248 30388
rect 87656 30348 88248 30376
rect 87656 30336 87662 30348
rect 88242 30336 88248 30348
rect 88300 30336 88306 30388
rect 91462 30336 91468 30388
rect 91520 30376 91526 30388
rect 92290 30376 92296 30388
rect 91520 30348 92296 30376
rect 91520 30336 91526 30348
rect 92290 30336 92296 30348
rect 92348 30336 92354 30388
rect 93210 30336 93216 30388
rect 93268 30376 93274 30388
rect 93762 30376 93768 30388
rect 93268 30348 93768 30376
rect 93268 30336 93274 30348
rect 93762 30336 93768 30348
rect 93820 30336 93826 30388
rect 94314 30336 94320 30388
rect 94372 30376 94378 30388
rect 94866 30376 94872 30388
rect 94372 30348 94872 30376
rect 94372 30336 94378 30348
rect 94866 30336 94872 30348
rect 94924 30336 94930 30388
rect 95970 30336 95976 30388
rect 96028 30376 96034 30388
rect 96522 30376 96528 30388
rect 96028 30348 96528 30376
rect 96028 30336 96034 30348
rect 96522 30336 96528 30348
rect 96580 30336 96586 30388
rect 97626 30336 97632 30388
rect 97684 30376 97690 30388
rect 97810 30376 97816 30388
rect 97684 30348 97816 30376
rect 97684 30336 97690 30348
rect 97810 30336 97816 30348
rect 97868 30336 97874 30388
rect 98730 30336 98736 30388
rect 98788 30376 98794 30388
rect 99282 30376 99288 30388
rect 98788 30348 99288 30376
rect 98788 30336 98794 30348
rect 99282 30336 99288 30348
rect 99340 30336 99346 30388
rect 99834 30336 99840 30388
rect 99892 30376 99898 30388
rect 100570 30376 100576 30388
rect 99892 30348 100576 30376
rect 99892 30336 99898 30348
rect 100570 30336 100576 30348
rect 100628 30336 100634 30388
rect 101490 30336 101496 30388
rect 101548 30376 101554 30388
rect 102042 30376 102048 30388
rect 101548 30348 102048 30376
rect 101548 30336 101554 30348
rect 102042 30336 102048 30348
rect 102100 30336 102106 30388
rect 102686 30336 102692 30388
rect 102744 30376 102750 30388
rect 103238 30376 103244 30388
rect 102744 30348 103244 30376
rect 102744 30336 102750 30348
rect 103238 30336 103244 30348
rect 103296 30336 103302 30388
rect 105446 30336 105452 30388
rect 105504 30376 105510 30388
rect 106182 30376 106188 30388
rect 105504 30348 106188 30376
rect 105504 30336 105510 30348
rect 106182 30336 106188 30348
rect 106240 30336 106246 30388
rect 107102 30336 107108 30388
rect 107160 30376 107166 30388
rect 107562 30376 107568 30388
rect 107160 30348 107568 30376
rect 107160 30336 107166 30348
rect 107562 30336 107568 30348
rect 107620 30336 107626 30388
rect 108206 30336 108212 30388
rect 108264 30376 108270 30388
rect 108942 30376 108948 30388
rect 108264 30348 108948 30376
rect 108264 30336 108270 30348
rect 108942 30336 108948 30348
rect 109000 30336 109006 30388
rect 113818 30336 113824 30388
rect 113876 30376 113882 30388
rect 114462 30376 114468 30388
rect 113876 30348 114468 30376
rect 113876 30336 113882 30348
rect 114462 30336 114468 30348
rect 114520 30336 114526 30388
rect 114922 30336 114928 30388
rect 114980 30376 114986 30388
rect 115474 30376 115480 30388
rect 114980 30348 115480 30376
rect 114980 30336 114986 30348
rect 115474 30336 115480 30348
rect 115532 30336 115538 30388
rect 116578 30336 116584 30388
rect 116636 30376 116642 30388
rect 117130 30376 117136 30388
rect 116636 30348 117136 30376
rect 116636 30336 116642 30348
rect 117130 30336 117136 30348
rect 117188 30336 117194 30388
rect 120442 30336 120448 30388
rect 120500 30376 120506 30388
rect 121362 30376 121368 30388
rect 120500 30348 121368 30376
rect 120500 30336 120506 30348
rect 121362 30336 121368 30348
rect 121420 30336 121426 30388
rect 122098 30336 122104 30388
rect 122156 30376 122162 30388
rect 122742 30376 122748 30388
rect 122156 30348 122748 30376
rect 122156 30336 122162 30348
rect 122742 30336 122748 30348
rect 122800 30336 122806 30388
rect 123202 30336 123208 30388
rect 123260 30376 123266 30388
rect 123938 30376 123944 30388
rect 123260 30348 123944 30376
rect 123260 30336 123266 30348
rect 123938 30336 123944 30348
rect 123996 30336 124002 30388
rect 124950 30336 124956 30388
rect 125008 30376 125014 30388
rect 125410 30376 125416 30388
rect 125008 30348 125416 30376
rect 125008 30336 125014 30348
rect 125410 30336 125416 30348
rect 125468 30336 125474 30388
rect 126054 30336 126060 30388
rect 126112 30376 126118 30388
rect 126790 30376 126796 30388
rect 126112 30348 126796 30376
rect 126112 30336 126118 30348
rect 126790 30336 126796 30348
rect 126848 30336 126854 30388
rect 127710 30336 127716 30388
rect 127768 30376 127774 30388
rect 128262 30376 128268 30388
rect 127768 30348 128268 30376
rect 127768 30336 127774 30348
rect 128262 30336 128268 30348
rect 128320 30336 128326 30388
rect 129366 30336 129372 30388
rect 129424 30376 129430 30388
rect 129550 30376 129556 30388
rect 129424 30348 129556 30376
rect 129424 30336 129430 30348
rect 129550 30336 129556 30348
rect 129608 30336 129614 30388
rect 130470 30336 130476 30388
rect 130528 30376 130534 30388
rect 131022 30376 131028 30388
rect 130528 30348 131028 30376
rect 130528 30336 130534 30348
rect 131022 30336 131028 30348
rect 131080 30336 131086 30388
rect 131574 30336 131580 30388
rect 131632 30376 131638 30388
rect 132218 30376 132224 30388
rect 131632 30348 132224 30376
rect 131632 30336 131638 30348
rect 132218 30336 132224 30348
rect 132276 30336 132282 30388
rect 133230 30336 133236 30388
rect 133288 30376 133294 30388
rect 133690 30376 133696 30388
rect 133288 30348 133696 30376
rect 133288 30336 133294 30348
rect 133690 30336 133696 30348
rect 133748 30336 133754 30388
rect 134426 30336 134432 30388
rect 134484 30376 134490 30388
rect 135070 30376 135076 30388
rect 134484 30348 135076 30376
rect 134484 30336 134490 30348
rect 135070 30336 135076 30348
rect 135128 30336 135134 30388
rect 136082 30336 136088 30388
rect 136140 30376 136146 30388
rect 136542 30376 136548 30388
rect 136140 30348 136548 30376
rect 136140 30336 136146 30348
rect 136542 30336 136548 30348
rect 136600 30336 136606 30388
rect 137186 30336 137192 30388
rect 137244 30376 137250 30388
rect 137922 30376 137928 30388
rect 137244 30348 137928 30376
rect 137244 30336 137250 30348
rect 137922 30336 137928 30348
rect 137980 30336 137986 30388
rect 140498 30336 140504 30388
rect 140556 30376 140562 30388
rect 140682 30376 140688 30388
rect 140556 30348 140688 30376
rect 140556 30336 140562 30348
rect 140682 30336 140688 30348
rect 140740 30336 140746 30388
rect 141602 30336 141608 30388
rect 141660 30376 141666 30388
rect 142062 30376 142068 30388
rect 141660 30348 142068 30376
rect 141660 30336 141666 30348
rect 142062 30336 142068 30348
rect 142120 30336 142126 30388
rect 142706 30336 142712 30388
rect 142764 30376 142770 30388
rect 142764 30348 143212 30376
rect 142764 30336 142770 30348
rect 143184 30240 143212 30348
rect 143258 30336 143264 30388
rect 143316 30376 143322 30388
rect 143442 30376 143448 30388
rect 143316 30348 143448 30376
rect 143316 30336 143322 30348
rect 143442 30336 143448 30348
rect 143500 30336 143506 30388
rect 144362 30336 144368 30388
rect 144420 30376 144426 30388
rect 144822 30376 144828 30388
rect 144420 30348 144828 30376
rect 144420 30336 144426 30348
rect 144822 30336 144828 30348
rect 144880 30336 144886 30388
rect 145558 30336 145564 30388
rect 145616 30376 145622 30388
rect 146110 30376 146116 30388
rect 145616 30348 146116 30376
rect 145616 30336 145622 30348
rect 146110 30336 146116 30348
rect 146168 30336 146174 30388
rect 146662 30336 146668 30388
rect 146720 30376 146726 30388
rect 147490 30376 147496 30388
rect 146720 30348 147496 30376
rect 146720 30336 146726 30348
rect 147490 30336 147496 30348
rect 147548 30336 147554 30388
rect 148318 30336 148324 30388
rect 148376 30376 148382 30388
rect 148962 30376 148968 30388
rect 148376 30348 148968 30376
rect 148376 30336 148382 30348
rect 148962 30336 148968 30348
rect 149020 30336 149026 30388
rect 149974 30336 149980 30388
rect 150032 30376 150038 30388
rect 150250 30376 150256 30388
rect 150032 30348 150256 30376
rect 150032 30336 150038 30348
rect 150250 30336 150256 30348
rect 150308 30336 150314 30388
rect 151078 30336 151084 30388
rect 151136 30376 151142 30388
rect 151722 30376 151728 30388
rect 151136 30348 151728 30376
rect 151136 30336 151142 30348
rect 151722 30336 151728 30348
rect 151780 30336 151786 30388
rect 152182 30336 152188 30388
rect 152240 30376 152246 30388
rect 152918 30376 152924 30388
rect 152240 30348 152924 30376
rect 152240 30336 152246 30348
rect 152918 30336 152924 30348
rect 152976 30336 152982 30388
rect 153838 30336 153844 30388
rect 153896 30376 153902 30388
rect 154390 30376 154396 30388
rect 153896 30348 154396 30376
rect 153896 30336 153902 30348
rect 154390 30336 154396 30348
rect 154448 30336 154454 30388
rect 154942 30336 154948 30388
rect 155000 30376 155006 30388
rect 155770 30376 155776 30388
rect 155000 30348 155776 30376
rect 155000 30336 155006 30348
rect 155770 30336 155776 30348
rect 155828 30336 155834 30388
rect 156690 30336 156696 30388
rect 156748 30376 156754 30388
rect 157242 30376 157248 30388
rect 156748 30348 157248 30376
rect 156748 30336 156754 30348
rect 157242 30336 157248 30348
rect 157300 30336 157306 30388
rect 157794 30336 157800 30388
rect 157852 30376 157858 30388
rect 158438 30376 158444 30388
rect 157852 30348 158444 30376
rect 157852 30336 157858 30348
rect 158438 30336 158444 30348
rect 158496 30336 158502 30388
rect 159450 30336 159456 30388
rect 159508 30376 159514 30388
rect 159910 30376 159916 30388
rect 159508 30348 159916 30376
rect 159508 30336 159514 30348
rect 159910 30336 159916 30348
rect 159968 30336 159974 30388
rect 160554 30336 160560 30388
rect 160612 30376 160618 30388
rect 161198 30376 161204 30388
rect 160612 30348 161204 30376
rect 160612 30336 160618 30348
rect 161198 30336 161204 30348
rect 161256 30336 161262 30388
rect 163866 30336 163872 30388
rect 163924 30376 163930 30388
rect 164050 30376 164056 30388
rect 163924 30348 164056 30376
rect 163924 30336 163930 30348
rect 164050 30336 164056 30348
rect 164108 30336 164114 30388
rect 164970 30336 164976 30388
rect 165028 30376 165034 30388
rect 165522 30376 165528 30388
rect 165028 30348 165528 30376
rect 165028 30336 165034 30348
rect 165522 30336 165528 30348
rect 165580 30336 165586 30388
rect 166166 30336 166172 30388
rect 166224 30376 166230 30388
rect 166902 30376 166908 30388
rect 166224 30348 166908 30376
rect 166224 30336 166230 30348
rect 166902 30336 166908 30348
rect 166960 30336 166966 30388
rect 168208 30376 168236 30416
rect 170582 30404 170588 30456
rect 170640 30444 170646 30456
rect 242158 30444 242164 30456
rect 170640 30416 242164 30444
rect 170640 30404 170646 30416
rect 242158 30404 242164 30416
rect 242216 30404 242222 30456
rect 242434 30404 242440 30456
rect 242492 30444 242498 30456
rect 245396 30444 245424 30484
rect 248233 30481 248245 30484
rect 248279 30481 248291 30515
rect 248233 30475 248291 30481
rect 250162 30472 250168 30524
rect 250220 30512 250226 30524
rect 250990 30512 250996 30524
rect 250220 30484 250996 30512
rect 250220 30472 250226 30484
rect 250990 30472 250996 30484
rect 251048 30472 251054 30524
rect 251910 30472 251916 30524
rect 251968 30512 251974 30524
rect 252462 30512 252468 30524
rect 251968 30484 252468 30512
rect 251968 30472 251974 30484
rect 252462 30472 252468 30484
rect 252520 30472 252526 30524
rect 253014 30472 253020 30524
rect 253072 30512 253078 30524
rect 253566 30512 253572 30524
rect 253072 30484 253572 30512
rect 253072 30472 253078 30484
rect 253566 30472 253572 30484
rect 253624 30472 253630 30524
rect 254670 30472 254676 30524
rect 254728 30512 254734 30524
rect 255130 30512 255136 30524
rect 254728 30484 255136 30512
rect 254728 30472 254734 30484
rect 255130 30472 255136 30484
rect 255188 30472 255194 30524
rect 255774 30472 255780 30524
rect 255832 30512 255838 30524
rect 256510 30512 256516 30524
rect 255832 30484 256516 30512
rect 255832 30472 255838 30484
rect 256510 30472 256516 30484
rect 256568 30472 256574 30524
rect 257430 30472 257436 30524
rect 257488 30512 257494 30524
rect 257982 30512 257988 30524
rect 257488 30484 257988 30512
rect 257488 30472 257494 30484
rect 257982 30472 257988 30484
rect 258040 30472 258046 30524
rect 259086 30472 259092 30524
rect 259144 30512 259150 30524
rect 259270 30512 259276 30524
rect 259144 30484 259276 30512
rect 259144 30472 259150 30484
rect 259270 30472 259276 30484
rect 259328 30472 259334 30524
rect 260190 30472 260196 30524
rect 260248 30512 260254 30524
rect 260742 30512 260748 30524
rect 260248 30484 260748 30512
rect 260248 30472 260254 30484
rect 260742 30472 260748 30484
rect 260800 30472 260806 30524
rect 261386 30472 261392 30524
rect 261444 30512 261450 30524
rect 261938 30512 261944 30524
rect 261444 30484 261944 30512
rect 261444 30472 261450 30484
rect 261938 30472 261944 30484
rect 261996 30472 262002 30524
rect 263042 30472 263048 30524
rect 263100 30512 263106 30524
rect 263502 30512 263508 30524
rect 263100 30484 263508 30512
rect 263100 30472 263106 30484
rect 263502 30472 263508 30484
rect 263560 30472 263566 30524
rect 264146 30472 264152 30524
rect 264204 30512 264210 30524
rect 264698 30512 264704 30524
rect 264204 30484 264704 30512
rect 264204 30472 264210 30484
rect 264698 30472 264704 30484
rect 264756 30472 264762 30524
rect 266906 30472 266912 30524
rect 266964 30512 266970 30524
rect 267550 30512 267556 30524
rect 266964 30484 267556 30512
rect 266964 30472 266970 30484
rect 267550 30472 267556 30484
rect 267608 30472 267614 30524
rect 268562 30472 268568 30524
rect 268620 30512 268626 30524
rect 269022 30512 269028 30524
rect 268620 30484 269028 30512
rect 268620 30472 268626 30484
rect 269022 30472 269028 30484
rect 269080 30472 269086 30524
rect 269592 30512 269620 30620
rect 269666 30608 269672 30660
rect 269724 30648 269730 30660
rect 270494 30648 270500 30660
rect 269724 30620 270500 30648
rect 269724 30608 269730 30620
rect 270494 30608 270500 30620
rect 270552 30608 270558 30660
rect 270589 30651 270647 30657
rect 270589 30617 270601 30651
rect 270635 30648 270647 30651
rect 276290 30648 276296 30660
rect 270635 30620 276296 30648
rect 270635 30617 270647 30620
rect 270589 30611 270647 30617
rect 276290 30608 276296 30620
rect 276348 30608 276354 30660
rect 276382 30608 276388 30660
rect 276440 30648 276446 30660
rect 277302 30648 277308 30660
rect 276440 30620 277308 30648
rect 276440 30608 276446 30620
rect 277302 30608 277308 30620
rect 277360 30608 277366 30660
rect 279694 30608 279700 30660
rect 279752 30648 279758 30660
rect 280062 30648 280068 30660
rect 279752 30620 280068 30648
rect 279752 30608 279758 30620
rect 280062 30608 280068 30620
rect 280120 30608 280126 30660
rect 284754 30608 284760 30660
rect 284812 30648 284818 30660
rect 285582 30648 285588 30660
rect 284812 30620 285588 30648
rect 284812 30608 284818 30620
rect 285582 30608 285588 30620
rect 285640 30608 285646 30660
rect 288066 30608 288072 30660
rect 288124 30648 288130 30660
rect 288342 30648 288348 30660
rect 288124 30620 288348 30648
rect 288124 30608 288130 30620
rect 288342 30608 288348 30620
rect 288400 30608 288406 30660
rect 293126 30608 293132 30660
rect 293184 30648 293190 30660
rect 293954 30648 293960 30660
rect 293184 30620 293960 30648
rect 293184 30608 293190 30620
rect 293954 30608 293960 30620
rect 294012 30608 294018 30660
rect 301406 30608 301412 30660
rect 301464 30648 301470 30660
rect 308398 30648 308404 30660
rect 301464 30620 308404 30648
rect 301464 30608 301470 30620
rect 308398 30608 308404 30620
rect 308456 30608 308462 30660
rect 269761 30583 269819 30589
rect 269761 30549 269773 30583
rect 269807 30580 269819 30583
rect 309778 30580 309784 30592
rect 269807 30552 309784 30580
rect 269807 30549 269819 30552
rect 269761 30543 269819 30549
rect 309778 30540 309784 30552
rect 309836 30540 309842 30592
rect 270129 30515 270187 30521
rect 270129 30512 270141 30515
rect 269592 30484 270141 30512
rect 270129 30481 270141 30484
rect 270175 30481 270187 30515
rect 270129 30475 270187 30481
rect 270218 30472 270224 30524
rect 270276 30512 270282 30524
rect 270402 30512 270408 30524
rect 270276 30484 270408 30512
rect 270276 30472 270282 30484
rect 270402 30472 270408 30484
rect 270460 30472 270466 30524
rect 271322 30472 271328 30524
rect 271380 30512 271386 30524
rect 271782 30512 271788 30524
rect 271380 30484 271788 30512
rect 271380 30472 271386 30484
rect 271782 30472 271788 30484
rect 271840 30472 271846 30524
rect 272518 30472 272524 30524
rect 272576 30512 272582 30524
rect 273070 30512 273076 30524
rect 272576 30484 273076 30512
rect 272576 30472 272582 30484
rect 273070 30472 273076 30484
rect 273128 30472 273134 30524
rect 273622 30472 273628 30524
rect 273680 30512 273686 30524
rect 274450 30512 274456 30524
rect 273680 30484 274456 30512
rect 273680 30472 273686 30484
rect 274450 30472 274456 30484
rect 274508 30472 274514 30524
rect 275278 30472 275284 30524
rect 275336 30512 275342 30524
rect 275922 30512 275928 30524
rect 275336 30484 275928 30512
rect 275336 30472 275342 30484
rect 275922 30472 275928 30484
rect 275980 30472 275986 30524
rect 276934 30472 276940 30524
rect 276992 30512 276998 30524
rect 277210 30512 277216 30524
rect 276992 30484 277216 30512
rect 276992 30472 276998 30484
rect 277210 30472 277216 30484
rect 277268 30472 277274 30524
rect 278038 30472 278044 30524
rect 278096 30512 278102 30524
rect 278682 30512 278688 30524
rect 278096 30484 278688 30512
rect 278096 30472 278102 30484
rect 278682 30472 278688 30484
rect 278740 30472 278746 30524
rect 279142 30472 279148 30524
rect 279200 30512 279206 30524
rect 279878 30512 279884 30524
rect 279200 30484 279884 30512
rect 279200 30472 279206 30484
rect 279878 30472 279884 30484
rect 279936 30472 279942 30524
rect 280798 30472 280804 30524
rect 280856 30512 280862 30524
rect 281350 30512 281356 30524
rect 280856 30484 281356 30512
rect 280856 30472 280862 30484
rect 281350 30472 281356 30484
rect 281408 30472 281414 30524
rect 281902 30472 281908 30524
rect 281960 30512 281966 30524
rect 282730 30512 282736 30524
rect 281960 30484 282736 30512
rect 281960 30472 281966 30484
rect 282730 30472 282736 30484
rect 282788 30472 282794 30524
rect 283650 30472 283656 30524
rect 283708 30512 283714 30524
rect 284202 30512 284208 30524
rect 283708 30484 284208 30512
rect 283708 30472 283714 30484
rect 284202 30472 284208 30484
rect 284260 30472 284266 30524
rect 285306 30472 285312 30524
rect 285364 30512 285370 30524
rect 285490 30512 285496 30524
rect 285364 30484 285496 30512
rect 285364 30472 285370 30484
rect 285490 30472 285496 30484
rect 285548 30472 285554 30524
rect 286410 30472 286416 30524
rect 286468 30512 286474 30524
rect 286962 30512 286968 30524
rect 286468 30484 286968 30512
rect 286468 30472 286474 30484
rect 286962 30472 286968 30484
rect 287020 30472 287026 30524
rect 287514 30472 287520 30524
rect 287572 30512 287578 30524
rect 288158 30512 288164 30524
rect 287572 30484 288164 30512
rect 287572 30472 287578 30484
rect 288158 30472 288164 30484
rect 288216 30472 288222 30524
rect 289170 30472 289176 30524
rect 289228 30512 289234 30524
rect 289630 30512 289636 30524
rect 289228 30484 289636 30512
rect 289228 30472 289234 30484
rect 289630 30472 289636 30484
rect 289688 30472 289694 30524
rect 290274 30472 290280 30524
rect 290332 30512 290338 30524
rect 291010 30512 291016 30524
rect 290332 30484 291016 30512
rect 290332 30472 290338 30484
rect 291010 30472 291016 30484
rect 291068 30472 291074 30524
rect 291930 30472 291936 30524
rect 291988 30512 291994 30524
rect 292390 30512 292396 30524
rect 291988 30484 292396 30512
rect 291988 30472 291994 30484
rect 292390 30472 292396 30484
rect 292448 30472 292454 30524
rect 293678 30472 293684 30524
rect 293736 30512 293742 30524
rect 293862 30512 293868 30524
rect 293736 30484 293868 30512
rect 293736 30472 293742 30484
rect 293862 30472 293868 30484
rect 293920 30472 293926 30524
rect 294782 30472 294788 30524
rect 294840 30512 294846 30524
rect 295242 30512 295248 30524
rect 294840 30484 295248 30512
rect 294840 30472 294846 30484
rect 295242 30472 295248 30484
rect 295300 30472 295306 30524
rect 295886 30472 295892 30524
rect 295944 30512 295950 30524
rect 296438 30512 296444 30524
rect 295944 30484 296444 30512
rect 295944 30472 295950 30484
rect 296438 30472 296444 30484
rect 296496 30472 296502 30524
rect 298646 30472 298652 30524
rect 298704 30512 298710 30524
rect 299290 30512 299296 30524
rect 298704 30484 299296 30512
rect 298704 30472 298710 30484
rect 299290 30472 299296 30484
rect 299348 30472 299354 30524
rect 301958 30472 301964 30524
rect 302016 30512 302022 30524
rect 304258 30512 304264 30524
rect 302016 30484 304264 30512
rect 302016 30472 302022 30484
rect 304258 30472 304264 30484
rect 304316 30472 304322 30524
rect 242492 30416 245424 30444
rect 242492 30404 242498 30416
rect 245470 30404 245476 30456
rect 245528 30444 245534 30456
rect 315390 30444 315396 30456
rect 245528 30416 315396 30444
rect 245528 30404 245534 30416
rect 315390 30404 315396 30416
rect 315448 30404 315454 30456
rect 200577 30379 200635 30385
rect 200577 30376 200589 30379
rect 168208 30348 200589 30376
rect 200577 30345 200589 30348
rect 200623 30345 200635 30379
rect 200577 30339 200635 30345
rect 200666 30336 200672 30388
rect 200724 30376 200730 30388
rect 200724 30348 201172 30376
rect 200724 30336 200730 30348
rect 143442 30240 143448 30252
rect 143184 30212 143448 30240
rect 143442 30200 143448 30212
rect 143500 30200 143506 30252
rect 201144 30240 201172 30348
rect 201218 30336 201224 30388
rect 201276 30376 201282 30388
rect 201402 30376 201408 30388
rect 201276 30348 201408 30376
rect 201276 30336 201282 30348
rect 201402 30336 201408 30348
rect 201460 30336 201466 30388
rect 203886 30336 203892 30388
rect 203944 30376 203950 30388
rect 204162 30376 204168 30388
rect 203944 30348 204168 30376
rect 203944 30336 203950 30348
rect 204162 30336 204168 30348
rect 204220 30336 204226 30388
rect 205082 30336 205088 30388
rect 205140 30376 205146 30388
rect 205542 30376 205548 30388
rect 205140 30348 205548 30376
rect 205140 30336 205146 30348
rect 205542 30336 205548 30348
rect 205600 30336 205606 30388
rect 206186 30336 206192 30388
rect 206244 30376 206250 30388
rect 206738 30376 206744 30388
rect 206244 30348 206744 30376
rect 206244 30336 206250 30348
rect 206738 30336 206744 30348
rect 206796 30336 206802 30388
rect 210142 30336 210148 30388
rect 210200 30376 210206 30388
rect 210878 30376 210884 30388
rect 210200 30348 210884 30376
rect 210200 30336 210206 30348
rect 210878 30336 210884 30348
rect 210936 30336 210942 30388
rect 211798 30336 211804 30388
rect 211856 30376 211862 30388
rect 212442 30376 212448 30388
rect 211856 30348 212448 30376
rect 211856 30336 211862 30348
rect 212442 30336 212448 30348
rect 212500 30336 212506 30388
rect 212902 30336 212908 30388
rect 212960 30376 212966 30388
rect 213730 30376 213736 30388
rect 212960 30348 213736 30376
rect 212960 30336 212966 30348
rect 213730 30336 213736 30348
rect 213788 30336 213794 30388
rect 214558 30336 214564 30388
rect 214616 30376 214622 30388
rect 215202 30376 215208 30388
rect 214616 30348 215208 30376
rect 214616 30336 214622 30348
rect 215202 30336 215208 30348
rect 215260 30336 215266 30388
rect 216214 30336 216220 30388
rect 216272 30376 216278 30388
rect 216582 30376 216588 30388
rect 216272 30348 216588 30376
rect 216272 30336 216278 30348
rect 216582 30336 216588 30348
rect 216640 30336 216646 30388
rect 217318 30336 217324 30388
rect 217376 30376 217382 30388
rect 217962 30376 217968 30388
rect 217376 30348 217968 30376
rect 217376 30336 217382 30348
rect 217962 30336 217968 30348
rect 218020 30336 218026 30388
rect 218422 30336 218428 30388
rect 218480 30376 218486 30388
rect 219250 30376 219256 30388
rect 218480 30348 219256 30376
rect 218480 30336 218486 30348
rect 219250 30336 219256 30348
rect 219308 30336 219314 30388
rect 220170 30336 220176 30388
rect 220228 30376 220234 30388
rect 220630 30376 220636 30388
rect 220228 30348 220636 30376
rect 220228 30336 220234 30348
rect 220630 30336 220636 30348
rect 220688 30336 220694 30388
rect 221274 30336 221280 30388
rect 221332 30376 221338 30388
rect 222102 30376 222108 30388
rect 221332 30348 222108 30376
rect 221332 30336 221338 30348
rect 222102 30336 222108 30348
rect 222160 30336 222166 30388
rect 222930 30336 222936 30388
rect 222988 30376 222994 30388
rect 223482 30376 223488 30388
rect 222988 30348 223488 30376
rect 222988 30336 222994 30348
rect 223482 30336 223488 30348
rect 223540 30336 223546 30388
rect 224586 30336 224592 30388
rect 224644 30376 224650 30388
rect 224770 30376 224776 30388
rect 224644 30348 224776 30376
rect 224644 30336 224650 30348
rect 224770 30336 224776 30348
rect 224828 30336 224834 30388
rect 226794 30336 226800 30388
rect 226852 30376 226858 30388
rect 227438 30376 227444 30388
rect 226852 30348 227444 30376
rect 226852 30336 226858 30348
rect 227438 30336 227444 30348
rect 227496 30336 227502 30388
rect 228450 30336 228456 30388
rect 228508 30376 228514 30388
rect 229002 30376 229008 30388
rect 228508 30348 229008 30376
rect 228508 30336 228514 30348
rect 229002 30336 229008 30348
rect 229060 30336 229066 30388
rect 229646 30336 229652 30388
rect 229704 30376 229710 30388
rect 230290 30376 230296 30388
rect 229704 30348 230296 30376
rect 229704 30336 229710 30348
rect 230290 30336 230296 30348
rect 230348 30336 230354 30388
rect 231302 30336 231308 30388
rect 231360 30376 231366 30388
rect 231762 30376 231768 30388
rect 231360 30348 231768 30376
rect 231360 30336 231366 30348
rect 231762 30336 231768 30348
rect 231820 30336 231826 30388
rect 232958 30336 232964 30388
rect 233016 30376 233022 30388
rect 233142 30376 233148 30388
rect 233016 30348 233148 30376
rect 233016 30336 233022 30348
rect 233142 30336 233148 30348
rect 233200 30336 233206 30388
rect 235166 30336 235172 30388
rect 235224 30376 235230 30388
rect 235810 30376 235816 30388
rect 235224 30348 235816 30376
rect 235224 30336 235230 30348
rect 235810 30336 235816 30348
rect 235868 30336 235874 30388
rect 239493 30379 239551 30385
rect 239493 30376 239505 30379
rect 235920 30348 239505 30376
rect 235718 30268 235724 30320
rect 235776 30308 235782 30320
rect 235920 30308 235948 30348
rect 239493 30345 239505 30348
rect 239539 30345 239551 30379
rect 239493 30339 239551 30345
rect 239582 30336 239588 30388
rect 239640 30376 239646 30388
rect 240042 30376 240048 30388
rect 239640 30348 240048 30376
rect 239640 30336 239646 30348
rect 240042 30336 240048 30348
rect 240100 30336 240106 30388
rect 240778 30336 240784 30388
rect 240836 30376 240842 30388
rect 241330 30376 241336 30388
rect 240836 30348 241336 30376
rect 240836 30336 240842 30348
rect 241330 30336 241336 30348
rect 241388 30336 241394 30388
rect 241882 30336 241888 30388
rect 241940 30376 241946 30388
rect 242710 30376 242716 30388
rect 241940 30348 242716 30376
rect 241940 30336 241946 30348
rect 242710 30336 242716 30348
rect 242768 30336 242774 30388
rect 243538 30336 243544 30388
rect 243596 30376 243602 30388
rect 244182 30376 244188 30388
rect 243596 30348 244188 30376
rect 243596 30336 243602 30348
rect 244182 30336 244188 30348
rect 244240 30336 244246 30388
rect 244642 30336 244648 30388
rect 244700 30376 244706 30388
rect 245562 30376 245568 30388
rect 244700 30348 245568 30376
rect 244700 30336 244706 30348
rect 245562 30336 245568 30348
rect 245620 30336 245626 30388
rect 246298 30336 246304 30388
rect 246356 30376 246362 30388
rect 246942 30376 246948 30388
rect 246356 30348 246948 30376
rect 246356 30336 246362 30348
rect 246942 30336 246948 30348
rect 247000 30336 247006 30388
rect 247402 30336 247408 30388
rect 247460 30376 247466 30388
rect 248138 30376 248144 30388
rect 247460 30348 248144 30376
rect 247460 30336 247466 30348
rect 248138 30336 248144 30348
rect 248196 30336 248202 30388
rect 248233 30379 248291 30385
rect 248233 30345 248245 30379
rect 248279 30376 248291 30379
rect 312538 30376 312544 30388
rect 248279 30348 312544 30376
rect 248279 30345 248291 30348
rect 248233 30339 248291 30345
rect 312538 30336 312544 30348
rect 312596 30336 312602 30388
rect 235776 30280 235948 30308
rect 235776 30268 235782 30280
rect 201402 30240 201408 30252
rect 201144 30212 201408 30240
rect 201402 30200 201408 30212
rect 201460 30200 201466 30252
rect 296622 30200 296628 30252
rect 296680 30200 296686 30252
rect 296530 29996 296536 30048
rect 296588 30036 296594 30048
rect 296640 30036 296668 30200
rect 296588 30008 296668 30036
rect 296588 29996 296594 30008
rect 258534 27276 258540 27328
rect 258592 27316 258598 27328
rect 259362 27316 259368 27328
rect 258592 27288 259368 27316
rect 258592 27276 258598 27288
rect 259362 27276 259368 27288
rect 259420 27276 259426 27328
rect 234430 16056 234436 16108
rect 234488 16096 234494 16108
rect 436738 16096 436744 16108
rect 234488 16068 436744 16096
rect 234488 16056 234494 16068
rect 436738 16056 436744 16068
rect 436796 16056 436802 16108
rect 241330 15988 241336 16040
rect 241388 16028 241394 16040
rect 450906 16028 450912 16040
rect 241388 16000 450912 16028
rect 241388 15988 241394 16000
rect 450906 15988 450912 16000
rect 450964 15988 450970 16040
rect 244090 15920 244096 15972
rect 244148 15960 244154 15972
rect 456794 15960 456800 15972
rect 244148 15932 456800 15960
rect 244148 15920 244154 15932
rect 456794 15920 456800 15932
rect 456852 15920 456858 15972
rect 248138 15852 248144 15904
rect 248196 15892 248202 15904
rect 465166 15892 465172 15904
rect 248196 15864 465172 15892
rect 248196 15852 248202 15864
rect 465166 15852 465172 15864
rect 465224 15852 465230 15904
rect 227438 15104 227444 15156
rect 227496 15144 227502 15156
rect 420914 15144 420920 15156
rect 227496 15116 420920 15144
rect 227496 15104 227502 15116
rect 420914 15104 420920 15116
rect 420972 15104 420978 15156
rect 229002 15036 229008 15088
rect 229060 15076 229066 15088
rect 423674 15076 423680 15088
rect 229060 15048 423680 15076
rect 229060 15036 229066 15048
rect 423674 15036 423680 15048
rect 423732 15036 423738 15088
rect 230198 14968 230204 15020
rect 230256 15008 230262 15020
rect 428458 15008 428464 15020
rect 230256 14980 428464 15008
rect 230256 14968 230262 14980
rect 428458 14968 428464 14980
rect 428516 14968 428522 15020
rect 231670 14900 231676 14952
rect 231728 14940 231734 14952
rect 432046 14940 432052 14952
rect 231728 14912 432052 14940
rect 231728 14900 231734 14912
rect 432046 14900 432052 14912
rect 432104 14900 432110 14952
rect 233050 14832 233056 14884
rect 233108 14872 233114 14884
rect 435082 14872 435088 14884
rect 233108 14844 435088 14872
rect 233108 14832 233114 14844
rect 435082 14832 435088 14844
rect 435140 14832 435146 14884
rect 248230 14764 248236 14816
rect 248288 14804 248294 14816
rect 465810 14804 465816 14816
rect 248288 14776 465816 14804
rect 248288 14764 248294 14776
rect 465810 14764 465816 14776
rect 465868 14764 465874 14816
rect 249702 14696 249708 14748
rect 249760 14736 249766 14748
rect 469858 14736 469864 14748
rect 249760 14708 469864 14736
rect 249760 14696 249766 14708
rect 469858 14696 469864 14708
rect 469916 14696 469922 14748
rect 253658 14628 253664 14680
rect 253716 14668 253722 14680
rect 476482 14668 476488 14680
rect 253716 14640 476488 14668
rect 253716 14628 253722 14640
rect 476482 14628 476488 14640
rect 476540 14628 476546 14680
rect 250898 14560 250904 14612
rect 250956 14600 250962 14612
rect 473446 14600 473452 14612
rect 250956 14572 473452 14600
rect 250956 14560 250962 14572
rect 473446 14560 473452 14572
rect 473504 14560 473510 14612
rect 290918 14492 290924 14544
rect 290976 14532 290982 14544
rect 556890 14532 556896 14544
rect 290976 14504 556896 14532
rect 290976 14492 290982 14504
rect 556890 14492 556896 14504
rect 556948 14492 556954 14544
rect 292390 14424 292396 14476
rect 292448 14464 292454 14476
rect 559282 14464 559288 14476
rect 292448 14436 559288 14464
rect 292448 14424 292454 14436
rect 559282 14424 559288 14436
rect 559340 14424 559346 14476
rect 208210 14356 208216 14408
rect 208268 14396 208274 14408
rect 381170 14396 381176 14408
rect 208268 14368 381176 14396
rect 208268 14356 208274 14368
rect 381170 14356 381176 14368
rect 381228 14356 381234 14408
rect 206738 14288 206744 14340
rect 206796 14328 206802 14340
rect 377674 14328 377680 14340
rect 206796 14300 377680 14328
rect 206796 14288 206802 14300
rect 377674 14288 377680 14300
rect 377732 14288 377738 14340
rect 187418 14220 187424 14272
rect 187476 14260 187482 14272
rect 336274 14260 336280 14272
rect 187476 14232 336280 14260
rect 187476 14220 187482 14232
rect 336274 14220 336280 14232
rect 336332 14220 336338 14272
rect 184658 14152 184664 14204
rect 184716 14192 184722 14204
rect 332686 14192 332692 14204
rect 184716 14164 332692 14192
rect 184716 14152 184722 14164
rect 332686 14152 332692 14164
rect 332744 14152 332750 14204
rect 183370 14084 183376 14136
rect 183428 14124 183434 14136
rect 328730 14124 328736 14136
rect 183428 14096 328736 14124
rect 183428 14084 183434 14096
rect 328730 14084 328736 14096
rect 328788 14084 328794 14136
rect 181990 14016 181996 14068
rect 182048 14056 182054 14068
rect 326338 14056 326344 14068
rect 182048 14028 326344 14056
rect 182048 14016 182054 14028
rect 326338 14016 326344 14028
rect 326396 14016 326402 14068
rect 181898 13948 181904 14000
rect 181956 13988 181962 14000
rect 324314 13988 324320 14000
rect 181956 13960 324320 13988
rect 181956 13948 181962 13960
rect 324314 13948 324320 13960
rect 324372 13948 324378 14000
rect 177850 13880 177856 13932
rect 177908 13920 177914 13932
rect 316034 13920 316040 13932
rect 177908 13892 316040 13920
rect 177908 13880 177914 13892
rect 316034 13880 316040 13892
rect 316092 13880 316098 13932
rect 173710 13812 173716 13864
rect 173768 13852 173774 13864
rect 307754 13852 307760 13864
rect 173768 13824 307760 13852
rect 173768 13812 173774 13824
rect 307754 13812 307760 13824
rect 307812 13812 307818 13864
rect 257890 13744 257896 13796
rect 257948 13784 257954 13796
rect 487154 13784 487160 13796
rect 257948 13756 487160 13784
rect 257948 13744 257954 13756
rect 487154 13744 487160 13756
rect 487212 13744 487218 13796
rect 259178 13676 259184 13728
rect 259236 13716 259242 13728
rect 489914 13716 489920 13728
rect 259236 13688 489920 13716
rect 259236 13676 259242 13688
rect 489914 13676 489920 13688
rect 489972 13676 489978 13728
rect 261938 13608 261944 13660
rect 261996 13648 262002 13660
rect 494698 13648 494704 13660
rect 261996 13620 494704 13648
rect 261996 13608 262002 13620
rect 494698 13608 494704 13620
rect 494756 13608 494762 13660
rect 275830 13540 275836 13592
rect 275888 13580 275894 13592
rect 525426 13580 525432 13592
rect 275888 13552 525432 13580
rect 275888 13540 275894 13552
rect 525426 13540 525432 13552
rect 525484 13540 525490 13592
rect 279878 13472 279884 13524
rect 279936 13512 279942 13524
rect 532050 13512 532056 13524
rect 279936 13484 532056 13512
rect 279936 13472 279942 13484
rect 532050 13472 532056 13484
rect 532108 13472 532114 13524
rect 158438 13404 158444 13456
rect 158496 13444 158502 13456
rect 274818 13444 274824 13456
rect 158496 13416 274824 13444
rect 158496 13404 158502 13416
rect 274818 13404 274824 13416
rect 274876 13404 274882 13456
rect 277118 13404 277124 13456
rect 277176 13444 277182 13456
rect 528554 13444 528560 13456
rect 277176 13416 528560 13444
rect 277176 13404 277182 13416
rect 528554 13404 528560 13416
rect 528612 13404 528618 13456
rect 159910 13336 159916 13388
rect 159968 13376 159974 13388
rect 278314 13376 278320 13388
rect 159968 13348 278320 13376
rect 159968 13336 159974 13348
rect 278314 13336 278320 13348
rect 278372 13336 278378 13388
rect 281350 13336 281356 13388
rect 281408 13376 281414 13388
rect 536098 13376 536104 13388
rect 281408 13348 536104 13376
rect 281408 13336 281414 13348
rect 536098 13336 536104 13348
rect 536156 13336 536162 13388
rect 162762 13268 162768 13320
rect 162820 13308 162826 13320
rect 284938 13308 284944 13320
rect 162820 13280 284944 13308
rect 162820 13268 162826 13280
rect 284938 13268 284944 13280
rect 284996 13268 285002 13320
rect 285398 13268 285404 13320
rect 285456 13308 285462 13320
rect 546678 13308 546684 13320
rect 285456 13280 546684 13308
rect 285456 13268 285462 13280
rect 546678 13268 546684 13280
rect 546736 13268 546742 13320
rect 163958 13200 163964 13252
rect 164016 13240 164022 13252
rect 288986 13240 288992 13252
rect 164016 13212 288992 13240
rect 164016 13200 164022 13212
rect 288986 13200 288992 13212
rect 289044 13200 289050 13252
rect 289630 13200 289636 13252
rect 289688 13240 289694 13252
rect 553762 13240 553768 13252
rect 289688 13212 553768 13240
rect 289688 13200 289694 13212
rect 553762 13200 553768 13212
rect 553820 13200 553826 13252
rect 169570 13132 169576 13184
rect 169628 13172 169634 13184
rect 299658 13172 299664 13184
rect 169628 13144 299664 13172
rect 169628 13132 169634 13144
rect 299658 13132 299664 13144
rect 299716 13132 299722 13184
rect 300670 13132 300676 13184
rect 300728 13172 300734 13184
rect 576946 13172 576952 13184
rect 300728 13144 576952 13172
rect 300728 13132 300734 13144
rect 576946 13132 576952 13144
rect 577004 13132 577010 13184
rect 171042 13064 171048 13116
rect 171100 13104 171106 13116
rect 303154 13104 303160 13116
rect 171100 13076 303160 13104
rect 171100 13064 171106 13076
rect 303154 13064 303160 13076
rect 303212 13064 303218 13116
rect 304258 13064 304264 13116
rect 304316 13104 304322 13116
rect 581730 13104 581736 13116
rect 304316 13076 581736 13104
rect 304316 13064 304322 13076
rect 581730 13064 581736 13076
rect 581788 13064 581794 13116
rect 256418 12996 256424 13048
rect 256476 13036 256482 13048
rect 484026 13036 484032 13048
rect 256476 13008 484032 13036
rect 256476 12996 256482 13008
rect 484026 12996 484032 13008
rect 484084 12996 484090 13048
rect 255130 12928 255136 12980
rect 255188 12968 255194 12980
rect 480530 12968 480536 12980
rect 255188 12940 480536 12968
rect 255188 12928 255194 12940
rect 480530 12928 480536 12940
rect 480588 12928 480594 12980
rect 203978 12860 203984 12912
rect 204036 12900 204042 12912
rect 374086 12900 374092 12912
rect 204036 12872 374092 12900
rect 204036 12860 204042 12872
rect 374086 12860 374092 12872
rect 374144 12860 374150 12912
rect 202782 12792 202788 12844
rect 202840 12832 202846 12844
rect 370130 12832 370136 12844
rect 202840 12804 370136 12832
rect 202840 12792 202846 12804
rect 370130 12792 370136 12804
rect 370188 12792 370194 12844
rect 177942 12724 177948 12776
rect 178000 12764 178006 12776
rect 317322 12764 317328 12776
rect 178000 12736 317328 12764
rect 178000 12724 178006 12736
rect 317322 12724 317328 12736
rect 317380 12724 317386 12776
rect 176470 12656 176476 12708
rect 176528 12696 176534 12708
rect 313826 12696 313832 12708
rect 176528 12668 313832 12696
rect 176528 12656 176534 12668
rect 313826 12656 313832 12668
rect 313884 12656 313890 12708
rect 172330 12588 172336 12640
rect 172388 12628 172394 12640
rect 306374 12628 306380 12640
rect 172388 12600 306380 12628
rect 172388 12588 172394 12600
rect 306374 12588 306380 12600
rect 306432 12588 306438 12640
rect 175090 12520 175096 12572
rect 175148 12560 175154 12572
rect 309686 12560 309692 12572
rect 175148 12532 309692 12560
rect 175148 12520 175154 12532
rect 309686 12520 309692 12532
rect 309744 12520 309750 12572
rect 168190 12452 168196 12504
rect 168248 12492 168254 12504
rect 295610 12492 295616 12504
rect 168248 12464 295616 12492
rect 168248 12452 168254 12464
rect 295610 12452 295616 12464
rect 295668 12452 295674 12504
rect 296438 12452 296444 12504
rect 296496 12492 296502 12504
rect 418798 12492 418804 12504
rect 296496 12464 418804 12492
rect 296496 12452 296502 12464
rect 418798 12452 418804 12464
rect 418856 12452 418862 12504
rect 250990 12384 250996 12436
rect 251048 12424 251054 12436
rect 470594 12424 470600 12436
rect 251048 12396 470600 12424
rect 251048 12384 251054 12396
rect 470594 12384 470600 12396
rect 470652 12384 470658 12436
rect 252462 12316 252468 12368
rect 252520 12356 252526 12368
rect 474090 12356 474096 12368
rect 252520 12328 474096 12356
rect 252520 12316 252526 12328
rect 474090 12316 474096 12328
rect 474148 12316 474154 12368
rect 253750 12248 253756 12300
rect 253808 12288 253814 12300
rect 478138 12288 478144 12300
rect 253808 12260 478144 12288
rect 253808 12248 253814 12260
rect 478138 12248 478144 12260
rect 478196 12248 478202 12300
rect 256510 12180 256516 12232
rect 256568 12220 256574 12232
rect 482370 12220 482376 12232
rect 256568 12192 482376 12220
rect 256568 12180 256574 12192
rect 482370 12180 482376 12192
rect 482428 12180 482434 12232
rect 257982 12112 257988 12164
rect 258040 12152 258046 12164
rect 486418 12152 486424 12164
rect 258040 12124 486424 12152
rect 258040 12112 258046 12124
rect 486418 12112 486424 12124
rect 486476 12112 486482 12164
rect 259270 12044 259276 12096
rect 259328 12084 259334 12096
rect 490006 12084 490012 12096
rect 259328 12056 490012 12084
rect 259328 12044 259334 12056
rect 490006 12044 490012 12056
rect 490064 12044 490070 12096
rect 260650 11976 260656 12028
rect 260708 12016 260714 12028
rect 493042 12016 493048 12028
rect 260708 11988 493048 12016
rect 260708 11976 260714 11988
rect 493042 11976 493048 11988
rect 493100 11976 493106 12028
rect 262030 11908 262036 11960
rect 262088 11948 262094 11960
rect 497090 11948 497096 11960
rect 262088 11920 497096 11948
rect 262088 11908 262094 11920
rect 497090 11908 497096 11920
rect 497148 11908 497154 11960
rect 264698 11840 264704 11892
rect 264756 11880 264762 11892
rect 500586 11880 500592 11892
rect 264756 11852 500592 11880
rect 264756 11840 264762 11852
rect 500586 11840 500592 11852
rect 500644 11840 500650 11892
rect 266170 11772 266176 11824
rect 266228 11812 266234 11824
rect 503714 11812 503720 11824
rect 266228 11784 503720 11812
rect 266228 11772 266234 11784
rect 503714 11772 503720 11784
rect 503772 11772 503778 11824
rect 267458 11704 267464 11756
rect 267516 11744 267522 11756
rect 507210 11744 507216 11756
rect 267516 11716 507216 11744
rect 267516 11704 267522 11716
rect 507210 11704 507216 11716
rect 507268 11704 507274 11756
rect 248322 11636 248328 11688
rect 248380 11676 248386 11688
rect 467466 11676 467472 11688
rect 248380 11648 467472 11676
rect 248380 11636 248386 11648
rect 467466 11636 467472 11648
rect 467524 11636 467530 11688
rect 246850 11568 246856 11620
rect 246908 11608 246914 11620
rect 463970 11608 463976 11620
rect 246908 11580 463976 11608
rect 246908 11568 246914 11580
rect 463970 11568 463976 11580
rect 464028 11568 464034 11620
rect 245470 11500 245476 11552
rect 245528 11540 245534 11552
rect 459922 11540 459928 11552
rect 245528 11512 459928 11540
rect 245528 11500 245534 11512
rect 459922 11500 459928 11512
rect 459980 11500 459986 11552
rect 244182 11432 244188 11484
rect 244240 11472 244246 11484
rect 456886 11472 456892 11484
rect 244240 11444 456892 11472
rect 244240 11432 244246 11444
rect 456886 11432 456892 11444
rect 456944 11432 456950 11484
rect 242710 11364 242716 11416
rect 242768 11404 242774 11416
rect 453298 11404 453304 11416
rect 242768 11376 453304 11404
rect 242768 11364 242774 11376
rect 453298 11364 453304 11376
rect 453356 11364 453362 11416
rect 239950 11296 239956 11348
rect 240008 11336 240014 11348
rect 448514 11336 448520 11348
rect 240008 11308 448520 11336
rect 240008 11296 240014 11308
rect 448514 11296 448520 11308
rect 448572 11296 448578 11348
rect 238570 11228 238576 11280
rect 238628 11268 238634 11280
rect 445754 11268 445760 11280
rect 238628 11240 445760 11268
rect 238628 11228 238634 11240
rect 445754 11228 445760 11240
rect 445812 11228 445818 11280
rect 235810 11160 235816 11212
rect 235868 11200 235874 11212
rect 439130 11200 439136 11212
rect 235868 11172 439136 11200
rect 235868 11160 235874 11172
rect 439130 11160 439136 11172
rect 439188 11160 439194 11212
rect 164050 11092 164056 11144
rect 164108 11132 164114 11144
rect 287330 11132 287336 11144
rect 164108 11104 287336 11132
rect 164108 11092 164114 11104
rect 287330 11092 287336 11104
rect 287388 11092 287394 11144
rect 201218 10956 201224 11008
rect 201276 10996 201282 11008
rect 367738 10996 367744 11008
rect 201276 10968 367744 10996
rect 201276 10956 201282 10968
rect 367738 10956 367744 10968
rect 367796 10956 367802 11008
rect 204070 10888 204076 10940
rect 204128 10928 204134 10940
rect 371234 10928 371240 10940
rect 204128 10900 371240 10928
rect 204128 10888 204134 10900
rect 371234 10888 371240 10900
rect 371292 10888 371298 10940
rect 205542 10820 205548 10872
rect 205600 10860 205606 10872
rect 375282 10860 375288 10872
rect 205600 10832 375288 10860
rect 205600 10820 205606 10832
rect 375282 10820 375288 10832
rect 375340 10820 375346 10872
rect 206830 10752 206836 10804
rect 206888 10792 206894 10804
rect 378410 10792 378416 10804
rect 206888 10764 378416 10792
rect 206888 10752 206894 10764
rect 378410 10752 378416 10764
rect 378468 10752 378474 10804
rect 208302 10684 208308 10736
rect 208360 10724 208366 10736
rect 382366 10724 382372 10736
rect 208360 10696 382372 10724
rect 208360 10684 208366 10696
rect 382366 10684 382372 10696
rect 382424 10684 382430 10736
rect 210878 10616 210884 10668
rect 210936 10656 210942 10668
rect 385954 10656 385960 10668
rect 210936 10628 385960 10656
rect 210936 10616 210942 10628
rect 385954 10616 385960 10628
rect 386012 10616 386018 10668
rect 212442 10548 212448 10600
rect 212500 10588 212506 10600
rect 389450 10588 389456 10600
rect 212500 10560 389456 10588
rect 212500 10548 212506 10560
rect 389450 10548 389456 10560
rect 389508 10548 389514 10600
rect 213638 10480 213644 10532
rect 213696 10520 213702 10532
rect 392578 10520 392584 10532
rect 213696 10492 392584 10520
rect 213696 10480 213702 10492
rect 392578 10480 392584 10492
rect 392636 10480 392642 10532
rect 215110 10412 215116 10464
rect 215168 10452 215174 10464
rect 396074 10452 396080 10464
rect 215168 10424 396080 10452
rect 215168 10412 215174 10424
rect 396074 10412 396080 10424
rect 396132 10412 396138 10464
rect 216490 10344 216496 10396
rect 216548 10384 216554 10396
rect 398834 10384 398840 10396
rect 216548 10356 398840 10384
rect 216548 10344 216554 10356
rect 398834 10344 398840 10356
rect 398892 10344 398898 10396
rect 219250 10276 219256 10328
rect 219308 10316 219314 10328
rect 403618 10316 403624 10328
rect 219308 10288 403624 10316
rect 219308 10276 219314 10288
rect 403618 10276 403624 10288
rect 403676 10276 403682 10328
rect 199930 10208 199936 10260
rect 199988 10248 199994 10260
rect 364610 10248 364616 10260
rect 199988 10220 364616 10248
rect 199988 10208 199994 10220
rect 364610 10208 364616 10220
rect 364668 10208 364674 10260
rect 198550 10140 198556 10192
rect 198608 10180 198614 10192
rect 361114 10180 361120 10192
rect 198608 10152 361120 10180
rect 198608 10140 198614 10152
rect 361114 10140 361120 10152
rect 361172 10140 361178 10192
rect 197170 10072 197176 10124
rect 197228 10112 197234 10124
rect 357526 10112 357532 10124
rect 197228 10084 357532 10112
rect 197228 10072 197234 10084
rect 357526 10072 357532 10084
rect 357584 10072 357590 10124
rect 195790 10004 195796 10056
rect 195848 10044 195854 10056
rect 353570 10044 353576 10056
rect 195848 10016 353576 10044
rect 195848 10004 195854 10016
rect 353570 10004 353576 10016
rect 353628 10004 353634 10056
rect 193030 9936 193036 9988
rect 193088 9976 193094 9988
rect 349154 9976 349160 9988
rect 193088 9948 349160 9976
rect 193088 9936 193094 9948
rect 349154 9936 349160 9948
rect 349212 9936 349218 9988
rect 191650 9868 191656 9920
rect 191708 9908 191714 9920
rect 346946 9908 346952 9920
rect 191708 9880 346952 9908
rect 191708 9868 191714 9880
rect 346946 9868 346952 9880
rect 347004 9868 347010 9920
rect 190178 9800 190184 9852
rect 190236 9840 190242 9852
rect 342898 9840 342904 9852
rect 190236 9812 342904 9840
rect 190236 9800 190242 9812
rect 342898 9800 342904 9812
rect 342956 9800 342962 9852
rect 188982 9732 188988 9784
rect 189040 9772 189046 9784
rect 339494 9772 339500 9784
rect 189040 9744 339500 9772
rect 189040 9732 189046 9744
rect 339494 9732 339500 9744
rect 339552 9732 339558 9784
rect 244918 9664 244924 9716
rect 244976 9704 244982 9716
rect 305546 9704 305552 9716
rect 244976 9676 305552 9704
rect 244976 9664 244982 9676
rect 305546 9664 305552 9676
rect 305604 9664 305610 9716
rect 157150 9596 157156 9648
rect 157208 9636 157214 9648
rect 273622 9636 273628 9648
rect 157208 9608 273628 9636
rect 157208 9596 157214 9608
rect 273622 9596 273628 9608
rect 273680 9596 273686 9648
rect 274450 9596 274456 9648
rect 274508 9636 274514 9648
rect 520734 9636 520740 9648
rect 274508 9608 520740 9636
rect 274508 9596 274514 9608
rect 520734 9596 520740 9608
rect 520792 9596 520798 9648
rect 158530 9528 158536 9580
rect 158588 9568 158594 9580
rect 277118 9568 277124 9580
rect 158588 9540 277124 9568
rect 158588 9528 158594 9540
rect 277118 9528 277124 9540
rect 277176 9528 277182 9580
rect 277210 9528 277216 9580
rect 277268 9568 277274 9580
rect 527818 9568 527824 9580
rect 277268 9540 527824 9568
rect 277268 9528 277274 9540
rect 527818 9528 527824 9540
rect 527876 9528 527882 9580
rect 160002 9460 160008 9512
rect 160060 9500 160066 9512
rect 279510 9500 279516 9512
rect 160060 9472 279516 9500
rect 160060 9460 160066 9472
rect 279510 9460 279516 9472
rect 279568 9460 279574 9512
rect 279970 9460 279976 9512
rect 280028 9500 280034 9512
rect 280028 9472 280844 9500
rect 280028 9460 280034 9472
rect 161198 9392 161204 9444
rect 161256 9432 161262 9444
rect 280706 9432 280712 9444
rect 161256 9404 280712 9432
rect 161256 9392 161262 9404
rect 280706 9392 280712 9404
rect 280764 9392 280770 9444
rect 280816 9432 280844 9472
rect 282730 9460 282736 9512
rect 282788 9500 282794 9512
rect 286873 9503 286931 9509
rect 282788 9472 286824 9500
rect 282788 9460 282794 9472
rect 280816 9404 283328 9432
rect 164142 9324 164148 9376
rect 164200 9364 164206 9376
rect 283193 9367 283251 9373
rect 283193 9364 283205 9367
rect 164200 9336 283205 9364
rect 164200 9324 164206 9336
rect 283193 9333 283205 9336
rect 283239 9333 283251 9367
rect 283193 9327 283251 9333
rect 161290 9256 161296 9308
rect 161348 9296 161354 9308
rect 283098 9296 283104 9308
rect 161348 9268 283104 9296
rect 161348 9256 161354 9268
rect 283098 9256 283104 9268
rect 283156 9256 283162 9308
rect 283300 9296 283328 9404
rect 284202 9392 284208 9444
rect 284260 9432 284266 9444
rect 286796 9432 286824 9472
rect 286873 9469 286885 9503
rect 286919 9500 286931 9503
rect 534902 9500 534908 9512
rect 286919 9472 534908 9500
rect 286919 9469 286931 9472
rect 286873 9463 286931 9469
rect 534902 9460 534908 9472
rect 534960 9460 534966 9512
rect 538398 9432 538404 9444
rect 284260 9404 286732 9432
rect 286796 9404 538404 9432
rect 284260 9392 284266 9404
rect 283377 9367 283435 9373
rect 283377 9333 283389 9367
rect 283423 9364 283435 9367
rect 286594 9364 286600 9376
rect 283423 9336 286600 9364
rect 283423 9333 283435 9336
rect 283377 9327 283435 9333
rect 286594 9324 286600 9336
rect 286652 9324 286658 9376
rect 286704 9364 286732 9404
rect 538398 9392 538404 9404
rect 538456 9392 538462 9444
rect 541986 9364 541992 9376
rect 286704 9336 541992 9364
rect 541986 9324 541992 9336
rect 542044 9324 542050 9376
rect 286781 9299 286839 9305
rect 286781 9296 286793 9299
rect 283300 9268 286793 9296
rect 286781 9265 286793 9268
rect 286827 9265 286839 9299
rect 286781 9259 286839 9265
rect 286870 9256 286876 9308
rect 286928 9296 286934 9308
rect 549070 9296 549076 9308
rect 286928 9268 549076 9296
rect 286928 9256 286934 9268
rect 549070 9256 549076 9268
rect 549128 9256 549134 9308
rect 165522 9188 165528 9240
rect 165580 9228 165586 9240
rect 290182 9228 290188 9240
rect 165580 9200 290188 9228
rect 165580 9188 165586 9200
rect 290182 9188 290188 9200
rect 290240 9188 290246 9240
rect 293770 9188 293776 9240
rect 293828 9228 293834 9240
rect 563238 9228 563244 9240
rect 293828 9200 563244 9228
rect 293828 9188 293834 9200
rect 563238 9188 563244 9200
rect 563296 9188 563302 9240
rect 166810 9120 166816 9172
rect 166868 9160 166874 9172
rect 293678 9160 293684 9172
rect 166868 9132 293684 9160
rect 166868 9120 166874 9132
rect 293678 9120 293684 9132
rect 293736 9120 293742 9172
rect 295150 9120 295156 9172
rect 295208 9160 295214 9172
rect 566826 9160 566832 9172
rect 295208 9132 566832 9160
rect 295208 9120 295214 9132
rect 566826 9120 566832 9132
rect 566884 9120 566890 9172
rect 173802 9052 173808 9104
rect 173860 9092 173866 9104
rect 307938 9092 307944 9104
rect 173860 9064 307944 9092
rect 173860 9052 173866 9064
rect 307938 9052 307944 9064
rect 307996 9052 308002 9104
rect 308398 9052 308404 9104
rect 308456 9092 308462 9104
rect 580994 9092 581000 9104
rect 308456 9064 581000 9092
rect 308456 9052 308462 9064
rect 580994 9052 581000 9064
rect 581052 9052 581058 9104
rect 168282 8984 168288 9036
rect 168340 9024 168346 9036
rect 297266 9024 297272 9036
rect 168340 8996 297272 9024
rect 168340 8984 168346 8996
rect 297266 8984 297272 8996
rect 297324 8984 297330 9036
rect 299290 8984 299296 9036
rect 299348 9024 299354 9036
rect 300581 9027 300639 9033
rect 300581 9024 300593 9027
rect 299348 8996 300593 9024
rect 299348 8984 299354 8996
rect 300581 8993 300593 8996
rect 300627 8993 300639 9027
rect 300581 8987 300639 8993
rect 300670 8984 300676 9036
rect 300728 9024 300734 9036
rect 300949 9027 301007 9033
rect 300728 8996 300900 9024
rect 300728 8984 300734 8996
rect 169662 8916 169668 8968
rect 169720 8956 169726 8968
rect 300762 8956 300768 8968
rect 169720 8928 300768 8956
rect 169720 8916 169726 8928
rect 300762 8916 300768 8928
rect 300820 8916 300826 8968
rect 300872 8956 300900 8996
rect 300949 8993 300961 9027
rect 300995 9024 301007 9027
rect 573910 9024 573916 9036
rect 300995 8996 573916 9024
rect 300995 8993 301007 8996
rect 300949 8987 301007 8993
rect 573910 8984 573916 8996
rect 573968 8984 573974 9036
rect 578602 8956 578608 8968
rect 300872 8928 578608 8956
rect 578602 8916 578608 8928
rect 578660 8916 578666 8968
rect 155678 8848 155684 8900
rect 155736 8888 155742 8900
rect 270034 8888 270040 8900
rect 155736 8860 270040 8888
rect 155736 8848 155742 8860
rect 270034 8848 270040 8860
rect 270092 8848 270098 8900
rect 270310 8848 270316 8900
rect 270368 8888 270374 8900
rect 513558 8888 513564 8900
rect 270368 8860 513564 8888
rect 270368 8848 270374 8860
rect 513558 8848 513564 8860
rect 513616 8848 513622 8900
rect 154390 8780 154396 8832
rect 154448 8820 154454 8832
rect 266538 8820 266544 8832
rect 154448 8792 266544 8820
rect 154448 8780 154454 8792
rect 266538 8780 266544 8792
rect 266596 8780 266602 8832
rect 267550 8780 267556 8832
rect 267608 8820 267614 8832
rect 506474 8820 506480 8832
rect 267608 8792 506480 8820
rect 267608 8780 267614 8792
rect 506474 8780 506480 8792
rect 506532 8780 506538 8832
rect 152918 8712 152924 8764
rect 152976 8752 152982 8764
rect 262950 8752 262956 8764
rect 152976 8724 262956 8752
rect 152976 8712 152982 8724
rect 262950 8712 262956 8724
rect 263008 8712 263014 8764
rect 263410 8712 263416 8764
rect 263468 8752 263474 8764
rect 499390 8752 499396 8764
rect 263468 8724 499396 8752
rect 263468 8712 263474 8724
rect 499390 8712 499396 8724
rect 499448 8712 499454 8764
rect 150158 8644 150164 8696
rect 150216 8684 150222 8696
rect 259454 8684 259460 8696
rect 150216 8656 259460 8684
rect 150216 8644 150222 8656
rect 259454 8644 259460 8656
rect 259512 8644 259518 8696
rect 262122 8644 262128 8696
rect 262180 8684 262186 8696
rect 495894 8684 495900 8696
rect 262180 8656 495900 8684
rect 262180 8644 262186 8656
rect 495894 8644 495900 8656
rect 495952 8644 495958 8696
rect 148870 8576 148876 8628
rect 148928 8616 148934 8628
rect 255866 8616 255872 8628
rect 148928 8588 255872 8616
rect 148928 8576 148934 8588
rect 255866 8576 255872 8588
rect 255924 8576 255930 8628
rect 259362 8576 259368 8628
rect 259420 8616 259426 8628
rect 488810 8616 488816 8628
rect 259420 8588 488816 8616
rect 259420 8576 259426 8588
rect 488810 8576 488816 8588
rect 488868 8576 488874 8628
rect 147398 8508 147404 8560
rect 147456 8548 147462 8560
rect 252370 8548 252376 8560
rect 147456 8520 252376 8548
rect 147456 8508 147462 8520
rect 252370 8508 252376 8520
rect 252428 8508 252434 8560
rect 256602 8508 256608 8560
rect 256660 8548 256666 8560
rect 485222 8548 485228 8560
rect 256660 8520 485228 8548
rect 256660 8508 256666 8520
rect 485222 8508 485228 8520
rect 485280 8508 485286 8560
rect 146110 8440 146116 8492
rect 146168 8480 146174 8492
rect 248782 8480 248788 8492
rect 146168 8452 248788 8480
rect 146168 8440 146174 8452
rect 248782 8440 248788 8452
rect 248840 8440 248846 8492
rect 255222 8440 255228 8492
rect 255280 8480 255286 8492
rect 481726 8480 481732 8492
rect 255280 8452 481732 8480
rect 255280 8440 255286 8452
rect 481726 8440 481732 8452
rect 481784 8440 481790 8492
rect 175182 8372 175188 8424
rect 175240 8412 175246 8424
rect 311434 8412 311440 8424
rect 175240 8384 311440 8412
rect 175240 8372 175246 8384
rect 311434 8372 311440 8384
rect 311492 8372 311498 8424
rect 172422 8304 172428 8356
rect 172480 8344 172486 8356
rect 304350 8344 304356 8356
rect 172480 8316 304356 8344
rect 172480 8304 172486 8316
rect 304350 8304 304356 8316
rect 304408 8304 304414 8356
rect 223482 8236 223488 8288
rect 223540 8276 223546 8288
rect 413094 8276 413100 8288
rect 223540 8248 413100 8276
rect 223540 8236 223546 8248
rect 413094 8236 413100 8248
rect 413152 8236 413158 8288
rect 123938 8168 123944 8220
rect 123996 8208 124002 8220
rect 201494 8208 201500 8220
rect 123996 8180 201500 8208
rect 123996 8168 124002 8180
rect 201494 8168 201500 8180
rect 201552 8168 201558 8220
rect 224770 8168 224776 8220
rect 224828 8208 224834 8220
rect 416682 8208 416688 8220
rect 224828 8180 416688 8208
rect 224828 8168 224834 8180
rect 416682 8168 416688 8180
rect 416740 8168 416746 8220
rect 125410 8100 125416 8152
rect 125468 8140 125474 8152
rect 205082 8140 205088 8152
rect 125468 8112 205088 8140
rect 125468 8100 125474 8112
rect 205082 8100 205088 8112
rect 205140 8100 205146 8152
rect 226242 8100 226248 8152
rect 226300 8140 226306 8152
rect 420178 8140 420184 8152
rect 226300 8112 420184 8140
rect 226300 8100 226306 8112
rect 420178 8100 420184 8112
rect 420236 8100 420242 8152
rect 126698 8032 126704 8084
rect 126756 8072 126762 8084
rect 208578 8072 208584 8084
rect 126756 8044 208584 8072
rect 126756 8032 126762 8044
rect 208578 8032 208584 8044
rect 208636 8032 208642 8084
rect 230290 8032 230296 8084
rect 230348 8072 230354 8084
rect 427262 8072 427268 8084
rect 230348 8044 427268 8072
rect 230348 8032 230354 8044
rect 427262 8032 427268 8044
rect 427320 8032 427326 8084
rect 132218 7964 132224 8016
rect 132276 8004 132282 8016
rect 219250 8004 219256 8016
rect 132276 7976 219256 8004
rect 132276 7964 132282 7976
rect 219250 7964 219256 7976
rect 219308 7964 219314 8016
rect 227530 7964 227536 8016
rect 227588 8004 227594 8016
rect 423766 8004 423772 8016
rect 227588 7976 423772 8004
rect 227588 7964 227594 7976
rect 423766 7964 423772 7976
rect 423824 7964 423830 8016
rect 129458 7896 129464 7948
rect 129516 7936 129522 7948
rect 215662 7936 215668 7948
rect 129516 7908 215668 7936
rect 129516 7896 129522 7908
rect 215662 7896 215668 7908
rect 215720 7896 215726 7948
rect 231762 7896 231768 7948
rect 231820 7936 231826 7948
rect 430850 7936 430856 7948
rect 231820 7908 430856 7936
rect 231820 7896 231826 7908
rect 430850 7896 430856 7908
rect 430908 7896 430914 7948
rect 133690 7828 133696 7880
rect 133748 7868 133754 7880
rect 222746 7868 222752 7880
rect 133748 7840 222752 7868
rect 133748 7828 133754 7840
rect 222746 7828 222752 7840
rect 222804 7828 222810 7880
rect 233142 7828 233148 7880
rect 233200 7868 233206 7880
rect 434438 7868 434444 7880
rect 233200 7840 434444 7868
rect 233200 7828 233206 7840
rect 434438 7828 434444 7840
rect 434496 7828 434502 7880
rect 134978 7760 134984 7812
rect 135036 7800 135042 7812
rect 226334 7800 226340 7812
rect 135036 7772 226340 7800
rect 135036 7760 135042 7772
rect 226334 7760 226340 7772
rect 226392 7760 226398 7812
rect 234522 7760 234528 7812
rect 234580 7800 234586 7812
rect 437934 7800 437940 7812
rect 234580 7772 437940 7800
rect 234580 7760 234586 7772
rect 437934 7760 437940 7772
rect 437992 7760 437998 7812
rect 139210 7692 139216 7744
rect 139268 7732 139274 7744
rect 234614 7732 234620 7744
rect 139268 7704 234620 7732
rect 139268 7692 139274 7704
rect 234614 7692 234620 7704
rect 234672 7692 234678 7744
rect 235902 7692 235908 7744
rect 235960 7732 235966 7744
rect 441522 7732 441528 7744
rect 235960 7704 441528 7732
rect 235960 7692 235966 7704
rect 441522 7692 441528 7704
rect 441580 7692 441586 7744
rect 141970 7624 141976 7676
rect 142028 7664 142034 7676
rect 241698 7664 241704 7676
rect 142028 7636 241704 7664
rect 142028 7624 142034 7636
rect 241698 7624 241704 7636
rect 241756 7624 241762 7676
rect 242802 7624 242808 7676
rect 242860 7664 242866 7676
rect 455690 7664 455696 7676
rect 242860 7636 455696 7664
rect 242860 7624 242866 7636
rect 455690 7624 455696 7636
rect 455748 7624 455754 7676
rect 143258 7556 143264 7608
rect 143316 7596 143322 7608
rect 245194 7596 245200 7608
rect 143316 7568 245200 7596
rect 143316 7556 143322 7568
rect 245194 7556 245200 7568
rect 245252 7556 245258 7608
rect 245562 7556 245568 7608
rect 245620 7596 245626 7608
rect 459186 7596 459192 7608
rect 245620 7568 459192 7596
rect 245620 7556 245626 7568
rect 459186 7556 459192 7568
rect 459244 7556 459250 7608
rect 219342 7488 219348 7540
rect 219400 7528 219406 7540
rect 406010 7528 406016 7540
rect 219400 7500 406016 7528
rect 219400 7488 219406 7500
rect 406010 7488 406016 7500
rect 406068 7488 406074 7540
rect 222102 7420 222108 7472
rect 222160 7460 222166 7472
rect 409598 7460 409604 7472
rect 222160 7432 409604 7460
rect 222160 7420 222166 7432
rect 409598 7420 409604 7432
rect 409656 7420 409662 7472
rect 217870 7352 217876 7404
rect 217928 7392 217934 7404
rect 402514 7392 402520 7404
rect 217928 7364 402520 7392
rect 217928 7352 217934 7364
rect 402514 7352 402520 7364
rect 402572 7352 402578 7404
rect 216582 7284 216588 7336
rect 216640 7324 216646 7336
rect 398926 7324 398932 7336
rect 216640 7296 398932 7324
rect 216640 7284 216646 7296
rect 398926 7284 398932 7296
rect 398984 7284 398990 7336
rect 215202 7216 215208 7268
rect 215260 7256 215266 7268
rect 395338 7256 395344 7268
rect 215260 7228 395344 7256
rect 215260 7216 215266 7228
rect 395338 7216 395344 7228
rect 395396 7216 395402 7268
rect 213730 7148 213736 7200
rect 213788 7188 213794 7200
rect 391842 7188 391848 7200
rect 213788 7160 391848 7188
rect 213788 7148 213794 7160
rect 391842 7148 391848 7160
rect 391900 7148 391906 7200
rect 210970 7080 210976 7132
rect 211028 7120 211034 7132
rect 388254 7120 388260 7132
rect 211028 7092 388260 7120
rect 211028 7080 211034 7092
rect 388254 7080 388260 7092
rect 388312 7080 388318 7132
rect 209682 7012 209688 7064
rect 209740 7052 209746 7064
rect 384758 7052 384764 7064
rect 209740 7024 384764 7052
rect 209740 7012 209746 7024
rect 384758 7012 384764 7024
rect 384816 7012 384822 7064
rect 158622 6944 158628 6996
rect 158680 6984 158686 6996
rect 276014 6984 276020 6996
rect 158680 6956 276020 6984
rect 158680 6944 158686 6956
rect 276014 6944 276020 6956
rect 276072 6944 276078 6996
rect 276658 6944 276664 6996
rect 276716 6984 276722 6996
rect 319714 6984 319720 6996
rect 276716 6956 319720 6984
rect 276716 6944 276722 6956
rect 319714 6944 319720 6956
rect 319772 6944 319778 6996
rect 142062 6808 142068 6860
rect 142120 6848 142126 6860
rect 240502 6848 240508 6860
rect 142120 6820 240508 6848
rect 142120 6808 142126 6820
rect 240502 6808 240508 6820
rect 240560 6808 240566 6860
rect 242158 6808 242164 6860
rect 242216 6848 242222 6860
rect 301406 6848 301412 6860
rect 242216 6820 301412 6848
rect 242216 6808 242222 6820
rect 301406 6808 301412 6820
rect 301464 6808 301470 6860
rect 301498 6808 301504 6860
rect 301556 6848 301562 6860
rect 312630 6848 312636 6860
rect 301556 6820 312636 6848
rect 301556 6808 301562 6820
rect 312630 6808 312636 6820
rect 312688 6808 312694 6860
rect 315298 6808 315304 6860
rect 315356 6848 315362 6860
rect 580166 6848 580172 6860
rect 315356 6820 580172 6848
rect 315356 6808 315362 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 117130 6740 117136 6792
rect 117188 6780 117194 6792
rect 187326 6780 187332 6792
rect 117188 6752 187332 6780
rect 117188 6740 117194 6752
rect 187326 6740 187332 6752
rect 187384 6740 187390 6792
rect 198642 6740 198648 6792
rect 198700 6780 198706 6792
rect 359918 6780 359924 6792
rect 198700 6752 359924 6780
rect 198700 6740 198706 6752
rect 359918 6740 359924 6752
rect 359976 6740 359982 6792
rect 118510 6672 118516 6724
rect 118568 6712 118574 6724
rect 190822 6712 190828 6724
rect 118568 6684 190828 6712
rect 118568 6672 118574 6684
rect 190822 6672 190828 6684
rect 190880 6672 190886 6724
rect 200022 6672 200028 6724
rect 200080 6712 200086 6724
rect 363506 6712 363512 6724
rect 200080 6684 363512 6712
rect 200080 6672 200086 6684
rect 363506 6672 363512 6684
rect 363564 6672 363570 6724
rect 119982 6604 119988 6656
rect 120040 6644 120046 6656
rect 194318 6644 194324 6656
rect 120040 6616 194324 6644
rect 120040 6604 120046 6616
rect 194318 6604 194324 6616
rect 194376 6604 194382 6656
rect 201310 6604 201316 6656
rect 201368 6644 201374 6656
rect 367002 6644 367008 6656
rect 201368 6616 367008 6644
rect 201368 6604 201374 6616
rect 367002 6604 367008 6616
rect 367060 6604 367066 6656
rect 121270 6536 121276 6588
rect 121328 6576 121334 6588
rect 197906 6576 197912 6588
rect 121328 6548 197912 6576
rect 121328 6536 121334 6548
rect 197906 6536 197912 6548
rect 197964 6536 197970 6588
rect 237190 6536 237196 6588
rect 237248 6576 237254 6588
rect 442626 6576 442632 6588
rect 237248 6548 442632 6576
rect 237248 6536 237254 6548
rect 442626 6536 442632 6548
rect 442684 6536 442690 6588
rect 143350 6468 143356 6520
rect 143408 6508 143414 6520
rect 244090 6508 244096 6520
rect 143408 6480 244096 6508
rect 143408 6468 143414 6480
rect 244090 6468 244096 6480
rect 244148 6468 244154 6520
rect 260742 6468 260748 6520
rect 260800 6508 260806 6520
rect 492306 6508 492312 6520
rect 260800 6480 492312 6508
rect 260800 6468 260806 6480
rect 492306 6468 492312 6480
rect 492364 6468 492370 6520
rect 144730 6400 144736 6452
rect 144788 6440 144794 6452
rect 247586 6440 247592 6452
rect 144788 6412 247592 6440
rect 144788 6400 144794 6412
rect 247586 6400 247592 6412
rect 247644 6400 247650 6452
rect 264790 6400 264796 6452
rect 264848 6440 264854 6452
rect 502978 6440 502984 6452
rect 264848 6412 502984 6440
rect 264848 6400 264854 6412
rect 502978 6400 502984 6412
rect 503036 6400 503042 6452
rect 147490 6332 147496 6384
rect 147548 6372 147554 6384
rect 251174 6372 251180 6384
rect 147548 6344 251180 6372
rect 147548 6332 147554 6344
rect 251174 6332 251180 6344
rect 251232 6332 251238 6384
rect 269022 6332 269028 6384
rect 269080 6372 269086 6384
rect 510062 6372 510068 6384
rect 269080 6344 510068 6372
rect 269080 6332 269086 6344
rect 510062 6332 510068 6344
rect 510120 6332 510126 6384
rect 99190 6264 99196 6316
rect 99248 6304 99254 6316
rect 150618 6304 150624 6316
rect 99248 6276 150624 6304
rect 99248 6264 99254 6276
rect 150618 6264 150624 6276
rect 150676 6264 150682 6316
rect 151630 6264 151636 6316
rect 151688 6304 151694 6316
rect 261754 6304 261760 6316
rect 151688 6276 261760 6304
rect 151688 6264 151694 6276
rect 261754 6264 261760 6276
rect 261812 6264 261818 6316
rect 271690 6264 271696 6316
rect 271748 6304 271754 6316
rect 517146 6304 517152 6316
rect 271748 6276 517152 6304
rect 271748 6264 271754 6276
rect 517146 6264 517152 6276
rect 517204 6264 517210 6316
rect 100478 6196 100484 6248
rect 100536 6236 100542 6248
rect 154206 6236 154212 6248
rect 100536 6208 154212 6236
rect 100536 6196 100542 6208
rect 154206 6196 154212 6208
rect 154264 6196 154270 6248
rect 155770 6196 155776 6248
rect 155828 6236 155834 6248
rect 268838 6236 268844 6248
rect 155828 6208 268844 6236
rect 155828 6196 155834 6208
rect 268838 6196 268844 6208
rect 268896 6196 268902 6248
rect 275922 6196 275928 6248
rect 275980 6236 275986 6248
rect 524230 6236 524236 6248
rect 275980 6208 524236 6236
rect 275980 6196 275986 6208
rect 524230 6196 524236 6208
rect 524288 6196 524294 6248
rect 111610 6128 111616 6180
rect 111668 6168 111674 6180
rect 176654 6168 176660 6180
rect 111668 6140 176660 6168
rect 111668 6128 111674 6140
rect 176654 6128 176660 6140
rect 176712 6128 176718 6180
rect 179322 6128 179328 6180
rect 179380 6168 179386 6180
rect 320910 6168 320916 6180
rect 179380 6140 320916 6168
rect 179380 6128 179386 6140
rect 320910 6128 320916 6140
rect 320968 6128 320974 6180
rect 322198 6128 322204 6180
rect 322256 6168 322262 6180
rect 583389 6171 583447 6177
rect 583389 6168 583401 6171
rect 322256 6140 583401 6168
rect 322256 6128 322262 6140
rect 583389 6137 583401 6140
rect 583435 6137 583447 6171
rect 583389 6131 583447 6137
rect 115750 6060 115756 6112
rect 115808 6100 115814 6112
rect 183738 6100 183744 6112
rect 115808 6072 183744 6100
rect 115808 6060 115814 6072
rect 183738 6060 183744 6072
rect 183796 6060 183802 6112
rect 194410 6060 194416 6112
rect 194468 6100 194474 6112
rect 352834 6100 352840 6112
rect 194468 6072 352840 6100
rect 194468 6060 194474 6072
rect 352834 6060 352840 6072
rect 352892 6060 352898 6112
rect 114462 5992 114468 6044
rect 114520 6032 114526 6044
rect 181438 6032 181444 6044
rect 114520 6004 181444 6032
rect 114520 5992 114526 6004
rect 181438 5992 181444 6004
rect 181496 5992 181502 6044
rect 193122 5992 193128 6044
rect 193180 6032 193186 6044
rect 349246 6032 349252 6044
rect 193180 6004 349252 6032
rect 193180 5992 193186 6004
rect 349246 5992 349252 6004
rect 349304 5992 349310 6044
rect 113082 5924 113088 5976
rect 113140 5964 113146 5976
rect 180242 5964 180248 5976
rect 113140 5936 180248 5964
rect 113140 5924 113146 5936
rect 180242 5924 180248 5936
rect 180300 5924 180306 5976
rect 191742 5924 191748 5976
rect 191800 5964 191806 5976
rect 345750 5964 345756 5976
rect 191800 5936 345756 5964
rect 191800 5924 191806 5936
rect 345750 5924 345756 5936
rect 345808 5924 345814 5976
rect 110230 5856 110236 5908
rect 110288 5896 110294 5908
rect 173158 5896 173164 5908
rect 110288 5868 173164 5896
rect 110288 5856 110294 5868
rect 173158 5856 173164 5868
rect 173216 5856 173222 5908
rect 190270 5856 190276 5908
rect 190328 5896 190334 5908
rect 342162 5896 342168 5908
rect 190328 5868 342168 5896
rect 190328 5856 190334 5868
rect 342162 5856 342168 5868
rect 342220 5856 342226 5908
rect 108850 5788 108856 5840
rect 108908 5828 108914 5840
rect 170766 5828 170772 5840
rect 108908 5800 170772 5828
rect 108908 5788 108914 5800
rect 170766 5788 170772 5800
rect 170824 5788 170830 5840
rect 187510 5788 187516 5840
rect 187568 5828 187574 5840
rect 338666 5828 338672 5840
rect 187568 5800 338672 5828
rect 187568 5788 187574 5800
rect 338666 5788 338672 5800
rect 338724 5788 338730 5840
rect 106090 5720 106096 5772
rect 106148 5760 106154 5772
rect 166074 5760 166080 5772
rect 106148 5732 166080 5760
rect 106148 5720 106154 5732
rect 166074 5720 166080 5732
rect 166132 5720 166138 5772
rect 186222 5720 186228 5772
rect 186280 5760 186286 5772
rect 335078 5760 335084 5772
rect 186280 5732 335084 5760
rect 186280 5720 186286 5732
rect 335078 5720 335084 5732
rect 335136 5720 335142 5772
rect 108942 5652 108948 5704
rect 109000 5692 109006 5704
rect 169570 5692 169576 5704
rect 109000 5664 169576 5692
rect 109000 5652 109006 5664
rect 169570 5652 169576 5664
rect 169628 5652 169634 5704
rect 184750 5652 184756 5704
rect 184808 5692 184814 5704
rect 331582 5692 331588 5704
rect 184808 5664 331588 5692
rect 184808 5652 184814 5664
rect 331582 5652 331588 5664
rect 331640 5652 331646 5704
rect 104802 5584 104808 5636
rect 104860 5624 104866 5636
rect 162486 5624 162492 5636
rect 104860 5596 162492 5624
rect 104860 5584 104866 5596
rect 162486 5584 162492 5596
rect 162544 5584 162550 5636
rect 183462 5584 183468 5636
rect 183520 5624 183526 5636
rect 327994 5624 328000 5636
rect 183520 5596 328000 5624
rect 183520 5584 183526 5596
rect 327994 5584 328000 5596
rect 328052 5584 328058 5636
rect 103238 5516 103244 5568
rect 103296 5556 103302 5568
rect 157794 5556 157800 5568
rect 103296 5528 157800 5556
rect 103296 5516 103302 5528
rect 157794 5516 157800 5528
rect 157852 5516 157858 5568
rect 182082 5516 182088 5568
rect 182140 5556 182146 5568
rect 324406 5556 324412 5568
rect 182140 5528 324412 5556
rect 182140 5516 182146 5528
rect 324406 5516 324412 5528
rect 324464 5516 324470 5568
rect 93762 5448 93768 5500
rect 93820 5488 93826 5500
rect 137646 5488 137652 5500
rect 93820 5460 137652 5488
rect 93820 5448 93826 5460
rect 137646 5448 137652 5460
rect 137704 5448 137710 5500
rect 137830 5448 137836 5500
rect 137888 5488 137894 5500
rect 232222 5488 232228 5500
rect 137888 5460 232228 5488
rect 137888 5448 137894 5460
rect 232222 5448 232228 5460
rect 232280 5448 232286 5500
rect 278682 5448 278688 5500
rect 278740 5488 278746 5500
rect 530118 5488 530124 5500
rect 278740 5460 530124 5488
rect 278740 5448 278746 5460
rect 530118 5448 530124 5460
rect 530176 5448 530182 5500
rect 94958 5380 94964 5432
rect 95016 5420 95022 5432
rect 140038 5420 140044 5432
rect 95016 5392 140044 5420
rect 95016 5380 95022 5392
rect 140038 5380 140044 5392
rect 140096 5380 140102 5432
rect 140590 5380 140596 5432
rect 140648 5420 140654 5432
rect 239306 5420 239312 5432
rect 140648 5392 239312 5420
rect 140648 5380 140654 5392
rect 239306 5380 239312 5392
rect 239364 5380 239370 5432
rect 280062 5380 280068 5432
rect 280120 5420 280126 5432
rect 533706 5420 533712 5432
rect 280120 5392 533712 5420
rect 280120 5380 280126 5392
rect 533706 5380 533712 5392
rect 533764 5380 533770 5432
rect 95050 5312 95056 5364
rect 95108 5352 95114 5364
rect 141234 5352 141240 5364
rect 95108 5324 141240 5352
rect 95108 5312 95114 5324
rect 141234 5312 141240 5324
rect 141292 5312 141298 5364
rect 143442 5312 143448 5364
rect 143500 5352 143506 5364
rect 242894 5352 242900 5364
rect 143500 5324 242900 5352
rect 143500 5312 143506 5324
rect 242894 5312 242900 5324
rect 242952 5312 242958 5364
rect 281442 5312 281448 5364
rect 281500 5352 281506 5364
rect 537202 5352 537208 5364
rect 281500 5324 537208 5352
rect 281500 5312 281506 5324
rect 537202 5312 537208 5324
rect 537260 5312 537266 5364
rect 96522 5244 96528 5296
rect 96580 5284 96586 5296
rect 143534 5284 143540 5296
rect 96580 5256 143540 5284
rect 96580 5244 96586 5256
rect 143534 5244 143540 5256
rect 143592 5244 143598 5296
rect 144822 5244 144828 5296
rect 144880 5284 144886 5296
rect 246390 5284 246396 5296
rect 144880 5256 246396 5284
rect 144880 5244 144886 5256
rect 246390 5244 246396 5256
rect 246448 5244 246454 5296
rect 282822 5244 282828 5296
rect 282880 5284 282886 5296
rect 540790 5284 540796 5296
rect 282880 5256 540796 5284
rect 282880 5244 282886 5256
rect 540790 5244 540796 5256
rect 540848 5244 540854 5296
rect 96430 5176 96436 5228
rect 96488 5216 96494 5228
rect 144730 5216 144736 5228
rect 96488 5188 144736 5216
rect 96488 5176 96494 5188
rect 144730 5176 144736 5188
rect 144788 5176 144794 5228
rect 146202 5176 146208 5228
rect 146260 5216 146266 5228
rect 249978 5216 249984 5228
rect 146260 5188 249984 5216
rect 146260 5176 146266 5188
rect 249978 5176 249984 5188
rect 250036 5176 250042 5228
rect 281905 5219 281963 5225
rect 281905 5185 281917 5219
rect 281951 5216 281963 5219
rect 284294 5216 284300 5228
rect 281951 5188 284300 5216
rect 281951 5185 281963 5188
rect 281905 5179 281963 5185
rect 284294 5176 284300 5188
rect 284352 5176 284358 5228
rect 285582 5176 285588 5228
rect 285640 5216 285646 5228
rect 544378 5216 544384 5228
rect 285640 5188 544384 5216
rect 285640 5176 285646 5188
rect 544378 5176 544384 5188
rect 544436 5176 544442 5228
rect 97810 5108 97816 5160
rect 97868 5148 97874 5160
rect 147122 5148 147128 5160
rect 97868 5120 147128 5148
rect 97868 5108 97874 5120
rect 147122 5108 147128 5120
rect 147180 5108 147186 5160
rect 147582 5108 147588 5160
rect 147640 5148 147646 5160
rect 253474 5148 253480 5160
rect 147640 5120 253480 5148
rect 147640 5108 147646 5120
rect 253474 5108 253480 5120
rect 253532 5108 253538 5160
rect 273162 5108 273168 5160
rect 273220 5148 273226 5160
rect 282549 5151 282607 5157
rect 282549 5148 282561 5151
rect 273220 5120 282561 5148
rect 273220 5108 273226 5120
rect 282549 5117 282561 5120
rect 282595 5117 282607 5151
rect 282549 5111 282607 5117
rect 286962 5108 286968 5160
rect 287020 5148 287026 5160
rect 547874 5148 547880 5160
rect 287020 5120 547880 5148
rect 287020 5108 287026 5120
rect 547874 5108 547880 5120
rect 547932 5108 547938 5160
rect 97718 5040 97724 5092
rect 97776 5080 97782 5092
rect 148318 5080 148324 5092
rect 97776 5052 148324 5080
rect 97776 5040 97782 5052
rect 148318 5040 148324 5052
rect 148376 5040 148382 5092
rect 150342 5040 150348 5092
rect 150400 5080 150406 5092
rect 257062 5080 257068 5092
rect 150400 5052 257068 5080
rect 150400 5040 150406 5052
rect 257062 5040 257068 5052
rect 257120 5040 257126 5092
rect 271782 5040 271788 5092
rect 271840 5080 271846 5092
rect 282457 5083 282515 5089
rect 282457 5080 282469 5083
rect 271840 5052 282469 5080
rect 271840 5040 271846 5052
rect 282457 5049 282469 5052
rect 282503 5049 282515 5083
rect 282457 5043 282515 5049
rect 288342 5040 288348 5092
rect 288400 5080 288406 5092
rect 551462 5080 551468 5092
rect 288400 5052 551468 5080
rect 288400 5040 288406 5052
rect 551462 5040 551468 5052
rect 551520 5040 551526 5092
rect 100570 4972 100576 5024
rect 100628 5012 100634 5024
rect 151814 5012 151820 5024
rect 100628 4984 151820 5012
rect 100628 4972 100634 4984
rect 151814 4972 151820 4984
rect 151872 4972 151878 5024
rect 153102 4972 153108 5024
rect 153160 5012 153166 5024
rect 264146 5012 264152 5024
rect 153160 4984 264152 5012
rect 153160 4972 153166 4984
rect 264146 4972 264152 4984
rect 264204 4972 264210 5024
rect 270402 4972 270408 5024
rect 270460 5012 270466 5024
rect 272889 5015 272947 5021
rect 272889 5012 272901 5015
rect 270460 4984 272901 5012
rect 270460 4972 270466 4984
rect 272889 4981 272901 4984
rect 272935 4981 272947 5015
rect 272889 4975 272947 4981
rect 274542 4972 274548 5024
rect 274600 5012 274606 5024
rect 282270 5012 282276 5024
rect 274600 4984 282276 5012
rect 274600 4972 274606 4984
rect 282270 4972 282276 4984
rect 282328 4972 282334 5024
rect 282365 5015 282423 5021
rect 282365 4981 282377 5015
rect 282411 5012 282423 5015
rect 298462 5012 298468 5024
rect 282411 4984 298468 5012
rect 282411 4981 282423 4984
rect 282365 4975 282423 4981
rect 298462 4972 298468 4984
rect 298520 4972 298526 5024
rect 299382 4972 299388 5024
rect 299440 5012 299446 5024
rect 301409 5015 301467 5021
rect 301409 5012 301421 5015
rect 299440 4984 301421 5012
rect 299440 4972 299446 4984
rect 301409 4981 301421 4984
rect 301455 4981 301467 5015
rect 301409 4975 301467 4981
rect 301501 5015 301559 5021
rect 301501 4981 301513 5015
rect 301547 5012 301559 5015
rect 562042 5012 562048 5024
rect 301547 4984 562048 5012
rect 301547 4981 301559 4984
rect 301501 4975 301559 4981
rect 562042 4972 562048 4984
rect 562100 4972 562106 5024
rect 102042 4904 102048 4956
rect 102100 4944 102106 4956
rect 155402 4944 155408 4956
rect 102100 4916 155408 4944
rect 102100 4904 102106 4916
rect 155402 4904 155408 4916
rect 155460 4904 155466 4956
rect 155862 4904 155868 4956
rect 155920 4944 155926 4956
rect 271230 4944 271236 4956
rect 155920 4916 271236 4944
rect 155920 4904 155926 4916
rect 271230 4904 271236 4916
rect 271288 4904 271294 4956
rect 277302 4904 277308 4956
rect 277360 4944 277366 4956
rect 281997 4947 282055 4953
rect 281997 4944 282009 4947
rect 277360 4916 282009 4944
rect 277360 4904 277366 4916
rect 281997 4913 282009 4916
rect 282043 4913 282055 4947
rect 281997 4907 282055 4913
rect 282086 4904 282092 4956
rect 282144 4944 282150 4956
rect 294874 4944 294880 4956
rect 282144 4916 294880 4944
rect 282144 4904 282150 4916
rect 294874 4904 294880 4916
rect 294932 4904 294938 4956
rect 295242 4904 295248 4956
rect 295300 4944 295306 4956
rect 565630 4944 565636 4956
rect 295300 4916 565636 4944
rect 295300 4904 295306 4916
rect 565630 4904 565636 4916
rect 565688 4904 565694 4956
rect 103330 4836 103336 4888
rect 103388 4876 103394 4888
rect 158898 4876 158904 4888
rect 103388 4848 158904 4876
rect 103388 4836 103394 4848
rect 158898 4836 158904 4848
rect 158956 4836 158962 4888
rect 161382 4836 161388 4888
rect 161440 4876 161446 4888
rect 281902 4876 281908 4888
rect 161440 4848 281908 4876
rect 161440 4836 161446 4848
rect 281902 4836 281908 4848
rect 281960 4836 281966 4888
rect 282181 4879 282239 4885
rect 282181 4845 282193 4879
rect 282227 4876 282239 4879
rect 291378 4876 291384 4888
rect 282227 4848 291384 4876
rect 282227 4845 282239 4848
rect 282181 4839 282239 4845
rect 291378 4836 291384 4848
rect 291436 4836 291442 4888
rect 296622 4836 296628 4888
rect 296680 4876 296686 4888
rect 569126 4876 569132 4888
rect 296680 4848 569132 4876
rect 296680 4836 296686 4848
rect 569126 4836 569132 4848
rect 569184 4836 569190 4888
rect 106182 4768 106188 4820
rect 106240 4808 106246 4820
rect 163682 4808 163688 4820
rect 106240 4780 163688 4808
rect 106240 4768 106246 4780
rect 163682 4768 163688 4780
rect 163740 4768 163746 4820
rect 166902 4768 166908 4820
rect 166960 4808 166966 4820
rect 292574 4808 292580 4820
rect 166960 4780 281948 4808
rect 166960 4768 166966 4780
rect 92290 4700 92296 4752
rect 92348 4740 92354 4752
rect 134150 4740 134156 4752
rect 92348 4712 134156 4740
rect 92348 4700 92354 4712
rect 134150 4700 134156 4712
rect 134208 4700 134214 4752
rect 136542 4700 136548 4752
rect 136600 4740 136606 4752
rect 228726 4740 228732 4752
rect 136600 4712 228732 4740
rect 136600 4700 136606 4712
rect 228726 4700 228732 4712
rect 228784 4700 228790 4752
rect 272429 4743 272487 4749
rect 272429 4709 272441 4743
rect 272475 4740 272487 4743
rect 281810 4740 281816 4752
rect 272475 4712 281816 4740
rect 272475 4709 272487 4712
rect 272429 4703 272487 4709
rect 281810 4700 281816 4712
rect 281868 4700 281874 4752
rect 281920 4740 281948 4780
rect 282288 4780 292580 4808
rect 282288 4740 282316 4780
rect 292574 4768 292580 4780
rect 292632 4768 292638 4820
rect 293862 4768 293868 4820
rect 293920 4808 293926 4820
rect 301501 4811 301559 4817
rect 301501 4808 301513 4811
rect 293920 4780 301513 4808
rect 293920 4768 293926 4780
rect 301501 4777 301513 4780
rect 301547 4777 301559 4811
rect 301501 4771 301559 4777
rect 301593 4811 301651 4817
rect 301593 4777 301605 4811
rect 301639 4808 301651 4811
rect 576302 4808 576308 4820
rect 301639 4780 576308 4808
rect 301639 4777 301651 4780
rect 301593 4771 301651 4777
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 281920 4712 282316 4740
rect 282362 4700 282368 4752
rect 282420 4740 282426 4752
rect 523034 4740 523040 4752
rect 282420 4712 523040 4740
rect 282420 4700 282426 4712
rect 523034 4700 523040 4712
rect 523092 4700 523098 4752
rect 89622 4632 89628 4684
rect 89680 4672 89686 4684
rect 129366 4672 129372 4684
rect 89680 4644 129372 4672
rect 89680 4632 89686 4644
rect 129366 4632 129372 4644
rect 129424 4632 129430 4684
rect 135070 4632 135076 4684
rect 135128 4672 135134 4684
rect 225138 4672 225144 4684
rect 135128 4644 225144 4672
rect 135128 4632 135134 4644
rect 225138 4632 225144 4644
rect 225196 4632 225202 4684
rect 263502 4632 263508 4684
rect 263560 4672 263566 4684
rect 272337 4675 272395 4681
rect 272337 4672 272349 4675
rect 263560 4644 272349 4672
rect 263560 4632 263566 4644
rect 272337 4641 272349 4644
rect 272383 4641 272395 4675
rect 272337 4635 272395 4641
rect 272521 4675 272579 4681
rect 272521 4641 272533 4675
rect 272567 4672 272579 4675
rect 282181 4675 282239 4681
rect 282181 4672 282193 4675
rect 272567 4644 282193 4672
rect 272567 4641 272579 4644
rect 272521 4635 272579 4641
rect 282181 4641 282193 4644
rect 282227 4641 282239 4675
rect 526622 4672 526628 4684
rect 282181 4635 282239 4641
rect 282288 4644 526628 4672
rect 88242 4564 88248 4616
rect 88300 4604 88306 4616
rect 125870 4604 125876 4616
rect 88300 4576 125876 4604
rect 88300 4564 88306 4576
rect 125870 4564 125876 4576
rect 125928 4564 125934 4616
rect 132310 4564 132316 4616
rect 132368 4604 132374 4616
rect 221550 4604 221556 4616
rect 132368 4576 221556 4604
rect 132368 4564 132374 4576
rect 221550 4564 221556 4576
rect 221608 4564 221614 4616
rect 264882 4564 264888 4616
rect 264940 4604 264946 4616
rect 272705 4607 272763 4613
rect 272705 4604 272717 4607
rect 264940 4576 272717 4604
rect 264940 4564 264946 4576
rect 272705 4573 272717 4576
rect 272751 4573 272763 4607
rect 272705 4567 272763 4573
rect 272797 4607 272855 4613
rect 272797 4573 272809 4607
rect 272843 4604 272855 4607
rect 281905 4607 281963 4613
rect 281905 4604 281917 4607
rect 272843 4576 281917 4604
rect 272843 4573 272855 4576
rect 272797 4567 272855 4573
rect 281905 4573 281917 4576
rect 281951 4573 281963 4607
rect 281905 4567 281963 4573
rect 281997 4607 282055 4613
rect 281997 4573 282009 4607
rect 282043 4604 282055 4607
rect 282288 4604 282316 4644
rect 526622 4632 526628 4644
rect 526680 4632 526686 4684
rect 282043 4576 282316 4604
rect 282549 4607 282607 4613
rect 282043 4573 282055 4576
rect 281997 4567 282055 4573
rect 282549 4573 282561 4607
rect 282595 4604 282607 4607
rect 519538 4604 519544 4616
rect 282595 4576 519544 4604
rect 282595 4573 282607 4576
rect 282549 4567 282607 4573
rect 519538 4564 519544 4576
rect 519596 4564 519602 4616
rect 130930 4496 130936 4548
rect 130988 4536 130994 4548
rect 218054 4536 218060 4548
rect 130988 4508 218060 4536
rect 130988 4496 130994 4508
rect 218054 4496 218060 4508
rect 218112 4496 218118 4548
rect 218149 4539 218207 4545
rect 218149 4505 218161 4539
rect 218195 4536 218207 4539
rect 282365 4539 282423 4545
rect 282365 4536 282377 4539
rect 218195 4508 282377 4536
rect 218195 4505 218207 4508
rect 218149 4499 218207 4505
rect 282365 4505 282377 4508
rect 282411 4505 282423 4539
rect 282365 4499 282423 4505
rect 282457 4539 282515 4545
rect 282457 4505 282469 4539
rect 282503 4536 282515 4539
rect 515950 4536 515956 4548
rect 282503 4508 515956 4536
rect 282503 4505 282515 4508
rect 282457 4499 282515 4505
rect 515950 4496 515956 4508
rect 516008 4496 516014 4548
rect 124030 4428 124036 4480
rect 124088 4468 124094 4480
rect 203886 4468 203892 4480
rect 124088 4440 203892 4468
rect 124088 4428 124094 4440
rect 203886 4428 203892 4440
rect 203944 4428 203950 4480
rect 204898 4428 204904 4480
rect 204956 4468 204962 4480
rect 272521 4471 272579 4477
rect 272521 4468 272533 4471
rect 204956 4440 272533 4468
rect 204956 4428 204962 4440
rect 272521 4437 272533 4440
rect 272567 4437 272579 4471
rect 272521 4431 272579 4437
rect 272613 4471 272671 4477
rect 272613 4437 272625 4471
rect 272659 4468 272671 4471
rect 272797 4471 272855 4477
rect 272797 4468 272809 4471
rect 272659 4440 272809 4468
rect 272659 4437 272671 4440
rect 272613 4431 272671 4437
rect 272797 4437 272809 4440
rect 272843 4437 272855 4471
rect 272797 4431 272855 4437
rect 272889 4471 272947 4477
rect 272889 4437 272901 4471
rect 272935 4468 272947 4471
rect 512454 4468 512460 4480
rect 272935 4440 512460 4468
rect 272935 4437 272947 4440
rect 272889 4431 272947 4437
rect 512454 4428 512460 4440
rect 512512 4428 512518 4480
rect 126790 4360 126796 4412
rect 126848 4400 126854 4412
rect 207382 4400 207388 4412
rect 126848 4372 207388 4400
rect 126848 4360 126854 4372
rect 207382 4360 207388 4372
rect 207440 4360 207446 4412
rect 209038 4360 209044 4412
rect 209096 4400 209102 4412
rect 272429 4403 272487 4409
rect 272429 4400 272441 4403
rect 209096 4372 272441 4400
rect 209096 4360 209102 4372
rect 272429 4369 272441 4372
rect 272475 4369 272487 4403
rect 508866 4400 508872 4412
rect 272429 4363 272487 4369
rect 272536 4372 508872 4400
rect 129550 4292 129556 4344
rect 129608 4332 129614 4344
rect 214466 4332 214472 4344
rect 129608 4304 214472 4332
rect 129608 4292 129614 4304
rect 214466 4292 214472 4304
rect 214524 4292 214530 4344
rect 267642 4292 267648 4344
rect 267700 4332 267706 4344
rect 272536 4332 272564 4372
rect 508866 4360 508872 4372
rect 508924 4360 508930 4412
rect 505370 4332 505376 4344
rect 267700 4304 272564 4332
rect 272628 4304 505376 4332
rect 267700 4292 267706 4304
rect 122650 4224 122656 4276
rect 122708 4264 122714 4276
rect 200298 4264 200304 4276
rect 122708 4236 200304 4264
rect 122708 4224 122714 4236
rect 200298 4224 200304 4236
rect 200356 4224 200362 4276
rect 200758 4224 200764 4276
rect 200816 4264 200822 4276
rect 272521 4267 272579 4273
rect 272521 4264 272533 4267
rect 200816 4236 272533 4264
rect 200816 4224 200822 4236
rect 272521 4233 272533 4236
rect 272567 4233 272579 4267
rect 272521 4227 272579 4233
rect 103885 4199 103943 4205
rect 103885 4165 103897 4199
rect 103931 4196 103943 4199
rect 111521 4199 111579 4205
rect 103931 4168 104664 4196
rect 103931 4165 103943 4168
rect 103885 4159 103943 4165
rect 55030 4088 55036 4140
rect 55088 4128 55094 4140
rect 56042 4128 56048 4140
rect 55088 4100 56048 4128
rect 55088 4088 55094 4100
rect 56042 4088 56048 4100
rect 56100 4088 56106 4140
rect 64690 4088 64696 4140
rect 64748 4128 64754 4140
rect 76190 4128 76196 4140
rect 64748 4100 76196 4128
rect 64748 4088 64754 4100
rect 76190 4088 76196 4100
rect 76248 4088 76254 4140
rect 77110 4088 77116 4140
rect 77168 4128 77174 4140
rect 104526 4128 104532 4140
rect 77168 4100 104532 4128
rect 77168 4088 77174 4100
rect 104526 4088 104532 4100
rect 104584 4088 104590 4140
rect 104636 4128 104664 4168
rect 111521 4165 111533 4199
rect 111567 4196 111579 4199
rect 111567 4168 112944 4196
rect 111567 4165 111579 4168
rect 111521 4159 111579 4165
rect 112806 4128 112812 4140
rect 104636 4100 112812 4128
rect 112806 4088 112812 4100
rect 112864 4088 112870 4140
rect 112916 4128 112944 4168
rect 117222 4156 117228 4208
rect 117280 4196 117286 4208
rect 118053 4199 118111 4205
rect 118053 4196 118065 4199
rect 117280 4168 118065 4196
rect 117280 4156 117286 4168
rect 118053 4165 118065 4168
rect 118099 4165 118111 4199
rect 118053 4159 118111 4165
rect 128262 4156 128268 4208
rect 128320 4196 128326 4208
rect 210970 4196 210976 4208
rect 128320 4168 210976 4196
rect 128320 4156 128326 4168
rect 210970 4156 210976 4168
rect 211028 4156 211034 4208
rect 213178 4156 213184 4208
rect 213236 4196 213242 4208
rect 218149 4199 218207 4205
rect 218149 4196 218161 4199
rect 213236 4168 218161 4196
rect 213236 4156 213242 4168
rect 218149 4165 218161 4168
rect 218195 4165 218207 4199
rect 218149 4159 218207 4165
rect 266262 4156 266268 4208
rect 266320 4196 266326 4208
rect 272628 4196 272656 4304
rect 505370 4292 505376 4304
rect 505428 4292 505434 4344
rect 272705 4267 272763 4273
rect 272705 4233 272717 4267
rect 272751 4264 272763 4267
rect 501782 4264 501788 4276
rect 272751 4236 501788 4264
rect 272751 4233 272763 4236
rect 272705 4227 272763 4233
rect 501782 4224 501788 4236
rect 501840 4224 501846 4276
rect 266320 4168 272656 4196
rect 272797 4199 272855 4205
rect 266320 4156 266326 4168
rect 272797 4165 272809 4199
rect 272843 4196 272855 4199
rect 498194 4196 498200 4208
rect 272843 4168 498200 4196
rect 272843 4165 272855 4168
rect 272797 4159 272855 4165
rect 498194 4156 498200 4168
rect 498252 4156 498258 4208
rect 119890 4128 119896 4140
rect 112916 4100 119896 4128
rect 119890 4088 119896 4100
rect 119948 4088 119954 4140
rect 184934 4128 184940 4140
rect 120000 4100 184940 4128
rect 55122 4020 55128 4072
rect 55180 4060 55186 4072
rect 57238 4060 57244 4072
rect 55180 4032 57244 4060
rect 55180 4020 55186 4032
rect 57238 4020 57244 4032
rect 57296 4020 57302 4072
rect 63310 4020 63316 4072
rect 63368 4060 63374 4072
rect 74994 4060 75000 4072
rect 63368 4032 75000 4060
rect 63368 4020 63374 4032
rect 74994 4020 75000 4032
rect 75052 4020 75058 4072
rect 79870 4020 79876 4072
rect 79928 4060 79934 4072
rect 108114 4060 108120 4072
rect 79928 4032 108120 4060
rect 79928 4020 79934 4032
rect 108114 4020 108120 4032
rect 108172 4020 108178 4072
rect 108209 4063 108267 4069
rect 108209 4029 108221 4063
rect 108255 4060 108267 4063
rect 108255 4032 109448 4060
rect 108255 4029 108267 4032
rect 108209 4023 108267 4029
rect 64782 3952 64788 4004
rect 64840 3992 64846 4004
rect 77386 3992 77392 4004
rect 64840 3964 77392 3992
rect 64840 3952 64846 3964
rect 77386 3952 77392 3964
rect 77444 3952 77450 4004
rect 79962 3952 79968 4004
rect 80020 3992 80026 4004
rect 109310 3992 109316 4004
rect 80020 3964 109316 3992
rect 80020 3952 80026 3964
rect 109310 3952 109316 3964
rect 109368 3952 109374 4004
rect 109420 3992 109448 4032
rect 110322 4020 110328 4072
rect 110380 4060 110386 4072
rect 111797 4063 111855 4069
rect 111797 4060 111809 4063
rect 110380 4032 111809 4060
rect 110380 4020 110386 4032
rect 111797 4029 111809 4032
rect 111843 4029 111855 4063
rect 111797 4023 111855 4029
rect 111889 4063 111947 4069
rect 111889 4029 111901 4063
rect 111935 4060 111947 4063
rect 114002 4060 114008 4072
rect 111935 4032 114008 4060
rect 111935 4029 111947 4032
rect 111889 4023 111947 4029
rect 114002 4020 114008 4032
rect 114060 4020 114066 4072
rect 115842 4020 115848 4072
rect 115900 4060 115906 4072
rect 120000 4060 120028 4100
rect 184934 4088 184940 4100
rect 184992 4088 184998 4140
rect 185578 4088 185584 4140
rect 185636 4128 185642 4140
rect 196897 4131 196955 4137
rect 196897 4128 196909 4131
rect 185636 4100 196909 4128
rect 185636 4088 185642 4100
rect 196897 4097 196909 4100
rect 196943 4097 196955 4131
rect 196897 4091 196955 4097
rect 201402 4088 201408 4140
rect 201460 4128 201466 4140
rect 365806 4128 365812 4140
rect 201460 4100 365812 4128
rect 201460 4088 201466 4100
rect 365806 4088 365812 4100
rect 365864 4088 365870 4140
rect 366358 4088 366364 4140
rect 366416 4128 366422 4140
rect 368845 4131 368903 4137
rect 368845 4128 368857 4131
rect 366416 4100 368857 4128
rect 366416 4088 366422 4100
rect 368845 4097 368857 4100
rect 368891 4097 368903 4131
rect 368845 4091 368903 4097
rect 368937 4131 368995 4137
rect 368937 4097 368949 4131
rect 368983 4128 368995 4131
rect 373077 4131 373135 4137
rect 368983 4100 373028 4128
rect 368983 4097 368995 4100
rect 368937 4091 368995 4097
rect 115900 4032 120028 4060
rect 115900 4020 115906 4032
rect 121362 4020 121368 4072
rect 121420 4060 121426 4072
rect 127713 4063 127771 4069
rect 121420 4032 127664 4060
rect 121420 4020 121426 4032
rect 111521 3995 111579 4001
rect 111521 3992 111533 3995
rect 109420 3964 111533 3992
rect 111521 3961 111533 3964
rect 111567 3961 111579 3995
rect 111521 3955 111579 3961
rect 111705 3995 111763 4001
rect 111705 3961 111717 3995
rect 111751 3992 111763 3995
rect 118053 3995 118111 4001
rect 111751 3964 118004 3992
rect 111751 3961 111763 3964
rect 111705 3955 111763 3961
rect 26237 3927 26295 3933
rect 26237 3893 26249 3927
rect 26283 3924 26295 3927
rect 33318 3924 33324 3936
rect 26283 3896 33324 3924
rect 26283 3893 26295 3896
rect 26237 3887 26295 3893
rect 33318 3884 33324 3896
rect 33376 3884 33382 3936
rect 59170 3884 59176 3936
rect 59228 3924 59234 3936
rect 65518 3924 65524 3936
rect 59228 3896 65524 3924
rect 59228 3884 59234 3896
rect 65518 3884 65524 3896
rect 65576 3884 65582 3936
rect 66070 3884 66076 3936
rect 66128 3924 66134 3936
rect 79686 3924 79692 3936
rect 66128 3896 79692 3924
rect 66128 3884 66134 3896
rect 79686 3884 79692 3896
rect 79744 3884 79750 3936
rect 81250 3884 81256 3936
rect 81308 3924 81314 3936
rect 111610 3924 111616 3936
rect 81308 3896 111616 3924
rect 81308 3884 81314 3896
rect 111610 3884 111616 3896
rect 111668 3884 111674 3936
rect 111797 3927 111855 3933
rect 111797 3893 111809 3927
rect 111843 3924 111855 3927
rect 117869 3927 117927 3933
rect 117869 3924 117881 3927
rect 111843 3896 117881 3924
rect 111843 3893 111855 3896
rect 111797 3887 111855 3893
rect 117869 3893 117881 3896
rect 117915 3893 117927 3927
rect 117976 3924 118004 3964
rect 118053 3961 118065 3995
rect 118099 3992 118111 3995
rect 121181 3995 121239 4001
rect 121181 3992 121193 3995
rect 118099 3964 121193 3992
rect 118099 3961 118111 3964
rect 118053 3955 118111 3961
rect 121181 3961 121193 3964
rect 121227 3961 121239 3995
rect 121181 3955 121239 3961
rect 122742 3952 122748 4004
rect 122800 3992 122806 4004
rect 127529 3995 127587 4001
rect 127529 3992 127541 3995
rect 122800 3964 127541 3992
rect 122800 3952 122806 3964
rect 127529 3961 127541 3964
rect 127575 3961 127587 3995
rect 127636 3992 127664 4032
rect 127713 4029 127725 4063
rect 127759 4060 127771 4063
rect 188522 4060 188528 4072
rect 127759 4032 188528 4060
rect 127759 4029 127771 4032
rect 127713 4023 127771 4029
rect 188522 4020 188528 4032
rect 188580 4020 188586 4072
rect 204162 4020 204168 4072
rect 204220 4060 204226 4072
rect 372890 4060 372896 4072
rect 204220 4032 372896 4060
rect 204220 4020 204226 4032
rect 372890 4020 372896 4032
rect 372948 4020 372954 4072
rect 373000 4060 373028 4100
rect 373077 4097 373089 4131
rect 373123 4128 373135 4131
rect 383470 4128 383476 4140
rect 373123 4100 383476 4128
rect 373123 4097 373135 4100
rect 373077 4091 373135 4097
rect 383470 4088 383476 4100
rect 383528 4088 383534 4140
rect 383565 4131 383623 4137
rect 383565 4097 383577 4131
rect 383611 4128 383623 4131
rect 433242 4128 433248 4140
rect 383611 4100 433248 4128
rect 383611 4097 383623 4100
rect 383565 4091 383623 4097
rect 433242 4088 433248 4100
rect 433300 4088 433306 4140
rect 376478 4060 376484 4072
rect 373000 4032 376484 4060
rect 376478 4020 376484 4032
rect 376536 4020 376542 4072
rect 376570 4020 376576 4072
rect 376628 4060 376634 4072
rect 376628 4032 380112 4060
rect 376628 4020 376634 4032
rect 195606 3992 195612 4004
rect 127636 3964 195612 3992
rect 127529 3955 127587 3961
rect 195606 3952 195612 3964
rect 195664 3952 195670 4004
rect 200117 3995 200175 4001
rect 200117 3961 200129 3995
rect 200163 3992 200175 3995
rect 206186 3992 206192 4004
rect 200163 3964 206192 3992
rect 200163 3961 200175 3964
rect 200117 3955 200175 3961
rect 206186 3952 206192 3964
rect 206244 3952 206250 4004
rect 206922 3952 206928 4004
rect 206980 3992 206986 4004
rect 379974 3992 379980 4004
rect 206980 3964 379980 3992
rect 206980 3952 206986 3964
rect 379974 3952 379980 3964
rect 380032 3952 380038 4004
rect 380084 3992 380112 4032
rect 380158 4020 380164 4072
rect 380216 4060 380222 4072
rect 383381 4063 383439 4069
rect 383381 4060 383393 4063
rect 380216 4032 383393 4060
rect 380216 4020 380222 4032
rect 383381 4029 383393 4032
rect 383427 4029 383439 4063
rect 383381 4023 383439 4029
rect 383657 4063 383715 4069
rect 383657 4029 383669 4063
rect 383703 4060 383715 4063
rect 447410 4060 447416 4072
rect 383703 4032 447416 4060
rect 383703 4029 383715 4032
rect 383657 4023 383715 4029
rect 447410 4020 447416 4032
rect 447468 4020 447474 4072
rect 382829 3995 382887 4001
rect 382829 3992 382841 3995
rect 380084 3964 382841 3992
rect 382829 3961 382841 3964
rect 382875 3961 382887 3995
rect 382829 3955 382887 3961
rect 382918 3952 382924 4004
rect 382976 3992 382982 4004
rect 475746 3992 475752 4004
rect 382976 3964 475752 3992
rect 382976 3952 382982 3964
rect 475746 3952 475752 3964
rect 475804 3952 475810 4004
rect 123478 3924 123484 3936
rect 117976 3896 123484 3924
rect 117869 3887 117927 3893
rect 123478 3884 123484 3896
rect 123536 3884 123542 3936
rect 124122 3884 124128 3936
rect 124180 3924 124186 3936
rect 127434 3924 127440 3936
rect 124180 3896 127440 3924
rect 124180 3884 124186 3896
rect 127434 3884 127440 3896
rect 127492 3884 127498 3936
rect 192018 3924 192024 3936
rect 127636 3896 192024 3924
rect 17034 3816 17040 3868
rect 17092 3856 17098 3868
rect 26421 3859 26479 3865
rect 17092 3828 26234 3856
rect 17092 3816 17098 3828
rect 19426 3748 19432 3800
rect 19484 3788 19490 3800
rect 20530 3788 20536 3800
rect 19484 3760 20536 3788
rect 19484 3748 19490 3760
rect 20530 3748 20536 3760
rect 20588 3748 20594 3800
rect 26206 3788 26234 3828
rect 26421 3825 26433 3859
rect 26467 3856 26479 3859
rect 27798 3856 27804 3868
rect 26467 3828 27804 3856
rect 26467 3825 26479 3828
rect 26421 3819 26479 3825
rect 27798 3816 27804 3828
rect 27856 3816 27862 3868
rect 67542 3816 67548 3868
rect 67600 3856 67606 3868
rect 71685 3859 71743 3865
rect 67600 3828 71636 3856
rect 67600 3816 67606 3828
rect 36078 3788 36084 3800
rect 26206 3760 36084 3788
rect 36078 3748 36084 3760
rect 36136 3748 36142 3800
rect 60458 3748 60464 3800
rect 60516 3788 60522 3800
rect 62117 3791 62175 3797
rect 62117 3788 62129 3791
rect 60516 3760 62129 3788
rect 60516 3748 60522 3760
rect 62117 3757 62129 3760
rect 62163 3757 62175 3791
rect 62117 3751 62175 3757
rect 70210 3748 70216 3800
rect 70268 3788 70274 3800
rect 71608 3788 71636 3828
rect 71685 3825 71697 3859
rect 71731 3856 71743 3859
rect 80882 3856 80888 3868
rect 71731 3828 80888 3856
rect 71731 3825 71743 3828
rect 71685 3819 71743 3825
rect 80882 3816 80888 3828
rect 80940 3816 80946 3868
rect 81342 3816 81348 3868
rect 81400 3856 81406 3868
rect 103885 3859 103943 3865
rect 103885 3856 103897 3859
rect 81400 3828 103897 3856
rect 81400 3816 81406 3828
rect 103885 3825 103897 3828
rect 103931 3825 103943 3859
rect 108301 3859 108359 3865
rect 108301 3856 108313 3859
rect 103885 3819 103943 3825
rect 103992 3828 108313 3856
rect 82078 3788 82084 3800
rect 70268 3760 71544 3788
rect 71608 3760 82084 3788
rect 70268 3748 70274 3760
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 26237 3723 26295 3729
rect 26237 3720 26249 3723
rect 12308 3692 26249 3720
rect 12308 3680 12314 3692
rect 26237 3689 26249 3692
rect 26283 3689 26295 3723
rect 30558 3720 30564 3732
rect 26237 3683 26295 3689
rect 26344 3692 30564 3720
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 26344 3652 26372 3692
rect 30558 3680 30564 3692
rect 30616 3680 30622 3732
rect 61930 3680 61936 3732
rect 61988 3720 61994 3732
rect 70302 3720 70308 3732
rect 61988 3692 70308 3720
rect 61988 3680 61994 3692
rect 70302 3680 70308 3692
rect 70360 3680 70366 3732
rect 71516 3720 71544 3760
rect 82078 3748 82084 3760
rect 82136 3748 82142 3800
rect 82722 3748 82728 3800
rect 82780 3788 82786 3800
rect 103992 3788 104020 3828
rect 108301 3825 108313 3828
rect 108347 3825 108359 3859
rect 108301 3819 108359 3825
rect 108390 3816 108396 3868
rect 108448 3856 108454 3868
rect 111889 3859 111947 3865
rect 111889 3856 111901 3859
rect 108448 3828 111901 3856
rect 108448 3816 108454 3828
rect 111889 3825 111901 3828
rect 111935 3825 111947 3859
rect 111889 3819 111947 3825
rect 111981 3859 112039 3865
rect 111981 3825 111993 3859
rect 112027 3856 112039 3859
rect 118053 3859 118111 3865
rect 118053 3856 118065 3859
rect 112027 3828 118065 3856
rect 112027 3825 112039 3828
rect 111981 3819 112039 3825
rect 118053 3825 118065 3828
rect 118099 3825 118111 3859
rect 118053 3819 118111 3825
rect 118602 3816 118608 3868
rect 118660 3856 118666 3868
rect 127636 3856 127664 3896
rect 192018 3884 192024 3896
rect 192076 3884 192082 3936
rect 194502 3884 194508 3936
rect 194560 3924 194566 3936
rect 204993 3927 205051 3933
rect 204993 3924 205005 3927
rect 194560 3896 205005 3924
rect 194560 3884 194566 3896
rect 204993 3893 205005 3896
rect 205039 3893 205051 3927
rect 204993 3887 205051 3893
rect 211062 3884 211068 3936
rect 211120 3924 211126 3936
rect 387150 3924 387156 3936
rect 211120 3896 387156 3924
rect 211120 3884 211126 3896
rect 387150 3884 387156 3896
rect 387208 3884 387214 3936
rect 199102 3856 199108 3868
rect 118660 3828 127664 3856
rect 127728 3828 199108 3856
rect 118660 3816 118666 3828
rect 82780 3760 104020 3788
rect 104069 3791 104127 3797
rect 82780 3748 82786 3760
rect 104069 3757 104081 3791
rect 104115 3788 104127 3791
rect 105722 3788 105728 3800
rect 104115 3760 105728 3788
rect 104115 3757 104127 3760
rect 104069 3751 104127 3757
rect 105722 3748 105728 3760
rect 105780 3748 105786 3800
rect 105814 3748 105820 3800
rect 105872 3788 105878 3800
rect 108117 3791 108175 3797
rect 108117 3788 108129 3791
rect 105872 3760 108129 3788
rect 105872 3748 105878 3760
rect 108117 3757 108129 3760
rect 108163 3757 108175 3791
rect 108117 3751 108175 3757
rect 108209 3791 108267 3797
rect 108209 3757 108221 3791
rect 108255 3788 108267 3791
rect 111705 3791 111763 3797
rect 111705 3788 111717 3791
rect 108255 3760 111717 3788
rect 108255 3757 108267 3760
rect 108209 3751 108267 3757
rect 111705 3757 111717 3760
rect 111751 3757 111763 3791
rect 111705 3751 111763 3757
rect 117961 3791 118019 3797
rect 117961 3757 117973 3791
rect 118007 3788 118019 3791
rect 124674 3788 124680 3800
rect 118007 3760 124680 3788
rect 118007 3757 118019 3760
rect 117961 3751 118019 3757
rect 124674 3748 124680 3760
rect 124732 3748 124738 3800
rect 125502 3748 125508 3800
rect 125560 3788 125566 3800
rect 127437 3791 127495 3797
rect 127437 3788 127449 3791
rect 125560 3760 127449 3788
rect 125560 3748 125566 3760
rect 127437 3757 127449 3760
rect 127483 3757 127495 3791
rect 127437 3751 127495 3757
rect 127529 3791 127587 3797
rect 127529 3757 127541 3791
rect 127575 3788 127587 3791
rect 127728 3788 127756 3828
rect 199102 3816 199108 3828
rect 199160 3816 199166 3868
rect 202690 3856 202696 3868
rect 200086 3828 202696 3856
rect 127575 3760 127756 3788
rect 127575 3757 127587 3760
rect 127529 3751 127587 3757
rect 127802 3748 127808 3800
rect 127860 3788 127866 3800
rect 200086 3788 200114 3828
rect 202690 3816 202696 3828
rect 202748 3816 202754 3868
rect 213822 3816 213828 3868
rect 213880 3856 213886 3868
rect 394234 3856 394240 3868
rect 213880 3828 394240 3856
rect 213880 3816 213886 3828
rect 394234 3816 394240 3828
rect 394292 3816 394298 3868
rect 401318 3856 401324 3868
rect 398668 3828 401324 3856
rect 209774 3788 209780 3800
rect 127860 3760 200114 3788
rect 200408 3760 209780 3788
rect 127860 3748 127866 3760
rect 89162 3720 89168 3732
rect 71516 3692 89168 3720
rect 89162 3680 89168 3692
rect 89220 3680 89226 3732
rect 89257 3723 89315 3729
rect 89257 3689 89269 3723
rect 89303 3720 89315 3723
rect 89303 3692 92980 3720
rect 89303 3689 89315 3692
rect 89257 3683 89315 3689
rect 29086 3652 29092 3664
rect 7708 3624 26372 3652
rect 26436 3624 29092 3652
rect 7708 3612 7714 3624
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 26436 3584 26464 3624
rect 29086 3612 29092 3624
rect 29144 3612 29150 3664
rect 57698 3612 57704 3664
rect 57756 3652 57762 3664
rect 63218 3652 63224 3664
rect 57756 3624 63224 3652
rect 57756 3612 57762 3624
rect 63218 3612 63224 3624
rect 63276 3612 63282 3664
rect 68922 3612 68928 3664
rect 68980 3652 68986 3664
rect 84470 3652 84476 3664
rect 68980 3624 84476 3652
rect 68980 3612 68986 3624
rect 84470 3612 84476 3624
rect 84528 3612 84534 3664
rect 86862 3612 86868 3664
rect 86920 3652 86926 3664
rect 87509 3655 87567 3661
rect 87509 3652 87521 3655
rect 86920 3624 87521 3652
rect 86920 3612 86926 3624
rect 87509 3621 87521 3624
rect 87555 3621 87567 3655
rect 87509 3615 87567 3621
rect 87598 3612 87604 3664
rect 87656 3652 87662 3664
rect 92952 3652 92980 3692
rect 93118 3680 93124 3732
rect 93176 3720 93182 3732
rect 128170 3720 128176 3732
rect 93176 3692 128176 3720
rect 93176 3680 93182 3692
rect 128170 3680 128176 3692
rect 128228 3680 128234 3732
rect 132037 3723 132095 3729
rect 128280 3692 131988 3720
rect 122282 3652 122288 3664
rect 87656 3624 92888 3652
rect 92952 3624 122288 3652
rect 87656 3612 87662 3624
rect 2924 3556 26464 3584
rect 2924 3544 2930 3556
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 37090 3584 37096 3596
rect 36044 3556 37096 3584
rect 36044 3544 36050 3556
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45370 3584 45376 3596
rect 44324 3556 45376 3584
rect 44324 3544 44330 3556
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 60550 3544 60556 3596
rect 60608 3584 60614 3596
rect 60608 3556 60964 3584
rect 60608 3544 60614 3556
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 26421 3519 26479 3525
rect 26421 3516 26433 3519
rect 1728 3488 26433 3516
rect 1728 3476 1734 3488
rect 26421 3485 26433 3488
rect 26467 3485 26479 3519
rect 26421 3479 26479 3485
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 28810 3516 28816 3528
rect 27764 3488 28816 3516
rect 27764 3476 27770 3488
rect 28810 3476 28816 3488
rect 28868 3476 28874 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53742 3516 53748 3528
rect 52512 3488 53748 3516
rect 52512 3476 52518 3488
rect 53742 3476 53748 3488
rect 53800 3476 53806 3528
rect 54018 3476 54024 3528
rect 54076 3516 54082 3528
rect 54938 3516 54944 3528
rect 54076 3488 54944 3516
rect 54076 3476 54082 3488
rect 54938 3476 54944 3488
rect 54996 3476 55002 3528
rect 57882 3476 57888 3528
rect 57940 3516 57946 3528
rect 60826 3516 60832 3528
rect 57940 3488 60832 3516
rect 57940 3476 57946 3488
rect 60826 3476 60832 3488
rect 60884 3476 60890 3528
rect 60936 3516 60964 3556
rect 62022 3544 62028 3596
rect 62080 3584 62086 3596
rect 71498 3584 71504 3596
rect 62080 3556 71504 3584
rect 62080 3544 62086 3556
rect 71498 3544 71504 3556
rect 71556 3544 71562 3596
rect 71682 3544 71688 3596
rect 71740 3584 71746 3596
rect 92750 3584 92756 3596
rect 71740 3556 92756 3584
rect 71740 3544 71746 3556
rect 92750 3544 92756 3556
rect 92808 3544 92814 3596
rect 92860 3584 92888 3624
rect 122282 3612 122288 3624
rect 122340 3612 122346 3664
rect 126882 3612 126888 3664
rect 126940 3652 126946 3664
rect 128280 3652 128308 3692
rect 126940 3624 128308 3652
rect 126940 3612 126946 3624
rect 129642 3612 129648 3664
rect 129700 3652 129706 3664
rect 131960 3652 131988 3692
rect 132037 3689 132049 3723
rect 132083 3720 132095 3723
rect 200117 3723 200175 3729
rect 200117 3720 200129 3723
rect 132083 3692 200129 3720
rect 132083 3689 132095 3692
rect 132037 3683 132095 3689
rect 200117 3689 200129 3692
rect 200163 3689 200175 3723
rect 200117 3683 200175 3689
rect 200408 3652 200436 3760
rect 209774 3748 209780 3760
rect 209832 3748 209838 3800
rect 217962 3748 217968 3800
rect 218020 3788 218026 3800
rect 398668 3788 398696 3828
rect 401318 3816 401324 3828
rect 401376 3816 401382 3868
rect 218020 3760 398696 3788
rect 218020 3748 218026 3760
rect 398834 3748 398840 3800
rect 398892 3788 398898 3800
rect 400122 3788 400128 3800
rect 398892 3760 400128 3788
rect 398892 3748 398898 3760
rect 400122 3748 400128 3760
rect 400180 3748 400186 3800
rect 220722 3680 220728 3732
rect 220780 3720 220786 3732
rect 408402 3720 408408 3732
rect 220780 3692 408408 3720
rect 220780 3680 220786 3692
rect 408402 3680 408408 3692
rect 408460 3680 408466 3732
rect 129700 3624 131896 3652
rect 131960 3624 200436 3652
rect 200577 3655 200635 3661
rect 129700 3612 129706 3624
rect 93946 3584 93952 3596
rect 92860 3556 93952 3584
rect 93946 3544 93952 3556
rect 94004 3544 94010 3596
rect 94498 3544 94504 3596
rect 94556 3584 94562 3596
rect 131758 3584 131764 3596
rect 94556 3556 131764 3584
rect 94556 3544 94562 3556
rect 131758 3544 131764 3556
rect 131816 3544 131822 3596
rect 131868 3584 131896 3624
rect 200577 3621 200589 3655
rect 200623 3652 200635 3655
rect 212166 3652 212172 3664
rect 200623 3624 212172 3652
rect 200623 3621 200635 3624
rect 200577 3615 200635 3621
rect 212166 3612 212172 3624
rect 212224 3612 212230 3664
rect 224862 3612 224868 3664
rect 224920 3652 224926 3664
rect 415486 3652 415492 3664
rect 224920 3624 415492 3652
rect 224920 3612 224926 3624
rect 415486 3612 415492 3624
rect 415544 3612 415550 3664
rect 418798 3612 418804 3664
rect 418856 3652 418862 3664
rect 568022 3652 568028 3664
rect 418856 3624 568028 3652
rect 418856 3612 418862 3624
rect 568022 3612 568028 3624
rect 568080 3612 568086 3664
rect 213362 3584 213368 3596
rect 131868 3556 213368 3584
rect 213362 3544 213368 3556
rect 213420 3544 213426 3596
rect 227622 3544 227628 3596
rect 227680 3584 227686 3596
rect 422570 3584 422576 3596
rect 227680 3556 422576 3584
rect 227680 3544 227686 3556
rect 422570 3544 422576 3556
rect 422628 3544 422634 3596
rect 429654 3584 429660 3596
rect 423600 3556 429660 3584
rect 67910 3516 67916 3528
rect 60936 3488 67916 3516
rect 67910 3476 67916 3488
rect 67968 3476 67974 3528
rect 68830 3476 68836 3528
rect 68888 3516 68894 3528
rect 85666 3516 85672 3528
rect 68888 3488 85672 3516
rect 68888 3476 68894 3488
rect 85666 3476 85672 3488
rect 85724 3476 85730 3528
rect 86770 3476 86776 3528
rect 86828 3516 86834 3528
rect 88889 3519 88947 3525
rect 88889 3516 88901 3519
rect 86828 3488 88901 3516
rect 86828 3476 86834 3488
rect 88889 3485 88901 3488
rect 88935 3485 88947 3519
rect 88889 3479 88947 3485
rect 88978 3476 88984 3528
rect 89036 3516 89042 3528
rect 90358 3516 90364 3528
rect 89036 3488 90364 3516
rect 89036 3476 89042 3488
rect 90358 3476 90364 3488
rect 90416 3476 90422 3528
rect 90453 3519 90511 3525
rect 90453 3485 90465 3519
rect 90499 3516 90511 3519
rect 117961 3519 118019 3525
rect 117961 3516 117973 3519
rect 90499 3488 117973 3516
rect 90499 3485 90511 3488
rect 90453 3479 90511 3485
rect 117961 3485 117973 3488
rect 118007 3485 118019 3519
rect 117961 3479 118019 3485
rect 119338 3476 119344 3528
rect 119396 3516 119402 3528
rect 121086 3516 121092 3528
rect 119396 3488 121092 3516
rect 119396 3476 119402 3488
rect 121086 3476 121092 3488
rect 121144 3476 121150 3528
rect 121181 3519 121239 3525
rect 121181 3485 121193 3519
rect 121227 3516 121239 3519
rect 127713 3519 127771 3525
rect 127713 3516 127725 3519
rect 121227 3488 127725 3516
rect 121227 3485 121239 3488
rect 121181 3479 121239 3485
rect 127713 3485 127725 3488
rect 127759 3485 127771 3519
rect 127713 3479 127771 3485
rect 127805 3519 127863 3525
rect 127805 3485 127817 3519
rect 127851 3516 127863 3519
rect 132037 3519 132095 3525
rect 132037 3516 132049 3519
rect 127851 3488 132049 3516
rect 127851 3485 127863 3488
rect 127805 3479 127863 3485
rect 132037 3485 132049 3488
rect 132083 3485 132095 3519
rect 132037 3479 132095 3485
rect 132402 3476 132408 3528
rect 132460 3516 132466 3528
rect 220446 3516 220452 3528
rect 132460 3488 220452 3516
rect 132460 3476 132466 3488
rect 220446 3476 220452 3488
rect 220504 3476 220510 3528
rect 230382 3476 230388 3528
rect 230440 3516 230446 3528
rect 423600 3516 423628 3556
rect 429654 3544 429660 3556
rect 429712 3544 429718 3596
rect 489914 3544 489920 3596
rect 489972 3584 489978 3596
rect 491110 3584 491116 3596
rect 489972 3556 491116 3584
rect 489972 3544 489978 3556
rect 491110 3544 491116 3556
rect 491168 3544 491174 3596
rect 230440 3488 423628 3516
rect 230440 3476 230446 3488
rect 423674 3476 423680 3528
rect 423732 3516 423738 3528
rect 424962 3516 424968 3528
rect 423732 3488 424968 3516
rect 423732 3476 423738 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 448514 3476 448520 3528
rect 448572 3516 448578 3528
rect 449802 3516 449808 3528
rect 448572 3488 449808 3516
rect 448572 3476 448578 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 456794 3476 456800 3528
rect 456852 3516 456858 3528
rect 458082 3516 458088 3528
rect 456852 3488 458088 3516
rect 456852 3476 456858 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 27614 3448 27620 3460
rect 624 3420 27620 3448
rect 624 3408 630 3420
rect 27614 3408 27620 3420
rect 27672 3408 27678 3460
rect 57790 3408 57796 3460
rect 57848 3448 57854 3460
rect 62022 3448 62028 3460
rect 57848 3420 62028 3448
rect 57848 3408 57854 3420
rect 62022 3408 62028 3420
rect 62080 3408 62086 3460
rect 62117 3451 62175 3457
rect 62117 3417 62129 3451
rect 62163 3448 62175 3451
rect 69106 3448 69112 3460
rect 62163 3420 69112 3448
rect 62163 3417 62175 3420
rect 62117 3411 62175 3417
rect 69106 3408 69112 3420
rect 69164 3408 69170 3460
rect 71590 3408 71596 3460
rect 71648 3448 71654 3460
rect 91554 3448 91560 3460
rect 71648 3420 91560 3448
rect 71648 3408 71654 3420
rect 91554 3408 91560 3420
rect 91612 3408 91618 3460
rect 92382 3408 92388 3460
rect 92440 3448 92446 3460
rect 135254 3448 135260 3460
rect 92440 3420 135260 3448
rect 92440 3408 92446 3420
rect 135254 3408 135260 3420
rect 135312 3408 135318 3460
rect 137922 3408 137928 3460
rect 137980 3448 137986 3460
rect 231026 3448 231032 3460
rect 137980 3420 231032 3448
rect 137980 3408 137986 3420
rect 231026 3408 231032 3420
rect 231084 3408 231090 3460
rect 237282 3408 237288 3460
rect 237340 3448 237346 3460
rect 443822 3448 443828 3460
rect 237340 3420 443828 3448
rect 237340 3408 237346 3420
rect 443822 3408 443828 3420
rect 443880 3408 443886 3460
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 9582 3380 9588 3392
rect 8812 3352 9588 3380
rect 8812 3340 8818 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 10962 3380 10968 3392
rect 10008 3352 10968 3380
rect 10008 3340 10014 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 12342 3380 12348 3392
rect 11204 3352 12348 3380
rect 11204 3340 11210 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 16482 3380 16488 3392
rect 15988 3352 16488 3380
rect 15988 3340 15994 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 19242 3380 19248 3392
rect 18288 3352 19248 3380
rect 18288 3340 18294 3352
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 24762 3380 24768 3392
rect 24268 3352 24768 3380
rect 24268 3340 24274 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25314 3340 25320 3392
rect 25372 3380 25378 3392
rect 26142 3380 26148 3392
rect 25372 3352 26148 3380
rect 25372 3340 25378 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 59262 3340 59268 3392
rect 59320 3380 59326 3392
rect 64322 3380 64328 3392
rect 59320 3352 64328 3380
rect 59320 3340 59326 3352
rect 64322 3340 64328 3352
rect 64380 3340 64386 3392
rect 66162 3340 66168 3392
rect 66220 3380 66226 3392
rect 71685 3383 71743 3389
rect 71685 3380 71697 3383
rect 66220 3352 71697 3380
rect 66220 3340 66226 3352
rect 71685 3349 71697 3352
rect 71731 3349 71743 3383
rect 78582 3380 78588 3392
rect 71685 3343 71743 3349
rect 73908 3352 78588 3380
rect 63126 3272 63132 3324
rect 63184 3312 63190 3324
rect 73798 3312 73804 3324
rect 63184 3284 73804 3312
rect 63184 3272 63190 3284
rect 73798 3272 73804 3284
rect 73856 3272 73862 3324
rect 63402 3204 63408 3256
rect 63460 3244 63466 3256
rect 72602 3244 72608 3256
rect 63460 3216 72608 3244
rect 63460 3204 63466 3216
rect 72602 3204 72608 3216
rect 72660 3204 72666 3256
rect 56410 3136 56416 3188
rect 56468 3176 56474 3188
rect 59630 3176 59636 3188
rect 56468 3148 59636 3176
rect 56468 3136 56474 3148
rect 59630 3136 59636 3148
rect 59688 3136 59694 3188
rect 60642 3136 60648 3188
rect 60700 3176 60706 3188
rect 66714 3176 66720 3188
rect 60700 3148 66720 3176
rect 60700 3136 60706 3148
rect 66714 3136 66720 3148
rect 66772 3136 66778 3188
rect 65978 3068 65984 3120
rect 66036 3108 66042 3120
rect 73908 3108 73936 3352
rect 78582 3340 78588 3352
rect 78640 3340 78646 3392
rect 78674 3340 78680 3392
rect 78732 3380 78738 3392
rect 104069 3383 104127 3389
rect 104069 3380 104081 3383
rect 78732 3352 104081 3380
rect 78732 3340 78738 3352
rect 104069 3349 104081 3352
rect 104115 3349 104127 3383
rect 104069 3343 104127 3349
rect 104158 3340 104164 3392
rect 104216 3380 104222 3392
rect 106918 3380 106924 3392
rect 104216 3352 106924 3380
rect 104216 3340 104222 3352
rect 106918 3340 106924 3352
rect 106976 3340 106982 3392
rect 107562 3340 107568 3392
rect 107620 3380 107626 3392
rect 108206 3380 108212 3392
rect 107620 3352 108212 3380
rect 107620 3340 107626 3352
rect 108206 3340 108212 3352
rect 108264 3340 108270 3392
rect 108301 3383 108359 3389
rect 108301 3349 108313 3383
rect 108347 3380 108359 3383
rect 115198 3380 115204 3392
rect 108347 3352 115204 3380
rect 108347 3349 108359 3352
rect 108301 3343 108359 3349
rect 115198 3340 115204 3352
rect 115256 3340 115262 3392
rect 177850 3380 177856 3392
rect 117792 3352 177856 3380
rect 87966 3312 87972 3324
rect 66036 3080 73936 3108
rect 74000 3284 87972 3312
rect 66036 3068 66042 3080
rect 70394 3000 70400 3052
rect 70452 3040 70458 3052
rect 74000 3040 74028 3284
rect 87966 3272 87972 3284
rect 88024 3272 88030 3324
rect 88061 3315 88119 3321
rect 88061 3281 88073 3315
rect 88107 3312 88119 3315
rect 90361 3315 90419 3321
rect 90361 3312 90373 3315
rect 88107 3284 90373 3312
rect 88107 3281 88119 3284
rect 88061 3275 88119 3281
rect 90361 3281 90373 3284
rect 90407 3281 90419 3315
rect 90361 3275 90419 3281
rect 90450 3272 90456 3324
rect 90508 3312 90514 3324
rect 116394 3312 116400 3324
rect 90508 3284 116400 3312
rect 90508 3272 90514 3284
rect 116394 3272 116400 3284
rect 116452 3272 116458 3324
rect 75730 3204 75736 3256
rect 75788 3244 75794 3256
rect 101030 3244 101036 3256
rect 75788 3216 101036 3244
rect 75788 3204 75794 3216
rect 101030 3204 101036 3216
rect 101088 3204 101094 3256
rect 101398 3204 101404 3256
rect 101456 3244 101462 3256
rect 104529 3247 104587 3253
rect 104529 3244 104541 3247
rect 101456 3216 104541 3244
rect 101456 3204 101462 3216
rect 104529 3213 104541 3216
rect 104575 3213 104587 3247
rect 108301 3247 108359 3253
rect 108301 3244 108313 3247
rect 104529 3207 104587 3213
rect 104636 3216 108313 3244
rect 77202 3136 77208 3188
rect 77260 3176 77266 3188
rect 102226 3176 102232 3188
rect 77260 3148 102232 3176
rect 77260 3136 77266 3148
rect 102226 3136 102232 3148
rect 102284 3136 102290 3188
rect 104636 3176 104664 3216
rect 108301 3213 108313 3216
rect 108347 3213 108359 3247
rect 108301 3207 108359 3213
rect 108390 3204 108396 3256
rect 108448 3244 108454 3256
rect 111981 3247 112039 3253
rect 111981 3244 111993 3247
rect 108448 3216 111993 3244
rect 108448 3204 108454 3216
rect 111981 3213 111993 3216
rect 112027 3213 112039 3247
rect 111981 3207 112039 3213
rect 112070 3204 112076 3256
rect 112128 3244 112134 3256
rect 117792 3244 117820 3352
rect 177850 3340 177856 3352
rect 177908 3340 177914 3392
rect 185673 3383 185731 3389
rect 177960 3352 185624 3380
rect 117869 3315 117927 3321
rect 117869 3281 117881 3315
rect 117915 3312 117927 3315
rect 174262 3312 174268 3324
rect 117915 3284 174268 3312
rect 117915 3281 117927 3284
rect 117869 3275 117927 3281
rect 174262 3272 174268 3284
rect 174320 3272 174326 3324
rect 175918 3272 175924 3324
rect 175976 3312 175982 3324
rect 177960 3312 177988 3352
rect 185489 3315 185547 3321
rect 185489 3312 185501 3315
rect 175976 3284 177988 3312
rect 178052 3284 185501 3312
rect 175976 3272 175982 3284
rect 112128 3216 117820 3244
rect 118053 3247 118111 3253
rect 112128 3204 112134 3216
rect 118053 3213 118065 3247
rect 118099 3244 118111 3247
rect 167178 3244 167184 3256
rect 118099 3216 167184 3244
rect 118099 3213 118111 3216
rect 118053 3207 118111 3213
rect 167178 3204 167184 3216
rect 167236 3204 167242 3256
rect 177298 3204 177304 3256
rect 177356 3244 177362 3256
rect 178052 3244 178080 3284
rect 185489 3281 185501 3284
rect 185535 3281 185547 3315
rect 185596 3312 185624 3352
rect 185673 3349 185685 3383
rect 185719 3380 185731 3383
rect 200577 3383 200635 3389
rect 200577 3380 200589 3383
rect 185719 3352 200589 3380
rect 185719 3349 185731 3352
rect 185673 3343 185731 3349
rect 200577 3349 200589 3352
rect 200623 3349 200635 3383
rect 355873 3383 355931 3389
rect 355873 3380 355885 3383
rect 200577 3343 200635 3349
rect 204916 3352 355885 3380
rect 194229 3315 194287 3321
rect 185596 3284 194180 3312
rect 185489 3275 185547 3281
rect 177356 3216 178080 3244
rect 178129 3247 178187 3253
rect 177356 3204 177362 3216
rect 178129 3213 178141 3247
rect 178175 3244 178187 3247
rect 193214 3244 193220 3256
rect 178175 3216 193220 3244
rect 178175 3213 178187 3216
rect 178129 3207 178187 3213
rect 193214 3204 193220 3216
rect 193272 3204 193278 3256
rect 194152 3244 194180 3284
rect 194229 3281 194241 3315
rect 194275 3312 194287 3315
rect 194275 3284 195376 3312
rect 194275 3281 194287 3284
rect 194229 3275 194287 3281
rect 195149 3247 195207 3253
rect 195149 3244 195161 3247
rect 194152 3216 195161 3244
rect 195149 3213 195161 3216
rect 195195 3213 195207 3247
rect 195149 3207 195207 3213
rect 160094 3176 160100 3188
rect 102336 3148 104664 3176
rect 104728 3148 160100 3176
rect 74350 3068 74356 3120
rect 74408 3108 74414 3120
rect 98638 3108 98644 3120
rect 74408 3080 98644 3108
rect 74408 3068 74414 3080
rect 98638 3068 98644 3080
rect 98696 3068 98702 3120
rect 102336 3108 102364 3148
rect 99944 3080 102364 3108
rect 70452 3012 74028 3040
rect 70452 3000 70458 3012
rect 75822 3000 75828 3052
rect 75880 3040 75886 3052
rect 99834 3040 99840 3052
rect 75880 3012 99840 3040
rect 75880 3000 75886 3012
rect 99834 3000 99840 3012
rect 99892 3000 99898 3052
rect 56502 2932 56508 2984
rect 56560 2972 56566 2984
rect 58434 2972 58440 2984
rect 56560 2944 58440 2972
rect 56560 2932 56566 2944
rect 58434 2932 58440 2944
rect 58492 2932 58498 2984
rect 74258 2932 74264 2984
rect 74316 2972 74322 2984
rect 97442 2972 97448 2984
rect 74316 2944 97448 2972
rect 74316 2932 74322 2944
rect 97442 2932 97448 2944
rect 97500 2932 97506 2984
rect 97902 2932 97908 2984
rect 97960 2972 97966 2984
rect 99944 2972 99972 3080
rect 103422 3068 103428 3120
rect 103480 3108 103486 3120
rect 104728 3108 104756 3148
rect 160094 3136 160100 3148
rect 160152 3136 160158 3188
rect 160738 3136 160744 3188
rect 160796 3176 160802 3188
rect 160796 3148 161474 3176
rect 160796 3136 160802 3148
rect 153010 3108 153016 3120
rect 103480 3080 104756 3108
rect 104820 3080 153016 3108
rect 103480 3068 103486 3080
rect 100662 3000 100668 3052
rect 100720 3040 100726 3052
rect 104820 3040 104848 3080
rect 153010 3068 153016 3080
rect 153068 3068 153074 3120
rect 155218 3068 155224 3120
rect 155276 3108 155282 3120
rect 161290 3108 161296 3120
rect 155276 3080 161296 3108
rect 155276 3068 155282 3080
rect 161290 3068 161296 3080
rect 161348 3068 161354 3120
rect 161446 3108 161474 3148
rect 170398 3136 170404 3188
rect 170456 3176 170462 3188
rect 189718 3176 189724 3188
rect 170456 3148 189724 3176
rect 170456 3136 170462 3148
rect 189718 3136 189724 3148
rect 189776 3136 189782 3188
rect 190362 3136 190368 3188
rect 190420 3176 190426 3188
rect 195241 3179 195299 3185
rect 195241 3176 195253 3179
rect 190420 3148 195253 3176
rect 190420 3136 190426 3148
rect 195241 3145 195253 3148
rect 195287 3145 195299 3179
rect 195348 3176 195376 3284
rect 197262 3272 197268 3324
rect 197320 3312 197326 3324
rect 204916 3312 204944 3352
rect 355873 3349 355885 3352
rect 355919 3349 355931 3383
rect 355873 3343 355931 3349
rect 355962 3340 355968 3392
rect 356020 3380 356026 3392
rect 356020 3352 356192 3380
rect 356020 3340 356026 3352
rect 197320 3284 204944 3312
rect 204993 3315 205051 3321
rect 197320 3272 197326 3284
rect 204993 3281 205005 3315
rect 205039 3312 205051 3315
rect 349065 3315 349123 3321
rect 349065 3312 349077 3315
rect 205039 3284 349077 3312
rect 205039 3281 205051 3284
rect 204993 3275 205051 3281
rect 349065 3281 349077 3284
rect 349111 3281 349123 3315
rect 349065 3275 349123 3281
rect 349154 3272 349160 3324
rect 349212 3312 349218 3324
rect 350442 3312 350448 3324
rect 349212 3284 350448 3312
rect 349212 3272 349218 3284
rect 350442 3272 350448 3284
rect 350500 3272 350506 3324
rect 351178 3272 351184 3324
rect 351236 3312 351242 3324
rect 351236 3284 351776 3312
rect 351236 3272 351242 3284
rect 195425 3247 195483 3253
rect 195425 3213 195437 3247
rect 195471 3244 195483 3247
rect 344554 3244 344560 3256
rect 195471 3216 344560 3244
rect 195471 3213 195483 3216
rect 195425 3207 195483 3213
rect 344554 3204 344560 3216
rect 344612 3204 344618 3256
rect 344649 3247 344707 3253
rect 344649 3213 344661 3247
rect 344695 3244 344707 3247
rect 349801 3247 349859 3253
rect 349801 3244 349813 3247
rect 344695 3216 349813 3244
rect 344695 3213 344707 3216
rect 344649 3207 344707 3213
rect 349801 3213 349813 3216
rect 349847 3213 349859 3247
rect 349801 3207 349859 3213
rect 349893 3247 349951 3253
rect 349893 3213 349905 3247
rect 349939 3244 349951 3247
rect 351638 3244 351644 3256
rect 349939 3216 351644 3244
rect 349939 3213 349951 3216
rect 349893 3207 349951 3213
rect 351638 3204 351644 3216
rect 351696 3204 351702 3256
rect 351748 3244 351776 3284
rect 351822 3272 351828 3324
rect 351880 3312 351886 3324
rect 356164 3312 356192 3352
rect 358078 3340 358084 3392
rect 358136 3380 358142 3392
rect 369213 3383 369271 3389
rect 369213 3380 369225 3383
rect 358136 3352 369225 3380
rect 358136 3340 358142 3352
rect 369213 3349 369225 3352
rect 369259 3349 369271 3383
rect 369213 3343 369271 3349
rect 369486 3340 369492 3392
rect 369544 3380 369550 3392
rect 373077 3383 373135 3389
rect 373077 3380 373089 3383
rect 369544 3352 373089 3380
rect 369544 3340 369550 3352
rect 373077 3349 373089 3352
rect 373123 3349 373135 3383
rect 373077 3343 373135 3349
rect 373258 3340 373264 3392
rect 373316 3380 373322 3392
rect 426158 3380 426164 3392
rect 373316 3352 426164 3380
rect 373316 3340 373322 3352
rect 426158 3340 426164 3352
rect 426216 3340 426222 3392
rect 383470 3312 383476 3324
rect 351880 3284 356100 3312
rect 356164 3284 383476 3312
rect 351880 3272 351886 3284
rect 355870 3244 355876 3256
rect 351748 3216 355876 3244
rect 355870 3204 355876 3216
rect 355928 3204 355934 3256
rect 356072 3244 356100 3284
rect 383470 3272 383476 3284
rect 383528 3272 383534 3324
rect 383562 3272 383568 3324
rect 383620 3312 383626 3324
rect 418982 3312 418988 3324
rect 383620 3284 418988 3312
rect 383620 3272 383626 3284
rect 418982 3272 418988 3284
rect 419040 3272 419046 3324
rect 368937 3247 368995 3253
rect 368937 3244 368949 3247
rect 356072 3216 368949 3244
rect 368937 3213 368949 3216
rect 368983 3213 368995 3247
rect 369394 3244 369400 3256
rect 368937 3207 368995 3213
rect 369044 3216 369400 3244
rect 337470 3176 337476 3188
rect 195348 3148 337476 3176
rect 195241 3139 195299 3145
rect 337470 3136 337476 3148
rect 337528 3136 337534 3188
rect 337562 3136 337568 3188
rect 337620 3176 337626 3188
rect 344189 3179 344247 3185
rect 344189 3176 344201 3179
rect 337620 3148 344201 3176
rect 337620 3136 337626 3148
rect 344189 3145 344201 3148
rect 344235 3145 344247 3179
rect 344189 3139 344247 3145
rect 344278 3136 344284 3188
rect 344336 3176 344342 3188
rect 369044 3176 369072 3216
rect 369394 3204 369400 3216
rect 369452 3204 369458 3256
rect 369489 3247 369547 3253
rect 369489 3213 369501 3247
rect 369535 3244 369547 3247
rect 411898 3244 411904 3256
rect 369535 3216 411904 3244
rect 369535 3213 369547 3216
rect 369489 3207 369547 3213
rect 411898 3204 411904 3216
rect 411956 3204 411962 3256
rect 344336 3148 369072 3176
rect 369121 3179 369179 3185
rect 344336 3136 344342 3148
rect 369121 3145 369133 3179
rect 369167 3176 369179 3179
rect 404814 3176 404820 3188
rect 369167 3148 404820 3176
rect 369167 3145 369179 3148
rect 369121 3139 369179 3145
rect 404814 3136 404820 3148
rect 404872 3136 404878 3188
rect 175458 3108 175464 3120
rect 161446 3080 175464 3108
rect 175458 3068 175464 3080
rect 175516 3068 175522 3120
rect 177390 3068 177396 3120
rect 177448 3108 177454 3120
rect 178221 3111 178279 3117
rect 178221 3108 178233 3111
rect 177448 3080 178233 3108
rect 177448 3068 177454 3080
rect 178221 3077 178233 3080
rect 178267 3077 178279 3111
rect 178221 3071 178279 3077
rect 181530 3068 181536 3120
rect 181588 3108 181594 3120
rect 237006 3108 237012 3120
rect 181588 3080 237012 3108
rect 181588 3068 181594 3080
rect 237006 3068 237012 3080
rect 237064 3068 237070 3120
rect 307754 3068 307760 3120
rect 307812 3108 307818 3120
rect 309042 3108 309048 3120
rect 307812 3080 309048 3108
rect 307812 3068 307818 3080
rect 309042 3068 309048 3080
rect 309100 3068 309106 3120
rect 309778 3068 309784 3120
rect 309836 3108 309842 3120
rect 320637 3111 320695 3117
rect 320637 3108 320649 3111
rect 309836 3080 320649 3108
rect 309836 3068 309842 3080
rect 320637 3077 320649 3080
rect 320683 3077 320695 3111
rect 320637 3071 320695 3077
rect 320729 3111 320787 3117
rect 320729 3077 320741 3111
rect 320775 3108 320787 3111
rect 461578 3108 461584 3120
rect 320775 3080 461584 3108
rect 320775 3077 320787 3080
rect 320729 3071 320787 3077
rect 461578 3068 461584 3080
rect 461636 3068 461642 3120
rect 583386 3108 583392 3120
rect 583347 3080 583392 3108
rect 583386 3068 583392 3080
rect 583444 3068 583450 3120
rect 149514 3040 149520 3052
rect 100720 3012 104848 3040
rect 104912 3012 149520 3040
rect 100720 3000 100726 3012
rect 104912 2972 104940 3012
rect 149514 3000 149520 3012
rect 149572 3000 149578 3052
rect 156598 3000 156604 3052
rect 156656 3040 156662 3052
rect 164878 3040 164884 3052
rect 156656 3012 164884 3040
rect 156656 3000 156662 3012
rect 164878 3000 164884 3012
rect 164936 3000 164942 3052
rect 167638 3000 167644 3052
rect 167696 3040 167702 3052
rect 182542 3040 182548 3052
rect 167696 3012 182548 3040
rect 167696 3000 167702 3012
rect 182542 3000 182548 3012
rect 182600 3000 182606 3052
rect 184842 3000 184848 3052
rect 184900 3040 184906 3052
rect 184900 3012 186360 3040
rect 184900 3000 184906 3012
rect 97960 2944 99972 2972
rect 100128 2944 104940 2972
rect 104989 2975 105047 2981
rect 97960 2932 97966 2944
rect 73062 2864 73068 2916
rect 73120 2904 73126 2916
rect 95142 2904 95148 2916
rect 73120 2876 95148 2904
rect 73120 2864 73126 2876
rect 95142 2864 95148 2876
rect 95200 2864 95206 2916
rect 95878 2864 95884 2916
rect 95936 2904 95942 2916
rect 96338 2904 96344 2916
rect 95936 2876 96344 2904
rect 95936 2864 95942 2876
rect 96338 2864 96344 2876
rect 96396 2864 96402 2916
rect 96448 2876 99236 2904
rect 74442 2796 74448 2848
rect 74500 2836 74506 2848
rect 96246 2836 96252 2848
rect 74500 2808 96252 2836
rect 74500 2796 74506 2808
rect 96246 2796 96252 2808
rect 96304 2796 96310 2848
rect 95234 2728 95240 2780
rect 95292 2768 95298 2780
rect 96448 2768 96476 2876
rect 96522 2796 96528 2848
rect 96580 2836 96586 2848
rect 96580 2808 99144 2836
rect 96580 2796 96586 2808
rect 95292 2740 96476 2768
rect 95292 2728 95298 2740
rect 99116 2700 99144 2808
rect 99208 2768 99236 2876
rect 99282 2864 99288 2916
rect 99340 2904 99346 2916
rect 100128 2904 100156 2944
rect 104989 2941 105001 2975
rect 105035 2972 105047 2975
rect 108209 2975 108267 2981
rect 108209 2972 108221 2975
rect 105035 2944 108221 2972
rect 105035 2941 105047 2944
rect 104989 2935 105047 2941
rect 108209 2941 108221 2944
rect 108255 2941 108267 2975
rect 108209 2935 108267 2941
rect 108301 2975 108359 2981
rect 108301 2941 108313 2975
rect 108347 2972 108359 2975
rect 145926 2972 145932 2984
rect 108347 2944 145932 2972
rect 108347 2941 108359 2944
rect 108301 2935 108359 2941
rect 145926 2932 145932 2944
rect 145984 2932 145990 2984
rect 166258 2932 166264 2984
rect 166316 2972 166322 2984
rect 179046 2972 179052 2984
rect 166316 2944 179052 2972
rect 166316 2932 166322 2944
rect 179046 2932 179052 2944
rect 179104 2932 179110 2984
rect 180058 2932 180064 2984
rect 180116 2972 180122 2984
rect 186225 2975 186283 2981
rect 186225 2972 186237 2975
rect 180116 2944 186237 2972
rect 180116 2932 180122 2944
rect 186225 2941 186237 2944
rect 186271 2941 186283 2975
rect 186225 2935 186283 2941
rect 142430 2904 142436 2916
rect 99340 2876 100156 2904
rect 100220 2876 142436 2904
rect 99340 2864 99346 2876
rect 100220 2768 100248 2876
rect 142430 2864 142436 2876
rect 142488 2864 142494 2916
rect 142798 2864 142804 2916
rect 142856 2904 142862 2916
rect 156598 2904 156604 2916
rect 142856 2876 156604 2904
rect 142856 2864 142862 2876
rect 156598 2864 156604 2876
rect 156656 2864 156662 2916
rect 157978 2864 157984 2916
rect 158036 2904 158042 2916
rect 168374 2904 168380 2916
rect 158036 2876 168380 2904
rect 158036 2864 158042 2876
rect 168374 2864 168380 2876
rect 168432 2864 168438 2916
rect 169018 2864 169024 2916
rect 169076 2904 169082 2916
rect 186130 2904 186136 2916
rect 169076 2876 186136 2904
rect 169076 2864 169082 2876
rect 186130 2864 186136 2876
rect 186188 2864 186194 2916
rect 186332 2904 186360 3012
rect 187602 3000 187608 3052
rect 187660 3040 187666 3052
rect 194229 3043 194287 3049
rect 194229 3040 194241 3043
rect 187660 3012 194241 3040
rect 187660 3000 187666 3012
rect 194229 3009 194241 3012
rect 194275 3009 194287 3043
rect 194229 3003 194287 3009
rect 194321 3043 194379 3049
rect 194321 3009 194333 3043
rect 194367 3040 194379 3043
rect 330386 3040 330392 3052
rect 194367 3012 330392 3040
rect 194367 3009 194379 3012
rect 194321 3003 194379 3009
rect 330386 3000 330392 3012
rect 330444 3000 330450 3052
rect 330478 3000 330484 3052
rect 330536 3040 330542 3052
rect 333149 3043 333207 3049
rect 333149 3040 333161 3043
rect 330536 3012 333161 3040
rect 330536 3000 330542 3012
rect 333149 3009 333161 3012
rect 333195 3009 333207 3043
rect 333149 3003 333207 3009
rect 333238 3000 333244 3052
rect 333296 3040 333302 3052
rect 348050 3040 348056 3052
rect 333296 3012 348056 3040
rect 333296 3000 333302 3012
rect 348050 3000 348056 3012
rect 348108 3000 348114 3052
rect 349065 3043 349123 3049
rect 349065 3009 349077 3043
rect 349111 3040 349123 3043
rect 349709 3043 349767 3049
rect 349709 3040 349721 3043
rect 349111 3012 349721 3040
rect 349111 3009 349123 3012
rect 349065 3003 349123 3009
rect 349709 3009 349721 3012
rect 349755 3009 349767 3043
rect 349709 3003 349767 3009
rect 349801 3043 349859 3049
rect 349801 3009 349813 3043
rect 349847 3040 349859 3043
rect 362310 3040 362316 3052
rect 349847 3012 362316 3040
rect 349847 3009 349859 3012
rect 349801 3003 349859 3009
rect 362310 3000 362316 3012
rect 362368 3000 362374 3052
rect 362402 3000 362408 3052
rect 362460 3040 362466 3052
rect 369121 3043 369179 3049
rect 369121 3040 369133 3043
rect 362460 3012 369133 3040
rect 362460 3000 362466 3012
rect 369121 3009 369133 3012
rect 369167 3009 369179 3043
rect 369121 3003 369179 3009
rect 369213 3043 369271 3049
rect 369213 3009 369225 3043
rect 369259 3040 369271 3043
rect 397730 3040 397736 3052
rect 369259 3012 397736 3040
rect 369259 3009 369271 3012
rect 369213 3003 369271 3009
rect 397730 3000 397736 3012
rect 397788 3000 397794 3052
rect 186501 2975 186559 2981
rect 186501 2941 186513 2975
rect 186547 2972 186559 2975
rect 233418 2972 233424 2984
rect 186547 2944 233424 2972
rect 186547 2941 186559 2944
rect 186501 2935 186559 2941
rect 233418 2932 233424 2944
rect 233476 2932 233482 2984
rect 315390 2932 315396 2984
rect 315448 2972 315454 2984
rect 320729 2975 320787 2981
rect 320729 2972 320741 2975
rect 315448 2944 320741 2972
rect 315448 2932 315454 2944
rect 320729 2941 320741 2944
rect 320775 2941 320787 2975
rect 320729 2935 320787 2941
rect 320821 2975 320879 2981
rect 320821 2941 320833 2975
rect 320867 2972 320879 2975
rect 454494 2972 454500 2984
rect 320867 2944 454500 2972
rect 320867 2941 320879 2944
rect 320821 2935 320879 2941
rect 454494 2932 454500 2944
rect 454552 2932 454558 2984
rect 194321 2907 194379 2913
rect 194321 2904 194333 2907
rect 186332 2876 194333 2904
rect 194321 2873 194333 2876
rect 194367 2873 194379 2907
rect 194321 2867 194379 2873
rect 195149 2907 195207 2913
rect 195149 2873 195161 2907
rect 195195 2904 195207 2907
rect 196802 2904 196808 2916
rect 195195 2876 196808 2904
rect 195195 2873 195207 2876
rect 195149 2867 195207 2873
rect 196802 2864 196808 2876
rect 196860 2864 196866 2916
rect 196897 2907 196955 2913
rect 196897 2873 196909 2907
rect 196943 2904 196955 2907
rect 323302 2904 323308 2916
rect 196943 2876 323308 2904
rect 196943 2873 196955 2876
rect 196897 2867 196955 2873
rect 323302 2864 323308 2876
rect 323360 2864 323366 2916
rect 323670 2864 323676 2916
rect 323728 2904 323734 2916
rect 333882 2904 333888 2916
rect 323728 2876 333888 2904
rect 323728 2864 323734 2876
rect 333882 2864 333888 2876
rect 333940 2864 333946 2916
rect 340966 2904 340972 2916
rect 334084 2876 340972 2904
rect 138842 2836 138848 2848
rect 99208 2740 100248 2768
rect 100312 2808 138848 2836
rect 100312 2700 100340 2808
rect 138842 2796 138848 2808
rect 138900 2796 138906 2848
rect 159358 2796 159364 2848
rect 159416 2836 159422 2848
rect 171962 2836 171968 2848
rect 159416 2808 171968 2836
rect 159416 2796 159422 2808
rect 171962 2796 171968 2808
rect 172020 2796 172026 2848
rect 173250 2796 173256 2848
rect 173308 2836 173314 2848
rect 178129 2839 178187 2845
rect 178129 2836 178141 2839
rect 173308 2808 178141 2836
rect 173308 2796 173314 2808
rect 178129 2805 178141 2808
rect 178175 2805 178187 2839
rect 178129 2799 178187 2805
rect 178221 2839 178279 2845
rect 178221 2805 178233 2839
rect 178267 2836 178279 2839
rect 229830 2836 229836 2848
rect 178267 2808 229836 2836
rect 178267 2805 178279 2808
rect 178221 2799 178279 2805
rect 229830 2796 229836 2808
rect 229888 2796 229894 2848
rect 312538 2796 312544 2848
rect 312596 2836 312602 2848
rect 320821 2839 320879 2845
rect 320821 2836 320833 2839
rect 312596 2808 320833 2836
rect 312596 2796 312602 2808
rect 320821 2805 320833 2808
rect 320867 2805 320879 2839
rect 333977 2839 334035 2845
rect 333977 2836 333989 2839
rect 320821 2799 320879 2805
rect 320928 2808 333989 2836
rect 320637 2771 320695 2777
rect 320637 2737 320649 2771
rect 320683 2768 320695 2771
rect 320928 2768 320956 2808
rect 333977 2805 333989 2808
rect 334023 2805 334035 2839
rect 333977 2799 334035 2805
rect 320683 2740 320956 2768
rect 320683 2737 320695 2740
rect 320637 2731 320695 2737
rect 324314 2728 324320 2780
rect 324372 2768 324378 2780
rect 325602 2768 325608 2780
rect 324372 2740 325608 2768
rect 324372 2728 324378 2740
rect 325602 2728 325608 2740
rect 325660 2728 325666 2780
rect 333149 2771 333207 2777
rect 333149 2737 333161 2771
rect 333195 2768 333207 2771
rect 334084 2768 334112 2876
rect 340966 2864 340972 2876
rect 341024 2864 341030 2916
rect 341518 2864 341524 2916
rect 341576 2904 341582 2916
rect 344649 2907 344707 2913
rect 344649 2904 344661 2907
rect 341576 2876 344661 2904
rect 341576 2864 341582 2876
rect 344649 2873 344661 2876
rect 344695 2873 344707 2907
rect 344649 2867 344707 2873
rect 344741 2907 344799 2913
rect 344741 2873 344753 2907
rect 344787 2904 344799 2907
rect 355226 2904 355232 2916
rect 344787 2876 355232 2904
rect 344787 2873 344799 2876
rect 344741 2867 344799 2873
rect 355226 2864 355232 2876
rect 355284 2864 355290 2916
rect 355318 2864 355324 2916
rect 355376 2904 355382 2916
rect 355873 2907 355931 2913
rect 355376 2876 355824 2904
rect 355376 2864 355382 2876
rect 334161 2839 334219 2845
rect 334161 2805 334173 2839
rect 334207 2836 334219 2839
rect 355689 2839 355747 2845
rect 355689 2836 355701 2839
rect 334207 2808 355701 2836
rect 334207 2805 334219 2808
rect 334161 2799 334219 2805
rect 355689 2805 355701 2808
rect 355735 2805 355747 2839
rect 355689 2799 355747 2805
rect 333195 2740 334112 2768
rect 355796 2768 355824 2876
rect 355873 2873 355885 2907
rect 355919 2904 355931 2907
rect 358722 2904 358728 2916
rect 355919 2876 358728 2904
rect 355919 2873 355931 2876
rect 355873 2867 355931 2873
rect 358722 2864 358728 2876
rect 358780 2864 358786 2916
rect 390646 2904 390652 2916
rect 358924 2876 390652 2904
rect 355965 2839 356023 2845
rect 355965 2805 355977 2839
rect 356011 2836 356023 2839
rect 358817 2839 358875 2845
rect 358817 2836 358829 2839
rect 356011 2808 358829 2836
rect 356011 2805 356023 2808
rect 355965 2799 356023 2805
rect 358817 2805 358829 2808
rect 358863 2805 358875 2839
rect 358817 2799 358875 2805
rect 358924 2768 358952 2876
rect 390646 2864 390652 2876
rect 390704 2864 390710 2916
rect 359001 2839 359059 2845
rect 359001 2805 359013 2839
rect 359047 2836 359059 2839
rect 440326 2836 440332 2848
rect 359047 2808 440332 2836
rect 359047 2805 359059 2808
rect 359001 2799 359059 2805
rect 440326 2796 440332 2808
rect 440384 2796 440390 2848
rect 355796 2740 358952 2768
rect 333195 2737 333207 2740
rect 333149 2731 333207 2737
rect 99116 2672 100340 2700
<< via1 >>
rect 24308 700952 24360 701004
rect 196348 700952 196400 701004
rect 8116 700884 8168 700936
rect 188988 700884 189040 700936
rect 164148 700816 164200 700868
rect 348792 700816 348844 700868
rect 40500 700748 40552 700800
rect 227720 700748 227772 700800
rect 154488 700680 154540 700732
rect 397460 700680 397512 700732
rect 157248 700612 157300 700664
rect 413652 700612 413704 700664
rect 148324 700544 148376 700596
rect 462320 700544 462372 700596
rect 150348 700476 150400 700528
rect 478512 700476 478564 700528
rect 144828 700408 144880 700460
rect 494796 700408 494848 700460
rect 140688 700340 140740 700392
rect 527180 700340 527232 700392
rect 89168 700272 89220 700324
rect 98644 700272 98696 700324
rect 137100 700272 137152 700324
rect 559656 700272 559708 700324
rect 162768 700204 162820 700256
rect 332508 700204 332560 700256
rect 72976 700136 73028 700188
rect 188344 700136 188396 700188
rect 188436 700136 188488 700188
rect 218980 700136 219032 700188
rect 172428 700068 172480 700120
rect 283840 700068 283892 700120
rect 169668 700000 169720 700052
rect 267648 700000 267700 700052
rect 105452 699932 105504 699984
rect 187976 699932 188028 699984
rect 173808 699864 173860 699916
rect 235172 699864 235224 699916
rect 175924 699796 175976 699848
rect 202788 699796 202840 699848
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 251456 699660 251508 699712
rect 252468 699660 252520 699712
rect 381176 699660 381228 699712
rect 382188 699660 382240 699712
rect 133604 696940 133656 696992
rect 580172 696940 580224 696992
rect 410616 692792 410668 692844
rect 463332 692792 463384 692844
rect 3516 670692 3568 670744
rect 188528 670692 188580 670744
rect 542360 670352 542412 670404
rect 542360 668380 542412 668432
rect 2872 657500 2924 657552
rect 197820 657500 197872 657552
rect 429200 648320 429252 648372
rect 429200 648048 429252 648100
rect 227720 647096 227772 647148
rect 226156 646348 226208 646400
rect 226156 646051 226208 646060
rect 4804 645872 4856 645924
rect 32036 645872 32088 645924
rect 188528 645872 188580 645924
rect 198188 645872 198240 645924
rect 226156 646017 226165 646051
rect 226165 646017 226199 646051
rect 226199 646017 226208 646051
rect 226156 646008 226208 646017
rect 580356 645804 580408 645856
rect 188068 645600 188120 645652
rect 188344 645643 188396 645652
rect 188344 645609 188353 645643
rect 188353 645609 188387 645643
rect 188387 645609 188396 645643
rect 188344 645600 188396 645609
rect 188436 645600 188488 645652
rect 187976 645328 188028 645380
rect 196348 645575 196400 645584
rect 196348 645541 196357 645575
rect 196357 645541 196391 645575
rect 196391 645541 196400 645575
rect 196348 645532 196400 645541
rect 188436 645328 188488 645380
rect 197912 645124 197964 645176
rect 471888 644852 471940 644904
rect 459560 644444 459612 644496
rect 124772 643288 124824 643340
rect 128912 643288 128964 643340
rect 129280 643288 129332 643340
rect 132776 643288 132828 643340
rect 133144 643288 133196 643340
rect 136640 643288 136692 643340
rect 137008 643288 137060 643340
rect 579620 643288 579672 643340
rect 443644 643195 443696 643204
rect 443644 643161 443653 643195
rect 443653 643161 443687 643195
rect 443687 643161 443696 643195
rect 443644 643152 443696 643161
rect 196900 642336 196952 642388
rect 199568 640976 199620 641028
rect 214564 640976 214616 641028
rect 196992 640704 197044 640756
rect 90824 639888 90876 639940
rect 96344 639888 96396 639940
rect 197452 639548 197504 639600
rect 233884 639548 233936 639600
rect 415308 639548 415360 639600
rect 194692 639480 194744 639532
rect 194600 639412 194652 639464
rect 182916 639072 182968 639124
rect 196348 639072 196400 639124
rect 197084 639072 197136 639124
rect 184020 639004 184072 639056
rect 182548 638936 182600 638988
rect 187976 638800 188028 638852
rect 188436 638800 188488 638852
rect 188988 638800 189040 638852
rect 188988 638528 189040 638580
rect 187976 638460 188028 638512
rect 188344 638503 188396 638512
rect 188344 638469 188353 638503
rect 188353 638469 188387 638503
rect 188387 638469 188396 638503
rect 188344 638460 188396 638469
rect 188436 638460 188488 638512
rect 196256 638392 196308 638444
rect 196992 638392 197044 638444
rect 188528 638324 188580 638376
rect 214564 637848 214616 637900
rect 218888 637848 218940 637900
rect 214564 637576 214616 637628
rect 218888 637576 218940 637628
rect 218888 635944 218940 635996
rect 196256 635604 196308 635656
rect 196348 635647 196400 635656
rect 196348 635613 196357 635647
rect 196357 635613 196391 635647
rect 196391 635613 196400 635647
rect 196348 635604 196400 635613
rect 196164 635332 196216 635384
rect 196348 635171 196400 635180
rect 196348 635137 196357 635171
rect 196357 635137 196391 635171
rect 196391 635137 196400 635171
rect 196348 635128 196400 635137
rect 90824 634924 90876 634976
rect 96988 634924 97040 634976
rect 120264 634856 120316 634908
rect 126796 634856 126848 634908
rect 189264 634856 189316 634908
rect 191564 634856 191616 634908
rect 198464 634015 198516 634024
rect 198464 633981 198473 634015
rect 198473 633981 198507 634015
rect 198507 633981 198516 634015
rect 198464 633972 198516 633981
rect 199568 634015 199620 634024
rect 199568 633981 199577 634015
rect 199577 633981 199611 634015
rect 199611 633981 199620 634015
rect 199568 633972 199620 633981
rect 202207 633700 202259 633752
rect 3240 633360 3292 633412
rect 97908 633360 97960 633412
rect 214564 632748 214616 632800
rect 99748 632680 99800 632732
rect 126888 632680 126940 632732
rect 198464 632519 198516 632528
rect 198464 632485 198473 632519
rect 198473 632485 198507 632519
rect 198507 632485 198516 632519
rect 198464 632476 198516 632485
rect 199568 632519 199620 632528
rect 199568 632485 199577 632519
rect 199577 632485 199611 632519
rect 199611 632485 199620 632519
rect 199568 632476 199620 632485
rect 189816 632408 189868 632460
rect 191564 632408 191616 632460
rect 201960 632247 202012 632256
rect 201960 632213 201969 632247
rect 201969 632213 202003 632247
rect 202003 632213 202012 632247
rect 201960 632204 202012 632213
rect 436744 631796 436796 631848
rect 215392 631728 215444 631780
rect 128268 631388 128320 631440
rect 128912 631388 128964 631440
rect 129280 631388 129332 631440
rect 132776 631388 132828 631440
rect 133144 631388 133196 631440
rect 136640 631388 136692 631440
rect 137008 631388 137060 631440
rect 191564 631388 191616 631440
rect 192944 631116 192996 631168
rect 506664 631184 506716 631236
rect 579804 631320 579856 631372
rect 221096 630640 221148 630692
rect 496084 630776 496136 630828
rect 218888 629076 218940 629128
rect 414664 628940 414716 628992
rect 198464 628260 198516 628312
rect 199568 628260 199620 628312
rect 201960 628192 202012 628244
rect 210240 628192 210292 628244
rect 197360 627963 197412 627972
rect 197360 627929 197369 627963
rect 197369 627929 197403 627963
rect 197403 627929 197412 627963
rect 197360 627920 197412 627929
rect 197820 627920 197872 627972
rect 199568 627920 199620 627972
rect 214564 628192 214616 628244
rect 210976 627988 211028 628040
rect 201960 627852 202012 627904
rect 218888 627759 218940 627768
rect 218888 627725 218897 627759
rect 218897 627725 218931 627759
rect 218931 627725 218940 627759
rect 218888 627716 218940 627725
rect 214564 626764 214616 626816
rect 214564 626560 214616 626612
rect 187976 624656 188028 624708
rect 188344 624656 188396 624708
rect 188436 624656 188488 624708
rect 188528 624656 188580 624708
rect 188988 624656 189040 624708
rect 187976 624316 188028 624368
rect 188344 624316 188396 624368
rect 188436 624316 188488 624368
rect 188528 624316 188580 624368
rect 188988 624316 189040 624368
rect 542360 623024 542412 623076
rect 128268 621868 128320 621920
rect 128268 621324 128320 621376
rect 3608 620984 3660 621036
rect 31760 620984 31812 621036
rect 218888 620007 218940 620016
rect 218888 619973 218897 620007
rect 218897 619973 218931 620007
rect 218931 619973 218940 620007
rect 218888 619964 218940 619973
rect 542452 619828 542504 619880
rect 3516 619624 3568 619676
rect 31760 619624 31812 619676
rect 382188 619624 382240 619676
rect 3424 618536 3476 618588
rect 79232 618536 79284 618588
rect 79784 618536 79836 618588
rect 137100 618919 137152 618928
rect 137100 618885 137109 618919
rect 137109 618885 137143 618919
rect 137143 618885 137152 618919
rect 137100 618876 137152 618885
rect 199568 618536 199620 618588
rect 137100 618307 137152 618316
rect 137100 618273 137109 618307
rect 137109 618273 137143 618307
rect 137143 618273 137152 618307
rect 137100 618264 137152 618273
rect 124128 617992 124180 618044
rect 131488 617992 131540 618044
rect 132040 617040 132092 617092
rect 580172 617040 580224 617092
rect 160100 607112 160152 607164
rect 160928 607112 160980 607164
rect 124128 601944 124180 601996
rect 124772 601944 124824 601996
rect 128268 601944 128320 601996
rect 133604 601944 133656 601996
rect 124128 601536 124180 601588
rect 124772 601536 124824 601588
rect 128268 601536 128320 601588
rect 133604 601536 133656 601588
rect 159548 591268 159600 591320
rect 580172 591268 580224 591320
rect 3516 578212 3568 578264
rect 31852 578212 31904 578264
rect 98644 577983 98696 577992
rect 98644 577949 98653 577983
rect 98653 577949 98687 577983
rect 98687 577949 98696 577983
rect 98644 577940 98696 577949
rect 98644 577575 98696 577584
rect 98644 577541 98653 577575
rect 98653 577541 98687 577575
rect 98687 577541 98696 577575
rect 98644 577532 98696 577541
rect 139492 577464 139544 577516
rect 579988 577464 580040 577516
rect 410340 569916 410392 569968
rect 410616 569916 410668 569968
rect 579620 569916 579672 569968
rect 404268 566856 404320 566908
rect 427820 566448 427872 566500
rect 92388 558900 92440 558952
rect 391848 558900 391900 558952
rect 3332 553392 3384 553444
rect 211804 553392 211856 553444
rect 99288 542376 99340 542428
rect 391388 542376 391440 542428
rect 391756 542376 391808 542428
rect 3332 540880 3384 540932
rect 31760 540880 31812 540932
rect 111708 536800 111760 536852
rect 580172 536800 580224 536852
rect 417700 534012 417752 534064
rect 580356 534012 580408 534064
rect 401600 533944 401652 533996
rect 402060 533944 402112 533996
rect 542360 533944 542412 533996
rect 143448 533400 143500 533452
rect 401600 533400 401652 533452
rect 115848 533332 115900 533384
rect 417700 533332 417752 533384
rect 3332 527144 3384 527196
rect 223580 527144 223632 527196
rect 114468 524424 114520 524476
rect 580172 524424 580224 524476
rect 3332 515380 3384 515432
rect 197360 515380 197412 515432
rect 197360 514768 197412 514820
rect 198004 514768 198056 514820
rect 108948 510620 109000 510672
rect 580172 510620 580224 510672
rect 2872 500964 2924 501016
rect 218704 500964 218756 501016
rect 104808 484372 104860 484424
rect 579988 484372 580040 484424
rect 3056 474716 3108 474768
rect 230480 474716 230532 474768
rect 106188 470568 106240 470620
rect 580172 470568 580224 470620
rect 3332 462340 3384 462392
rect 200764 462340 200816 462392
rect 100760 457444 100812 457496
rect 579620 457444 579672 457496
rect 3332 448536 3384 448588
rect 226984 448536 227036 448588
rect 96528 430584 96580 430636
rect 579896 430584 579948 430636
rect 3516 422288 3568 422340
rect 237380 422288 237432 422340
rect 391756 419432 391808 419484
rect 580172 419432 580224 419484
rect 2872 409844 2924 409896
rect 221464 409844 221516 409896
rect 95148 404336 95200 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 233884 397468 233936 397520
rect 89628 378156 89680 378208
rect 580172 378156 580224 378208
rect 3516 371220 3568 371272
rect 245660 371220 245712 371272
rect 391848 365644 391900 365696
rect 580172 365644 580224 365696
rect 88248 351908 88300 351960
rect 580172 351908 580224 351960
rect 82544 324300 82596 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 252744 318792 252796 318844
rect 171048 314236 171100 314288
rect 180892 314236 180944 314288
rect 98644 314168 98696 314220
rect 192576 314168 192628 314220
rect 198004 314168 198056 314220
rect 228732 314168 228784 314220
rect 166816 314100 166868 314152
rect 299480 314100 299532 314152
rect 3424 314032 3476 314084
rect 216680 314032 216732 314084
rect 135076 313964 135128 314016
rect 443644 313964 443696 314016
rect 130660 313896 130712 313948
rect 580264 313896 580316 313948
rect 188344 313216 188396 313268
rect 190460 313216 190512 313268
rect 196348 313216 196400 313268
rect 200120 313216 200172 313268
rect 204904 313216 204956 313268
rect 211896 313216 211948 313268
rect 218888 313216 218940 313268
rect 221556 313216 221608 313268
rect 233884 313216 233936 313268
rect 240784 313216 240836 313268
rect 154396 313148 154448 313200
rect 142712 313080 142764 313132
rect 143448 313080 143500 313132
rect 147496 313080 147548 313132
rect 148324 313080 148376 313132
rect 149888 313080 149940 313132
rect 150348 313080 150400 313132
rect 152280 313080 152332 313132
rect 153108 313080 153160 313132
rect 159548 313080 159600 313132
rect 160008 313080 160060 313132
rect 161940 313148 161992 313200
rect 162768 313148 162820 313200
rect 169208 313148 169260 313200
rect 169668 313148 169720 313200
rect 171600 313148 171652 313200
rect 172428 313148 172480 313200
rect 178776 313148 178828 313200
rect 188436 313148 188488 313200
rect 197452 313148 197504 313200
rect 197820 313148 197872 313200
rect 204628 313148 204680 313200
rect 218704 313148 218756 313200
rect 226340 313148 226392 313200
rect 226984 313148 227036 313200
rect 233516 313148 233568 313200
rect 185400 313080 185452 313132
rect 188528 313080 188580 313132
rect 207020 313080 207072 313132
rect 211804 313080 211856 313132
rect 219072 313080 219124 313132
rect 221464 313080 221516 313132
rect 243176 313080 243228 313132
rect 87328 313012 87380 313064
rect 88248 313012 88300 313064
rect 94504 313012 94556 313064
rect 95148 313012 95200 313064
rect 104164 313012 104216 313064
rect 104808 313012 104860 313064
rect 113824 313012 113876 313064
rect 114468 313012 114520 313064
rect 123392 313012 123444 313064
rect 124128 313012 124180 313064
rect 124772 313012 124824 313064
rect 125232 313012 125284 313064
rect 133052 313012 133104 313064
rect 133604 313012 133656 313064
rect 137928 313012 137980 313064
rect 183008 313012 183060 313064
rect 188988 313012 189040 313064
rect 195704 313012 195756 313064
rect 196256 313012 196308 313064
rect 200764 313012 200816 313064
rect 236000 313012 236052 313064
rect 77668 312944 77720 312996
rect 303436 312944 303488 312996
rect 75276 312876 75328 312928
rect 303528 312876 303580 312928
rect 3976 312808 4028 312860
rect 247960 312808 248012 312860
rect 3608 312740 3660 312792
rect 250444 312740 250496 312792
rect 6368 312672 6420 312724
rect 257620 312672 257672 312724
rect 5356 312604 5408 312656
rect 262496 312604 262548 312656
rect 6276 312536 6328 312588
rect 264980 312536 265032 312588
rect 3332 312468 3384 312520
rect 272064 312468 272116 312520
rect 3884 312400 3936 312452
rect 276940 312400 276992 312452
rect 6184 312332 6236 312384
rect 279332 312332 279384 312384
rect 5172 312264 5224 312316
rect 281724 312264 281776 312316
rect 5080 312196 5132 312248
rect 284300 312196 284352 312248
rect 3792 312128 3844 312180
rect 286508 312128 286560 312180
rect 4988 312060 5040 312112
rect 288900 312060 288952 312112
rect 4896 311992 4948 312044
rect 291384 311992 291436 312044
rect 3700 311924 3752 311976
rect 293960 311924 294012 311976
rect 84936 311856 84988 311908
rect 580172 311856 580224 311908
rect 31760 310496 31812 310548
rect 302884 310496 302936 310548
rect 79968 310428 80020 310480
rect 304632 310428 304684 310480
rect 65616 310360 65668 310412
rect 60648 310335 60700 310344
rect 60648 310301 60657 310335
rect 60657 310301 60691 310335
rect 60691 310301 60700 310335
rect 60648 310292 60700 310301
rect 63224 310335 63276 310344
rect 63224 310301 63233 310335
rect 63233 310301 63267 310335
rect 63267 310301 63276 310335
rect 63224 310292 63276 310301
rect 70308 310335 70360 310344
rect 70308 310301 70317 310335
rect 70317 310301 70351 310335
rect 70351 310301 70360 310335
rect 70308 310292 70360 310301
rect 72884 310360 72936 310412
rect 304540 310360 304592 310412
rect 303344 310292 303396 310344
rect 55956 310267 56008 310276
rect 55956 310233 55965 310267
rect 55965 310233 55999 310267
rect 55999 310233 56008 310267
rect 55956 310224 56008 310233
rect 58440 310224 58492 310276
rect 303160 310224 303212 310276
rect 39120 310199 39172 310208
rect 39120 310165 39129 310199
rect 39129 310165 39163 310199
rect 39163 310165 39172 310199
rect 39120 310156 39172 310165
rect 41328 310199 41380 310208
rect 41328 310165 41337 310199
rect 41337 310165 41371 310199
rect 41371 310165 41380 310199
rect 41328 310156 41380 310165
rect 46388 310199 46440 310208
rect 46388 310165 46397 310199
rect 46397 310165 46431 310199
rect 46431 310165 46440 310199
rect 46388 310156 46440 310165
rect 48780 310199 48832 310208
rect 48780 310165 48789 310199
rect 48789 310165 48823 310199
rect 48823 310165 48832 310199
rect 48780 310156 48832 310165
rect 53564 310156 53616 310208
rect 304356 310156 304408 310208
rect 4712 310088 4764 310140
rect 255320 310088 255372 310140
rect 5448 310020 5500 310072
rect 260012 310020 260064 310072
rect 5264 309952 5316 310004
rect 267280 309952 267332 310004
rect 269672 309995 269724 310004
rect 269672 309961 269681 309995
rect 269681 309961 269715 309995
rect 269715 309961 269724 309995
rect 269672 309952 269724 309961
rect 274640 309995 274692 310004
rect 274640 309961 274649 309995
rect 274649 309961 274683 309995
rect 274683 309961 274692 309995
rect 274640 309952 274692 309961
rect 296168 309995 296220 310004
rect 296168 309961 296177 309995
rect 296177 309961 296211 309995
rect 296211 309961 296220 309995
rect 296168 309952 296220 309961
rect 304264 310020 304316 310072
rect 298560 309952 298612 310004
rect 4068 309816 4120 309868
rect 3976 309748 4028 309800
rect 3608 309680 3660 309732
rect 3424 309612 3476 309664
rect 580908 309544 580960 309596
rect 580724 309476 580776 309528
rect 580816 309408 580868 309460
rect 580632 309340 580684 309392
rect 580448 309272 580500 309324
rect 580540 309204 580592 309256
rect 580356 309136 580408 309188
rect 2964 306212 3016 306264
rect 6368 306212 6420 306264
rect 304632 299412 304684 299464
rect 580172 299412 580224 299464
rect 2780 293224 2832 293276
rect 4712 293224 4764 293276
rect 303528 273164 303580 273216
rect 579988 273164 580040 273216
rect 2780 267180 2832 267232
rect 5448 267180 5500 267232
rect 303436 259360 303488 259412
rect 580172 259360 580224 259412
rect 3148 255144 3200 255196
rect 6276 255144 6328 255196
rect 304540 245556 304592 245608
rect 580172 245556 580224 245608
rect 2780 241068 2832 241120
rect 5356 241068 5408 241120
rect 304448 233180 304500 233232
rect 579988 233180 580040 233232
rect 2780 214956 2832 215008
rect 5264 214956 5316 215008
rect 303344 206932 303396 206984
rect 580172 206932 580224 206984
rect 303160 166948 303212 167000
rect 579620 166948 579672 167000
rect 304356 153144 304408 153196
rect 579804 153144 579856 153196
rect 3148 150220 3200 150272
rect 6184 150220 6236 150272
rect 303252 126896 303304 126948
rect 579712 126896 579764 126948
rect 2780 123836 2832 123888
rect 4804 123836 4856 123888
rect 2780 111460 2832 111512
rect 5172 111460 5224 111512
rect 303068 86912 303120 86964
rect 579620 86912 579672 86964
rect 2780 85144 2832 85196
rect 5080 85144 5132 85196
rect 304264 73108 304316 73160
rect 580172 73108 580224 73160
rect 2780 71612 2832 71664
rect 4988 71612 5040 71664
rect 302976 46860 303028 46912
rect 580172 46860 580224 46912
rect 2780 45500 2832 45552
rect 4896 45500 4948 45552
rect 302884 33056 302936 33108
rect 580172 33056 580224 33108
rect 250812 31764 250864 31816
rect 251088 31764 251140 31816
rect 261944 31764 261996 31816
rect 262128 31764 262180 31816
rect 264704 31764 264756 31816
rect 264888 31764 264940 31816
rect 20536 31696 20588 31748
rect 37372 31696 37424 31748
rect 41328 31696 41380 31748
rect 46940 31696 46992 31748
rect 88156 31696 88208 31748
rect 127164 31696 127216 31748
rect 19248 31628 19300 31680
rect 36268 31628 36320 31680
rect 44088 31628 44140 31680
rect 47952 31628 48004 31680
rect 68836 31628 68888 31680
rect 16488 31560 16540 31612
rect 35164 31560 35216 31612
rect 42708 31560 42760 31612
rect 47400 31560 47452 31612
rect 83188 31628 83240 31680
rect 90272 31628 90324 31680
rect 90364 31628 90416 31680
rect 94504 31628 94556 31680
rect 108948 31628 109000 31680
rect 159364 31628 159416 31680
rect 162216 31628 162268 31680
rect 200764 31696 200816 31748
rect 215668 31696 215720 31748
rect 358084 31696 358136 31748
rect 202328 31628 202380 31680
rect 344284 31628 344336 31680
rect 85764 31560 85816 31612
rect 93676 31560 93728 31612
rect 95884 31560 95936 31612
rect 157984 31560 158036 31612
rect 188988 31560 189040 31612
rect 330484 31560 330536 31612
rect 13728 31492 13780 31544
rect 34060 31492 34112 31544
rect 72608 31492 72660 31544
rect 87512 31492 87564 31544
rect 104348 31492 104400 31544
rect 155224 31492 155276 31544
rect 166908 31492 166960 31544
rect 208952 31492 209004 31544
rect 15108 31424 15160 31476
rect 34612 31424 34664 31476
rect 38568 31424 38620 31476
rect 45744 31424 45796 31476
rect 86500 31424 86552 31476
rect 101404 31424 101456 31476
rect 106004 31424 106056 31476
rect 156604 31424 156656 31476
rect 168932 31424 168984 31476
rect 213184 31424 213236 31476
rect 219072 31424 219124 31476
rect 362224 31492 362276 31544
rect 237932 31424 237984 31476
rect 238668 31424 238720 31476
rect 376024 31424 376076 31476
rect 10968 31356 11020 31408
rect 32404 31356 32456 31408
rect 70952 31356 71004 31408
rect 88984 31356 89036 31408
rect 107568 31356 107620 31408
rect 170404 31356 170456 31408
rect 225696 31356 225748 31408
rect 369124 31356 369176 31408
rect 12348 31288 12400 31340
rect 33140 31288 33192 31340
rect 34428 31288 34480 31340
rect 43536 31288 43588 31340
rect 84844 31288 84896 31340
rect 105544 31288 105596 31340
rect 119344 31288 119396 31340
rect 173164 31288 173216 31340
rect 212356 31288 212408 31340
rect 355324 31288 355376 31340
rect 9588 31220 9640 31272
rect 31852 31220 31904 31272
rect 35808 31220 35860 31272
rect 44180 31220 44232 31272
rect 45468 31220 45520 31272
rect 48504 31220 48556 31272
rect 77024 31220 77076 31272
rect 102324 31220 102376 31272
rect 114376 31220 114428 31272
rect 167644 31220 167696 31272
rect 205548 31220 205600 31272
rect 348424 31220 348476 31272
rect 6828 31152 6880 31204
rect 30748 31152 30800 31204
rect 33048 31152 33100 31204
rect 42984 31152 43036 31204
rect 78588 31152 78640 31204
rect 112628 31152 112680 31204
rect 166264 31152 166316 31204
rect 198648 31152 198700 31204
rect 341524 31152 341576 31204
rect 4068 31084 4120 31136
rect 29644 31084 29696 31136
rect 30288 31084 30340 31136
rect 41880 31084 41932 31136
rect 45376 31084 45428 31136
rect 49148 31084 49200 31136
rect 82084 31084 82136 31136
rect 108304 31084 108356 31136
rect 115848 31084 115900 31136
rect 169024 31084 169076 31136
rect 222016 31084 222068 31136
rect 366364 31084 366416 31136
rect 5448 31016 5500 31068
rect 30380 31016 30432 31068
rect 31668 31016 31720 31068
rect 42432 31016 42484 31068
rect 67548 31016 67600 31068
rect 83004 31016 83056 31068
rect 85396 31016 85448 31068
rect 119344 31016 119396 31068
rect 121000 31016 121052 31068
rect 175924 31016 175976 31068
rect 180524 31016 180576 31068
rect 185492 31016 185544 31068
rect 228916 31016 228968 31068
rect 373264 31016 373316 31068
rect 23388 30948 23440 31000
rect 38660 30948 38712 31000
rect 39948 30948 40000 31000
rect 46296 30948 46348 31000
rect 104164 30948 104216 31000
rect 110972 30948 111024 31000
rect 160744 30948 160796 31000
rect 195612 30948 195664 31000
rect 337384 30948 337436 31000
rect 20628 30880 20680 30932
rect 36820 30880 36872 30932
rect 92296 30880 92348 30932
rect 135444 30880 135496 30932
rect 22008 30812 22060 30864
rect 37924 30812 37976 30864
rect 90916 30812 90968 30864
rect 132500 30812 132552 30864
rect 137928 30812 137980 30864
rect 179972 30880 180024 30932
rect 192300 30880 192352 30932
rect 24768 30744 24820 30796
rect 39120 30744 39172 30796
rect 102048 30744 102100 30796
rect 142804 30744 142856 30796
rect 28908 30676 28960 30728
rect 41420 30676 41472 30728
rect 89628 30676 89680 30728
rect 129740 30676 129792 30728
rect 136548 30676 136600 30728
rect 177396 30812 177448 30864
rect 185584 30812 185636 30864
rect 172244 30744 172296 30796
rect 180064 30744 180116 30796
rect 180708 30744 180760 30796
rect 181168 30744 181220 30796
rect 182088 30744 182140 30796
rect 183928 30744 183980 30796
rect 184848 30744 184900 30796
rect 187332 30812 187384 30864
rect 187608 30812 187660 30864
rect 189540 30812 189592 30864
rect 190276 30812 190328 30864
rect 191196 30812 191248 30864
rect 191748 30812 191800 30864
rect 193956 30812 194008 30864
rect 194508 30812 194560 30864
rect 204904 30880 204956 30932
rect 209044 30880 209096 30932
rect 351184 30880 351236 30932
rect 333244 30812 333296 30864
rect 323676 30744 323728 30796
rect 175188 30676 175240 30728
rect 301504 30676 301556 30728
rect 27528 30608 27580 30660
rect 40224 30608 40276 30660
rect 117688 30608 117740 30660
rect 128268 30608 128320 30660
rect 177212 30608 177264 30660
rect 178960 30608 179012 30660
rect 26148 30540 26200 30592
rect 39672 30540 39724 30592
rect 139952 30540 140004 30592
rect 181444 30540 181496 30592
rect 182824 30540 182876 30592
rect 183468 30540 183520 30592
rect 184480 30540 184532 30592
rect 184756 30540 184808 30592
rect 186688 30540 186740 30592
rect 187424 30540 187476 30592
rect 188436 30540 188488 30592
rect 188988 30540 189040 30592
rect 192852 30540 192904 30592
rect 193128 30540 193180 30592
rect 195060 30540 195112 30592
rect 195796 30540 195848 30592
rect 196716 30540 196768 30592
rect 197176 30540 197228 30592
rect 197912 30540 197964 30592
rect 198648 30540 198700 30592
rect 199568 30540 199620 30592
rect 200028 30540 200080 30592
rect 203432 30540 203484 30592
rect 204076 30540 204128 30592
rect 210700 30540 210752 30592
rect 211068 30540 211120 30592
rect 224040 30540 224092 30592
rect 224868 30540 224920 30592
rect 227352 30540 227404 30592
rect 227628 30540 227680 30592
rect 232412 30540 232464 30592
rect 28816 30472 28868 30524
rect 40776 30472 40828 30524
rect 49608 30472 49660 30524
rect 51080 30472 51132 30524
rect 171692 30472 171744 30524
rect 172428 30472 172480 30524
rect 173348 30472 173400 30524
rect 173808 30472 173860 30524
rect 174452 30472 174504 30524
rect 175004 30472 175056 30524
rect 177304 30472 177356 30524
rect 177856 30472 177908 30524
rect 178408 30472 178460 30524
rect 179236 30472 179288 30524
rect 244924 30472 244976 30524
rect 37096 30404 37148 30456
rect 45192 30404 45244 30456
rect 46848 30404 46900 30456
rect 49700 30404 49752 30456
rect 56968 30404 57020 30456
rect 57888 30404 57940 30456
rect 59728 30404 59780 30456
rect 60648 30404 60700 30456
rect 79232 30404 79284 30456
rect 79876 30404 79928 30456
rect 88708 30404 88760 30456
rect 93124 30404 93176 30456
rect 97080 30404 97132 30456
rect 97908 30404 97960 30456
rect 100300 30404 100352 30456
rect 100668 30404 100720 30456
rect 123852 30404 123904 30456
rect 124128 30404 124180 30456
rect 128820 30404 128872 30456
rect 129648 30404 129700 30456
rect 132132 30404 132184 30456
rect 132408 30404 132460 30456
rect 149428 30404 149480 30456
rect 150348 30404 150400 30456
rect 152740 30404 152792 30456
rect 153108 30404 153160 30456
rect 158352 30404 158404 30456
rect 158628 30404 158680 30456
rect 161112 30404 161164 30456
rect 161388 30404 161440 30456
rect 163320 30404 163372 30456
rect 164148 30404 164200 30456
rect 165436 30404 165488 30456
rect 37188 30336 37240 30388
rect 44640 30336 44692 30388
rect 48228 30336 48280 30388
rect 50252 30336 50304 30388
rect 52460 30336 52512 30388
rect 53012 30336 53064 30388
rect 55864 30336 55916 30388
rect 56508 30336 56560 30388
rect 57520 30336 57572 30388
rect 57796 30336 57848 30388
rect 58624 30336 58676 30388
rect 59268 30336 59320 30388
rect 60372 30336 60424 30388
rect 60556 30336 60608 30388
rect 61476 30336 61528 30388
rect 61936 30336 61988 30388
rect 62580 30336 62632 30388
rect 63408 30336 63460 30388
rect 64236 30336 64288 30388
rect 64696 30336 64748 30388
rect 65340 30336 65392 30388
rect 65892 30336 65944 30388
rect 66996 30336 67048 30388
rect 67548 30336 67600 30388
rect 68100 30336 68152 30388
rect 68928 30336 68980 30388
rect 69756 30336 69808 30388
rect 70308 30336 70360 30388
rect 73712 30336 73764 30388
rect 74448 30336 74500 30388
rect 75368 30336 75420 30388
rect 75828 30336 75880 30388
rect 76472 30336 76524 30388
rect 77208 30336 77260 30388
rect 78128 30336 78180 30388
rect 78588 30336 78640 30388
rect 79692 30336 79744 30388
rect 79968 30336 80020 30388
rect 85948 30336 86000 30388
rect 86776 30336 86828 30388
rect 87604 30336 87656 30388
rect 88248 30336 88300 30388
rect 91468 30336 91520 30388
rect 92296 30336 92348 30388
rect 93216 30336 93268 30388
rect 93768 30336 93820 30388
rect 94320 30336 94372 30388
rect 94872 30336 94924 30388
rect 95976 30336 96028 30388
rect 96528 30336 96580 30388
rect 97632 30336 97684 30388
rect 97816 30336 97868 30388
rect 98736 30336 98788 30388
rect 99288 30336 99340 30388
rect 99840 30336 99892 30388
rect 100576 30336 100628 30388
rect 101496 30336 101548 30388
rect 102048 30336 102100 30388
rect 102692 30336 102744 30388
rect 103244 30336 103296 30388
rect 105452 30336 105504 30388
rect 106188 30336 106240 30388
rect 107108 30336 107160 30388
rect 107568 30336 107620 30388
rect 108212 30336 108264 30388
rect 108948 30336 109000 30388
rect 113824 30336 113876 30388
rect 114468 30336 114520 30388
rect 114928 30336 114980 30388
rect 115480 30336 115532 30388
rect 116584 30336 116636 30388
rect 117136 30336 117188 30388
rect 120448 30336 120500 30388
rect 121368 30336 121420 30388
rect 122104 30336 122156 30388
rect 122748 30336 122800 30388
rect 123208 30336 123260 30388
rect 123944 30336 123996 30388
rect 124956 30336 125008 30388
rect 125416 30336 125468 30388
rect 126060 30336 126112 30388
rect 126796 30336 126848 30388
rect 127716 30336 127768 30388
rect 128268 30336 128320 30388
rect 129372 30336 129424 30388
rect 129556 30336 129608 30388
rect 130476 30336 130528 30388
rect 131028 30336 131080 30388
rect 131580 30336 131632 30388
rect 132224 30336 132276 30388
rect 133236 30336 133288 30388
rect 133696 30336 133748 30388
rect 134432 30336 134484 30388
rect 135076 30336 135128 30388
rect 136088 30336 136140 30388
rect 136548 30336 136600 30388
rect 137192 30336 137244 30388
rect 137928 30336 137980 30388
rect 140504 30336 140556 30388
rect 140688 30336 140740 30388
rect 141608 30336 141660 30388
rect 142068 30336 142120 30388
rect 142712 30336 142764 30388
rect 143264 30336 143316 30388
rect 143448 30336 143500 30388
rect 144368 30336 144420 30388
rect 144828 30336 144880 30388
rect 145564 30336 145616 30388
rect 146116 30336 146168 30388
rect 146668 30336 146720 30388
rect 147496 30336 147548 30388
rect 148324 30336 148376 30388
rect 148968 30336 149020 30388
rect 149980 30336 150032 30388
rect 150256 30336 150308 30388
rect 151084 30336 151136 30388
rect 151728 30336 151780 30388
rect 152188 30336 152240 30388
rect 152924 30336 152976 30388
rect 153844 30336 153896 30388
rect 154396 30336 154448 30388
rect 154948 30336 155000 30388
rect 155776 30336 155828 30388
rect 156696 30336 156748 30388
rect 157248 30336 157300 30388
rect 157800 30336 157852 30388
rect 158444 30336 158496 30388
rect 159456 30336 159508 30388
rect 159916 30336 159968 30388
rect 160560 30336 160612 30388
rect 161204 30336 161256 30388
rect 163872 30336 163924 30388
rect 164056 30336 164108 30388
rect 164976 30336 165028 30388
rect 165528 30336 165580 30388
rect 166172 30336 166224 30388
rect 166908 30336 166960 30388
rect 170588 30404 170640 30456
rect 242164 30404 242216 30456
rect 242440 30404 242492 30456
rect 250168 30472 250220 30524
rect 250996 30472 251048 30524
rect 251916 30472 251968 30524
rect 252468 30472 252520 30524
rect 253020 30472 253072 30524
rect 253572 30472 253624 30524
rect 254676 30472 254728 30524
rect 255136 30472 255188 30524
rect 255780 30472 255832 30524
rect 256516 30472 256568 30524
rect 257436 30472 257488 30524
rect 257988 30472 258040 30524
rect 259092 30472 259144 30524
rect 259276 30472 259328 30524
rect 260196 30472 260248 30524
rect 260748 30472 260800 30524
rect 261392 30472 261444 30524
rect 261944 30472 261996 30524
rect 263048 30472 263100 30524
rect 263508 30472 263560 30524
rect 264152 30472 264204 30524
rect 264704 30472 264756 30524
rect 266912 30472 266964 30524
rect 267556 30472 267608 30524
rect 268568 30472 268620 30524
rect 269028 30472 269080 30524
rect 269672 30608 269724 30660
rect 270500 30608 270552 30660
rect 276296 30608 276348 30660
rect 276388 30608 276440 30660
rect 277308 30608 277360 30660
rect 279700 30608 279752 30660
rect 280068 30608 280120 30660
rect 284760 30608 284812 30660
rect 285588 30608 285640 30660
rect 288072 30608 288124 30660
rect 288348 30608 288400 30660
rect 293132 30608 293184 30660
rect 293960 30608 294012 30660
rect 301412 30608 301464 30660
rect 308404 30608 308456 30660
rect 309784 30540 309836 30592
rect 270224 30472 270276 30524
rect 270408 30472 270460 30524
rect 271328 30472 271380 30524
rect 271788 30472 271840 30524
rect 272524 30472 272576 30524
rect 273076 30472 273128 30524
rect 273628 30472 273680 30524
rect 274456 30472 274508 30524
rect 275284 30472 275336 30524
rect 275928 30472 275980 30524
rect 276940 30472 276992 30524
rect 277216 30472 277268 30524
rect 278044 30472 278096 30524
rect 278688 30472 278740 30524
rect 279148 30472 279200 30524
rect 279884 30472 279936 30524
rect 280804 30472 280856 30524
rect 281356 30472 281408 30524
rect 281908 30472 281960 30524
rect 282736 30472 282788 30524
rect 283656 30472 283708 30524
rect 284208 30472 284260 30524
rect 285312 30472 285364 30524
rect 285496 30472 285548 30524
rect 286416 30472 286468 30524
rect 286968 30472 287020 30524
rect 287520 30472 287572 30524
rect 288164 30472 288216 30524
rect 289176 30472 289228 30524
rect 289636 30472 289688 30524
rect 290280 30472 290332 30524
rect 291016 30472 291068 30524
rect 291936 30472 291988 30524
rect 292396 30472 292448 30524
rect 293684 30472 293736 30524
rect 293868 30472 293920 30524
rect 294788 30472 294840 30524
rect 295248 30472 295300 30524
rect 295892 30472 295944 30524
rect 296444 30472 296496 30524
rect 298652 30472 298704 30524
rect 299296 30472 299348 30524
rect 301964 30472 302016 30524
rect 304264 30472 304316 30524
rect 245476 30404 245528 30456
rect 315396 30404 315448 30456
rect 200672 30336 200724 30388
rect 143448 30200 143500 30252
rect 201224 30336 201276 30388
rect 201408 30336 201460 30388
rect 203892 30336 203944 30388
rect 204168 30336 204220 30388
rect 205088 30336 205140 30388
rect 205548 30336 205600 30388
rect 206192 30336 206244 30388
rect 206744 30336 206796 30388
rect 210148 30336 210200 30388
rect 210884 30336 210936 30388
rect 211804 30336 211856 30388
rect 212448 30336 212500 30388
rect 212908 30336 212960 30388
rect 213736 30336 213788 30388
rect 214564 30336 214616 30388
rect 215208 30336 215260 30388
rect 216220 30336 216272 30388
rect 216588 30336 216640 30388
rect 217324 30336 217376 30388
rect 217968 30336 218020 30388
rect 218428 30336 218480 30388
rect 219256 30336 219308 30388
rect 220176 30336 220228 30388
rect 220636 30336 220688 30388
rect 221280 30336 221332 30388
rect 222108 30336 222160 30388
rect 222936 30336 222988 30388
rect 223488 30336 223540 30388
rect 224592 30336 224644 30388
rect 224776 30336 224828 30388
rect 226800 30336 226852 30388
rect 227444 30336 227496 30388
rect 228456 30336 228508 30388
rect 229008 30336 229060 30388
rect 229652 30336 229704 30388
rect 230296 30336 230348 30388
rect 231308 30336 231360 30388
rect 231768 30336 231820 30388
rect 232964 30336 233016 30388
rect 233148 30336 233200 30388
rect 235172 30336 235224 30388
rect 235816 30336 235868 30388
rect 235724 30268 235776 30320
rect 239588 30336 239640 30388
rect 240048 30336 240100 30388
rect 240784 30336 240836 30388
rect 241336 30336 241388 30388
rect 241888 30336 241940 30388
rect 242716 30336 242768 30388
rect 243544 30336 243596 30388
rect 244188 30336 244240 30388
rect 244648 30336 244700 30388
rect 245568 30336 245620 30388
rect 246304 30336 246356 30388
rect 246948 30336 247000 30388
rect 247408 30336 247460 30388
rect 248144 30336 248196 30388
rect 312544 30336 312596 30388
rect 201408 30200 201460 30252
rect 296628 30200 296680 30252
rect 296536 29996 296588 30048
rect 258540 27276 258592 27328
rect 259368 27276 259420 27328
rect 234436 16056 234488 16108
rect 436744 16056 436796 16108
rect 241336 15988 241388 16040
rect 450912 15988 450964 16040
rect 244096 15920 244148 15972
rect 456800 15920 456852 15972
rect 248144 15852 248196 15904
rect 465172 15852 465224 15904
rect 227444 15104 227496 15156
rect 420920 15104 420972 15156
rect 229008 15036 229060 15088
rect 423680 15036 423732 15088
rect 230204 14968 230256 15020
rect 428464 14968 428516 15020
rect 231676 14900 231728 14952
rect 432052 14900 432104 14952
rect 233056 14832 233108 14884
rect 435088 14832 435140 14884
rect 248236 14764 248288 14816
rect 465816 14764 465868 14816
rect 249708 14696 249760 14748
rect 469864 14696 469916 14748
rect 253664 14628 253716 14680
rect 476488 14628 476540 14680
rect 250904 14560 250956 14612
rect 473452 14560 473504 14612
rect 290924 14492 290976 14544
rect 556896 14492 556948 14544
rect 292396 14424 292448 14476
rect 559288 14424 559340 14476
rect 208216 14356 208268 14408
rect 381176 14356 381228 14408
rect 206744 14288 206796 14340
rect 377680 14288 377732 14340
rect 187424 14220 187476 14272
rect 336280 14220 336332 14272
rect 184664 14152 184716 14204
rect 332692 14152 332744 14204
rect 183376 14084 183428 14136
rect 328736 14084 328788 14136
rect 181996 14016 182048 14068
rect 326344 14016 326396 14068
rect 181904 13948 181956 14000
rect 324320 13948 324372 14000
rect 177856 13880 177908 13932
rect 316040 13880 316092 13932
rect 173716 13812 173768 13864
rect 307760 13812 307812 13864
rect 257896 13744 257948 13796
rect 487160 13744 487212 13796
rect 259184 13676 259236 13728
rect 489920 13676 489972 13728
rect 261944 13608 261996 13660
rect 494704 13608 494756 13660
rect 275836 13540 275888 13592
rect 525432 13540 525484 13592
rect 279884 13472 279936 13524
rect 532056 13472 532108 13524
rect 158444 13404 158496 13456
rect 274824 13404 274876 13456
rect 277124 13404 277176 13456
rect 528560 13404 528612 13456
rect 159916 13336 159968 13388
rect 278320 13336 278372 13388
rect 281356 13336 281408 13388
rect 536104 13336 536156 13388
rect 162768 13268 162820 13320
rect 284944 13268 284996 13320
rect 285404 13268 285456 13320
rect 546684 13268 546736 13320
rect 163964 13200 164016 13252
rect 288992 13200 289044 13252
rect 289636 13200 289688 13252
rect 553768 13200 553820 13252
rect 169576 13132 169628 13184
rect 299664 13132 299716 13184
rect 300676 13132 300728 13184
rect 576952 13132 577004 13184
rect 171048 13064 171100 13116
rect 303160 13064 303212 13116
rect 304264 13064 304316 13116
rect 581736 13064 581788 13116
rect 256424 12996 256476 13048
rect 484032 12996 484084 13048
rect 255136 12928 255188 12980
rect 480536 12928 480588 12980
rect 203984 12860 204036 12912
rect 374092 12860 374144 12912
rect 202788 12792 202840 12844
rect 370136 12792 370188 12844
rect 177948 12724 178000 12776
rect 317328 12724 317380 12776
rect 176476 12656 176528 12708
rect 313832 12656 313884 12708
rect 172336 12588 172388 12640
rect 306380 12588 306432 12640
rect 175096 12520 175148 12572
rect 309692 12520 309744 12572
rect 168196 12452 168248 12504
rect 295616 12452 295668 12504
rect 296444 12452 296496 12504
rect 418804 12452 418856 12504
rect 250996 12384 251048 12436
rect 470600 12384 470652 12436
rect 252468 12316 252520 12368
rect 474096 12316 474148 12368
rect 253756 12248 253808 12300
rect 478144 12248 478196 12300
rect 256516 12180 256568 12232
rect 482376 12180 482428 12232
rect 257988 12112 258040 12164
rect 486424 12112 486476 12164
rect 259276 12044 259328 12096
rect 490012 12044 490064 12096
rect 260656 11976 260708 12028
rect 493048 11976 493100 12028
rect 262036 11908 262088 11960
rect 497096 11908 497148 11960
rect 264704 11840 264756 11892
rect 500592 11840 500644 11892
rect 266176 11772 266228 11824
rect 503720 11772 503772 11824
rect 267464 11704 267516 11756
rect 507216 11704 507268 11756
rect 248328 11636 248380 11688
rect 467472 11636 467524 11688
rect 246856 11568 246908 11620
rect 463976 11568 464028 11620
rect 245476 11500 245528 11552
rect 459928 11500 459980 11552
rect 244188 11432 244240 11484
rect 456892 11432 456944 11484
rect 242716 11364 242768 11416
rect 453304 11364 453356 11416
rect 239956 11296 240008 11348
rect 448520 11296 448572 11348
rect 238576 11228 238628 11280
rect 445760 11228 445812 11280
rect 235816 11160 235868 11212
rect 439136 11160 439188 11212
rect 164056 11092 164108 11144
rect 287336 11092 287388 11144
rect 201224 10956 201276 11008
rect 367744 10956 367796 11008
rect 204076 10888 204128 10940
rect 371240 10888 371292 10940
rect 205548 10820 205600 10872
rect 375288 10820 375340 10872
rect 206836 10752 206888 10804
rect 378416 10752 378468 10804
rect 208308 10684 208360 10736
rect 382372 10684 382424 10736
rect 210884 10616 210936 10668
rect 385960 10616 386012 10668
rect 212448 10548 212500 10600
rect 389456 10548 389508 10600
rect 213644 10480 213696 10532
rect 392584 10480 392636 10532
rect 215116 10412 215168 10464
rect 396080 10412 396132 10464
rect 216496 10344 216548 10396
rect 398840 10344 398892 10396
rect 219256 10276 219308 10328
rect 403624 10276 403676 10328
rect 199936 10208 199988 10260
rect 364616 10208 364668 10260
rect 198556 10140 198608 10192
rect 361120 10140 361172 10192
rect 197176 10072 197228 10124
rect 357532 10072 357584 10124
rect 195796 10004 195848 10056
rect 353576 10004 353628 10056
rect 193036 9936 193088 9988
rect 349160 9936 349212 9988
rect 191656 9868 191708 9920
rect 346952 9868 347004 9920
rect 190184 9800 190236 9852
rect 342904 9800 342956 9852
rect 188988 9732 189040 9784
rect 339500 9732 339552 9784
rect 244924 9664 244976 9716
rect 305552 9664 305604 9716
rect 157156 9596 157208 9648
rect 273628 9596 273680 9648
rect 274456 9596 274508 9648
rect 520740 9596 520792 9648
rect 158536 9528 158588 9580
rect 277124 9528 277176 9580
rect 277216 9528 277268 9580
rect 527824 9528 527876 9580
rect 160008 9460 160060 9512
rect 279516 9460 279568 9512
rect 279976 9460 280028 9512
rect 161204 9392 161256 9444
rect 280712 9392 280764 9444
rect 282736 9460 282788 9512
rect 164148 9324 164200 9376
rect 161296 9256 161348 9308
rect 283104 9256 283156 9308
rect 284208 9392 284260 9444
rect 534908 9460 534960 9512
rect 286600 9324 286652 9376
rect 538404 9392 538456 9444
rect 541992 9324 542044 9376
rect 286876 9256 286928 9308
rect 549076 9256 549128 9308
rect 165528 9188 165580 9240
rect 290188 9188 290240 9240
rect 293776 9188 293828 9240
rect 563244 9188 563296 9240
rect 166816 9120 166868 9172
rect 293684 9120 293736 9172
rect 295156 9120 295208 9172
rect 566832 9120 566884 9172
rect 173808 9052 173860 9104
rect 307944 9052 307996 9104
rect 308404 9052 308456 9104
rect 581000 9052 581052 9104
rect 168288 8984 168340 9036
rect 297272 8984 297324 9036
rect 299296 8984 299348 9036
rect 300676 8984 300728 9036
rect 169668 8916 169720 8968
rect 300768 8916 300820 8968
rect 573916 8984 573968 9036
rect 578608 8916 578660 8968
rect 155684 8848 155736 8900
rect 270040 8848 270092 8900
rect 270316 8848 270368 8900
rect 513564 8848 513616 8900
rect 154396 8780 154448 8832
rect 266544 8780 266596 8832
rect 267556 8780 267608 8832
rect 506480 8780 506532 8832
rect 152924 8712 152976 8764
rect 262956 8712 263008 8764
rect 263416 8712 263468 8764
rect 499396 8712 499448 8764
rect 150164 8644 150216 8696
rect 259460 8644 259512 8696
rect 262128 8644 262180 8696
rect 495900 8644 495952 8696
rect 148876 8576 148928 8628
rect 255872 8576 255924 8628
rect 259368 8576 259420 8628
rect 488816 8576 488868 8628
rect 147404 8508 147456 8560
rect 252376 8508 252428 8560
rect 256608 8508 256660 8560
rect 485228 8508 485280 8560
rect 146116 8440 146168 8492
rect 248788 8440 248840 8492
rect 255228 8440 255280 8492
rect 481732 8440 481784 8492
rect 175188 8372 175240 8424
rect 311440 8372 311492 8424
rect 172428 8304 172480 8356
rect 304356 8304 304408 8356
rect 223488 8236 223540 8288
rect 413100 8236 413152 8288
rect 123944 8168 123996 8220
rect 201500 8168 201552 8220
rect 224776 8168 224828 8220
rect 416688 8168 416740 8220
rect 125416 8100 125468 8152
rect 205088 8100 205140 8152
rect 226248 8100 226300 8152
rect 420184 8100 420236 8152
rect 126704 8032 126756 8084
rect 208584 8032 208636 8084
rect 230296 8032 230348 8084
rect 427268 8032 427320 8084
rect 132224 7964 132276 8016
rect 219256 7964 219308 8016
rect 227536 7964 227588 8016
rect 423772 7964 423824 8016
rect 129464 7896 129516 7948
rect 215668 7896 215720 7948
rect 231768 7896 231820 7948
rect 430856 7896 430908 7948
rect 133696 7828 133748 7880
rect 222752 7828 222804 7880
rect 233148 7828 233200 7880
rect 434444 7828 434496 7880
rect 134984 7760 135036 7812
rect 226340 7760 226392 7812
rect 234528 7760 234580 7812
rect 437940 7760 437992 7812
rect 139216 7692 139268 7744
rect 234620 7692 234672 7744
rect 235908 7692 235960 7744
rect 441528 7692 441580 7744
rect 141976 7624 142028 7676
rect 241704 7624 241756 7676
rect 242808 7624 242860 7676
rect 455696 7624 455748 7676
rect 143264 7556 143316 7608
rect 245200 7556 245252 7608
rect 245568 7556 245620 7608
rect 459192 7556 459244 7608
rect 219348 7488 219400 7540
rect 406016 7488 406068 7540
rect 222108 7420 222160 7472
rect 409604 7420 409656 7472
rect 217876 7352 217928 7404
rect 402520 7352 402572 7404
rect 216588 7284 216640 7336
rect 398932 7284 398984 7336
rect 215208 7216 215260 7268
rect 395344 7216 395396 7268
rect 213736 7148 213788 7200
rect 391848 7148 391900 7200
rect 210976 7080 211028 7132
rect 388260 7080 388312 7132
rect 209688 7012 209740 7064
rect 384764 7012 384816 7064
rect 158628 6944 158680 6996
rect 276020 6944 276072 6996
rect 276664 6944 276716 6996
rect 319720 6944 319772 6996
rect 142068 6808 142120 6860
rect 240508 6808 240560 6860
rect 242164 6808 242216 6860
rect 301412 6808 301464 6860
rect 301504 6808 301556 6860
rect 312636 6808 312688 6860
rect 315304 6808 315356 6860
rect 580172 6808 580224 6860
rect 117136 6740 117188 6792
rect 187332 6740 187384 6792
rect 198648 6740 198700 6792
rect 359924 6740 359976 6792
rect 118516 6672 118568 6724
rect 190828 6672 190880 6724
rect 200028 6672 200080 6724
rect 363512 6672 363564 6724
rect 119988 6604 120040 6656
rect 194324 6604 194376 6656
rect 201316 6604 201368 6656
rect 367008 6604 367060 6656
rect 121276 6536 121328 6588
rect 197912 6536 197964 6588
rect 237196 6536 237248 6588
rect 442632 6536 442684 6588
rect 143356 6468 143408 6520
rect 244096 6468 244148 6520
rect 260748 6468 260800 6520
rect 492312 6468 492364 6520
rect 144736 6400 144788 6452
rect 247592 6400 247644 6452
rect 264796 6400 264848 6452
rect 502984 6400 503036 6452
rect 147496 6332 147548 6384
rect 251180 6332 251232 6384
rect 269028 6332 269080 6384
rect 510068 6332 510120 6384
rect 99196 6264 99248 6316
rect 150624 6264 150676 6316
rect 151636 6264 151688 6316
rect 261760 6264 261812 6316
rect 271696 6264 271748 6316
rect 517152 6264 517204 6316
rect 100484 6196 100536 6248
rect 154212 6196 154264 6248
rect 155776 6196 155828 6248
rect 268844 6196 268896 6248
rect 275928 6196 275980 6248
rect 524236 6196 524288 6248
rect 111616 6128 111668 6180
rect 176660 6128 176712 6180
rect 179328 6128 179380 6180
rect 320916 6128 320968 6180
rect 322204 6128 322256 6180
rect 115756 6060 115808 6112
rect 183744 6060 183796 6112
rect 194416 6060 194468 6112
rect 352840 6060 352892 6112
rect 114468 5992 114520 6044
rect 181444 5992 181496 6044
rect 193128 5992 193180 6044
rect 349252 5992 349304 6044
rect 113088 5924 113140 5976
rect 180248 5924 180300 5976
rect 191748 5924 191800 5976
rect 345756 5924 345808 5976
rect 110236 5856 110288 5908
rect 173164 5856 173216 5908
rect 190276 5856 190328 5908
rect 342168 5856 342220 5908
rect 108856 5788 108908 5840
rect 170772 5788 170824 5840
rect 187516 5788 187568 5840
rect 338672 5788 338724 5840
rect 106096 5720 106148 5772
rect 166080 5720 166132 5772
rect 186228 5720 186280 5772
rect 335084 5720 335136 5772
rect 108948 5652 109000 5704
rect 169576 5652 169628 5704
rect 184756 5652 184808 5704
rect 331588 5652 331640 5704
rect 104808 5584 104860 5636
rect 162492 5584 162544 5636
rect 183468 5584 183520 5636
rect 328000 5584 328052 5636
rect 103244 5516 103296 5568
rect 157800 5516 157852 5568
rect 182088 5516 182140 5568
rect 324412 5516 324464 5568
rect 93768 5448 93820 5500
rect 137652 5448 137704 5500
rect 137836 5448 137888 5500
rect 232228 5448 232280 5500
rect 278688 5448 278740 5500
rect 530124 5448 530176 5500
rect 94964 5380 95016 5432
rect 140044 5380 140096 5432
rect 140596 5380 140648 5432
rect 239312 5380 239364 5432
rect 280068 5380 280120 5432
rect 533712 5380 533764 5432
rect 95056 5312 95108 5364
rect 141240 5312 141292 5364
rect 143448 5312 143500 5364
rect 242900 5312 242952 5364
rect 281448 5312 281500 5364
rect 537208 5312 537260 5364
rect 96528 5244 96580 5296
rect 143540 5244 143592 5296
rect 144828 5244 144880 5296
rect 246396 5244 246448 5296
rect 282828 5244 282880 5296
rect 540796 5244 540848 5296
rect 96436 5176 96488 5228
rect 144736 5176 144788 5228
rect 146208 5176 146260 5228
rect 249984 5176 250036 5228
rect 284300 5176 284352 5228
rect 285588 5176 285640 5228
rect 544384 5176 544436 5228
rect 97816 5108 97868 5160
rect 147128 5108 147180 5160
rect 147588 5108 147640 5160
rect 253480 5108 253532 5160
rect 273168 5108 273220 5160
rect 286968 5108 287020 5160
rect 547880 5108 547932 5160
rect 97724 5040 97776 5092
rect 148324 5040 148376 5092
rect 150348 5040 150400 5092
rect 257068 5040 257120 5092
rect 271788 5040 271840 5092
rect 288348 5040 288400 5092
rect 551468 5040 551520 5092
rect 100576 4972 100628 5024
rect 151820 4972 151872 5024
rect 153108 4972 153160 5024
rect 264152 4972 264204 5024
rect 270408 4972 270460 5024
rect 274548 4972 274600 5024
rect 282276 4972 282328 5024
rect 298468 4972 298520 5024
rect 299388 4972 299440 5024
rect 562048 4972 562100 5024
rect 102048 4904 102100 4956
rect 155408 4904 155460 4956
rect 155868 4904 155920 4956
rect 271236 4904 271288 4956
rect 277308 4904 277360 4956
rect 282092 4904 282144 4956
rect 294880 4904 294932 4956
rect 295248 4904 295300 4956
rect 565636 4904 565688 4956
rect 103336 4836 103388 4888
rect 158904 4836 158956 4888
rect 161388 4836 161440 4888
rect 281908 4836 281960 4888
rect 291384 4836 291436 4888
rect 296628 4836 296680 4888
rect 569132 4836 569184 4888
rect 106188 4768 106240 4820
rect 163688 4768 163740 4820
rect 166908 4768 166960 4820
rect 92296 4700 92348 4752
rect 134156 4700 134208 4752
rect 136548 4700 136600 4752
rect 228732 4700 228784 4752
rect 281816 4700 281868 4752
rect 292580 4768 292632 4820
rect 293868 4768 293920 4820
rect 576308 4768 576360 4820
rect 282368 4700 282420 4752
rect 523040 4700 523092 4752
rect 89628 4632 89680 4684
rect 129372 4632 129424 4684
rect 135076 4632 135128 4684
rect 225144 4632 225196 4684
rect 263508 4632 263560 4684
rect 88248 4564 88300 4616
rect 125876 4564 125928 4616
rect 132316 4564 132368 4616
rect 221556 4564 221608 4616
rect 264888 4564 264940 4616
rect 526628 4632 526680 4684
rect 519544 4564 519596 4616
rect 130936 4496 130988 4548
rect 218060 4496 218112 4548
rect 515956 4496 516008 4548
rect 124036 4428 124088 4480
rect 203892 4428 203944 4480
rect 204904 4428 204956 4480
rect 512460 4428 512512 4480
rect 126796 4360 126848 4412
rect 207388 4360 207440 4412
rect 209044 4360 209096 4412
rect 129556 4292 129608 4344
rect 214472 4292 214524 4344
rect 267648 4292 267700 4344
rect 508872 4360 508924 4412
rect 122656 4224 122708 4276
rect 200304 4224 200356 4276
rect 200764 4224 200816 4276
rect 55036 4088 55088 4140
rect 56048 4088 56100 4140
rect 64696 4088 64748 4140
rect 76196 4088 76248 4140
rect 77116 4088 77168 4140
rect 104532 4088 104584 4140
rect 112812 4088 112864 4140
rect 117228 4156 117280 4208
rect 128268 4156 128320 4208
rect 210976 4156 211028 4208
rect 213184 4156 213236 4208
rect 266268 4156 266320 4208
rect 505376 4292 505428 4344
rect 501788 4224 501840 4276
rect 498200 4156 498252 4208
rect 119896 4088 119948 4140
rect 55128 4020 55180 4072
rect 57244 4020 57296 4072
rect 63316 4020 63368 4072
rect 75000 4020 75052 4072
rect 79876 4020 79928 4072
rect 108120 4020 108172 4072
rect 64788 3952 64840 4004
rect 77392 3952 77444 4004
rect 79968 3952 80020 4004
rect 109316 3952 109368 4004
rect 110328 4020 110380 4072
rect 114008 4020 114060 4072
rect 115848 4020 115900 4072
rect 184940 4088 184992 4140
rect 185584 4088 185636 4140
rect 201408 4088 201460 4140
rect 365812 4088 365864 4140
rect 366364 4088 366416 4140
rect 121368 4020 121420 4072
rect 33324 3884 33376 3936
rect 59176 3884 59228 3936
rect 65524 3884 65576 3936
rect 66076 3884 66128 3936
rect 79692 3884 79744 3936
rect 81256 3884 81308 3936
rect 111616 3884 111668 3936
rect 122748 3952 122800 4004
rect 188528 4020 188580 4072
rect 204168 4020 204220 4072
rect 372896 4020 372948 4072
rect 383476 4088 383528 4140
rect 433248 4088 433300 4140
rect 376484 4020 376536 4072
rect 376576 4020 376628 4072
rect 195612 3952 195664 4004
rect 206192 3952 206244 4004
rect 206928 3952 206980 4004
rect 379980 3952 380032 4004
rect 380164 4020 380216 4072
rect 447416 4020 447468 4072
rect 382924 3952 382976 4004
rect 475752 3952 475804 4004
rect 123484 3884 123536 3936
rect 124128 3884 124180 3936
rect 127440 3884 127492 3936
rect 17040 3816 17092 3868
rect 19432 3748 19484 3800
rect 20536 3748 20588 3800
rect 27804 3816 27856 3868
rect 67548 3816 67600 3868
rect 36084 3748 36136 3800
rect 60464 3748 60516 3800
rect 70216 3748 70268 3800
rect 80888 3816 80940 3868
rect 81348 3816 81400 3868
rect 12256 3680 12308 3732
rect 7656 3612 7708 3664
rect 30564 3680 30616 3732
rect 61936 3680 61988 3732
rect 70308 3680 70360 3732
rect 82084 3748 82136 3800
rect 82728 3748 82780 3800
rect 108396 3816 108448 3868
rect 118608 3816 118660 3868
rect 192024 3884 192076 3936
rect 194508 3884 194560 3936
rect 211068 3884 211120 3936
rect 387156 3884 387208 3936
rect 105728 3748 105780 3800
rect 105820 3748 105872 3800
rect 124680 3748 124732 3800
rect 125508 3748 125560 3800
rect 199108 3816 199160 3868
rect 127808 3748 127860 3800
rect 202696 3816 202748 3868
rect 213828 3816 213880 3868
rect 394240 3816 394292 3868
rect 89168 3680 89220 3732
rect 2872 3544 2924 3596
rect 29092 3612 29144 3664
rect 57704 3612 57756 3664
rect 63224 3612 63276 3664
rect 68928 3612 68980 3664
rect 84476 3612 84528 3664
rect 86868 3612 86920 3664
rect 87604 3612 87656 3664
rect 93124 3680 93176 3732
rect 128176 3680 128228 3732
rect 35992 3544 36044 3596
rect 37096 3544 37148 3596
rect 44272 3544 44324 3596
rect 45376 3544 45428 3596
rect 60556 3544 60608 3596
rect 1676 3476 1728 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 27712 3476 27764 3528
rect 28816 3476 28868 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 52460 3476 52512 3528
rect 53748 3476 53800 3528
rect 54024 3476 54076 3528
rect 54944 3476 54996 3528
rect 57888 3476 57940 3528
rect 60832 3476 60884 3528
rect 62028 3544 62080 3596
rect 71504 3544 71556 3596
rect 71688 3544 71740 3596
rect 92756 3544 92808 3596
rect 122288 3612 122340 3664
rect 126888 3612 126940 3664
rect 129648 3612 129700 3664
rect 209780 3748 209832 3800
rect 217968 3748 218020 3800
rect 401324 3816 401376 3868
rect 398840 3748 398892 3800
rect 400128 3748 400180 3800
rect 220728 3680 220780 3732
rect 408408 3680 408460 3732
rect 93952 3544 94004 3596
rect 94504 3544 94556 3596
rect 131764 3544 131816 3596
rect 212172 3612 212224 3664
rect 224868 3612 224920 3664
rect 415492 3612 415544 3664
rect 418804 3612 418856 3664
rect 568028 3612 568080 3664
rect 213368 3544 213420 3596
rect 227628 3544 227680 3596
rect 422576 3544 422628 3596
rect 67916 3476 67968 3528
rect 68836 3476 68888 3528
rect 85672 3476 85724 3528
rect 86776 3476 86828 3528
rect 88984 3476 89036 3528
rect 90364 3476 90416 3528
rect 119344 3476 119396 3528
rect 121092 3476 121144 3528
rect 132408 3476 132460 3528
rect 220452 3476 220504 3528
rect 230388 3476 230440 3528
rect 429660 3544 429712 3596
rect 489920 3544 489972 3596
rect 491116 3544 491168 3596
rect 423680 3476 423732 3528
rect 424968 3476 425020 3528
rect 448520 3476 448572 3528
rect 449808 3476 449860 3528
rect 456800 3476 456852 3528
rect 458088 3476 458140 3528
rect 572 3408 624 3460
rect 27620 3408 27672 3460
rect 57796 3408 57848 3460
rect 62028 3408 62080 3460
rect 69112 3408 69164 3460
rect 71596 3408 71648 3460
rect 91560 3408 91612 3460
rect 92388 3408 92440 3460
rect 135260 3408 135312 3460
rect 137928 3408 137980 3460
rect 231032 3408 231084 3460
rect 237288 3408 237340 3460
rect 443828 3408 443880 3460
rect 8760 3340 8812 3392
rect 9588 3340 9640 3392
rect 9956 3340 10008 3392
rect 10968 3340 11020 3392
rect 11152 3340 11204 3392
rect 12348 3340 12400 3392
rect 15936 3340 15988 3392
rect 16488 3340 16540 3392
rect 18236 3340 18288 3392
rect 19248 3340 19300 3392
rect 24216 3340 24268 3392
rect 24768 3340 24820 3392
rect 25320 3340 25372 3392
rect 26148 3340 26200 3392
rect 59268 3340 59320 3392
rect 64328 3340 64380 3392
rect 66168 3340 66220 3392
rect 63132 3272 63184 3324
rect 73804 3272 73856 3324
rect 63408 3204 63460 3256
rect 72608 3204 72660 3256
rect 56416 3136 56468 3188
rect 59636 3136 59688 3188
rect 60648 3136 60700 3188
rect 66720 3136 66772 3188
rect 65984 3068 66036 3120
rect 78588 3340 78640 3392
rect 78680 3340 78732 3392
rect 104164 3340 104216 3392
rect 106924 3340 106976 3392
rect 107568 3340 107620 3392
rect 108212 3340 108264 3392
rect 115204 3340 115256 3392
rect 70400 3000 70452 3052
rect 87972 3272 88024 3324
rect 90456 3272 90508 3324
rect 116400 3272 116452 3324
rect 75736 3204 75788 3256
rect 101036 3204 101088 3256
rect 101404 3204 101456 3256
rect 77208 3136 77260 3188
rect 102232 3136 102284 3188
rect 108396 3204 108448 3256
rect 112076 3204 112128 3256
rect 177856 3340 177908 3392
rect 174268 3272 174320 3324
rect 175924 3272 175976 3324
rect 167184 3204 167236 3256
rect 177304 3204 177356 3256
rect 193220 3204 193272 3256
rect 74356 3068 74408 3120
rect 98644 3068 98696 3120
rect 75828 3000 75880 3052
rect 99840 3000 99892 3052
rect 56508 2932 56560 2984
rect 58440 2932 58492 2984
rect 74264 2932 74316 2984
rect 97448 2932 97500 2984
rect 97908 2932 97960 2984
rect 103428 3068 103480 3120
rect 160100 3136 160152 3188
rect 160744 3136 160796 3188
rect 100668 3000 100720 3052
rect 153016 3068 153068 3120
rect 155224 3068 155276 3120
rect 161296 3068 161348 3120
rect 170404 3136 170456 3188
rect 189724 3136 189776 3188
rect 190368 3136 190420 3188
rect 197268 3272 197320 3324
rect 355968 3340 356020 3392
rect 349160 3272 349212 3324
rect 350448 3272 350500 3324
rect 351184 3272 351236 3324
rect 344560 3204 344612 3256
rect 351644 3204 351696 3256
rect 351828 3272 351880 3324
rect 358084 3340 358136 3392
rect 369492 3340 369544 3392
rect 373264 3340 373316 3392
rect 426164 3340 426216 3392
rect 355876 3204 355928 3256
rect 383476 3272 383528 3324
rect 383568 3272 383620 3324
rect 418988 3272 419040 3324
rect 337476 3136 337528 3188
rect 337568 3136 337620 3188
rect 344284 3136 344336 3188
rect 369400 3204 369452 3256
rect 411904 3204 411956 3256
rect 404820 3136 404872 3188
rect 175464 3068 175516 3120
rect 177396 3068 177448 3120
rect 181536 3068 181588 3120
rect 237012 3068 237064 3120
rect 307760 3068 307812 3120
rect 309048 3068 309100 3120
rect 309784 3068 309836 3120
rect 461584 3068 461636 3120
rect 583392 3111 583444 3120
rect 583392 3077 583401 3111
rect 583401 3077 583435 3111
rect 583435 3077 583444 3111
rect 583392 3068 583444 3077
rect 149520 3000 149572 3052
rect 156604 3000 156656 3052
rect 164884 3000 164936 3052
rect 167644 3000 167696 3052
rect 182548 3000 182600 3052
rect 184848 3000 184900 3052
rect 73068 2864 73120 2916
rect 95148 2864 95200 2916
rect 95884 2864 95936 2916
rect 96344 2864 96396 2916
rect 74448 2796 74500 2848
rect 96252 2796 96304 2848
rect 95240 2728 95292 2780
rect 96528 2796 96580 2848
rect 99288 2864 99340 2916
rect 145932 2932 145984 2984
rect 166264 2932 166316 2984
rect 179052 2932 179104 2984
rect 180064 2932 180116 2984
rect 142436 2864 142488 2916
rect 142804 2864 142856 2916
rect 156604 2864 156656 2916
rect 157984 2864 158036 2916
rect 168380 2864 168432 2916
rect 169024 2864 169076 2916
rect 186136 2864 186188 2916
rect 187608 3000 187660 3052
rect 330392 3000 330444 3052
rect 330484 3000 330536 3052
rect 333244 3000 333296 3052
rect 348056 3000 348108 3052
rect 362316 3000 362368 3052
rect 362408 3000 362460 3052
rect 397736 3000 397788 3052
rect 233424 2932 233476 2984
rect 315396 2932 315448 2984
rect 454500 2932 454552 2984
rect 196808 2864 196860 2916
rect 323308 2864 323360 2916
rect 323676 2864 323728 2916
rect 333888 2864 333940 2916
rect 138848 2796 138900 2848
rect 159364 2796 159416 2848
rect 171968 2796 172020 2848
rect 173256 2796 173308 2848
rect 229836 2796 229888 2848
rect 312544 2796 312596 2848
rect 324320 2728 324372 2780
rect 325608 2728 325660 2780
rect 340972 2864 341024 2916
rect 341524 2864 341576 2916
rect 355232 2864 355284 2916
rect 355324 2864 355376 2916
rect 358728 2864 358780 2916
rect 390652 2864 390704 2916
rect 440332 2796 440384 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700942 8156 703520
rect 24320 701010 24348 703520
rect 24308 701004 24360 701010
rect 24308 700946 24360 700952
rect 8116 700936 8168 700942
rect 8116 700878 8168 700884
rect 40512 700806 40540 703520
rect 40500 700800 40552 700806
rect 40500 700742 40552 700748
rect 72988 700194 73016 703520
rect 89180 700330 89208 703520
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 98644 700324 98696 700330
rect 98644 700266 98696 700272
rect 72976 700188 73028 700194
rect 72976 700130 73028 700136
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2870 658200 2926 658209
rect 2870 658135 2926 658144
rect 2884 657558 2912 658135
rect 2872 657552 2924 657558
rect 2872 657494 2924 657500
rect 3436 634953 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 32034 645960 32090 645969
rect 4804 645924 4856 645930
rect 32034 645895 32036 645904
rect 4804 645866 4856 645872
rect 32088 645895 32090 645904
rect 32036 645866 32088 645872
rect 3698 639976 3754 639985
rect 3698 639911 3754 639920
rect 3422 634944 3478 634953
rect 3422 634879 3478 634888
rect 3240 633412 3292 633418
rect 3240 633354 3292 633360
rect 3252 632097 3280 633354
rect 3238 632088 3294 632097
rect 3238 632023 3294 632032
rect 3608 621036 3660 621042
rect 3608 620978 3660 620984
rect 3516 619676 3568 619682
rect 3516 619618 3568 619624
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3436 618594 3464 619103
rect 3424 618588 3476 618594
rect 3424 618530 3476 618536
rect 3422 607200 3478 607209
rect 3422 607135 3478 607144
rect 3436 606121 3464 607135
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 3528 605834 3556 619618
rect 3436 605806 3556 605834
rect 3436 593065 3464 605806
rect 3422 593056 3478 593065
rect 3422 592991 3478 593000
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3332 540932 3384 540938
rect 3332 540874 3384 540880
rect 3344 540841 3372 540874
rect 3330 540832 3386 540841
rect 3330 540767 3386 540776
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3332 515432 3384 515438
rect 3332 515374 3384 515380
rect 3344 514865 3372 515374
rect 3330 514856 3386 514865
rect 3330 514791 3386 514800
rect 2870 501800 2926 501809
rect 2870 501735 2926 501744
rect 2884 501022 2912 501735
rect 2872 501016 2924 501022
rect 2872 500958 2924 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3436 314090 3464 579935
rect 3516 578264 3568 578270
rect 3516 578206 3568 578212
rect 3528 436665 3556 578206
rect 3620 488753 3648 620978
rect 3712 566953 3740 639911
rect 3698 566944 3754 566953
rect 3698 566879 3754 566888
rect 3606 488744 3662 488753
rect 3606 488679 3662 488688
rect 3514 436656 3570 436665
rect 3514 436591 3570 436600
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3528 371278 3556 371311
rect 3516 371272 3568 371278
rect 3516 371214 3568 371220
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 3424 314084 3476 314090
rect 3424 314026 3476 314032
rect 3620 312798 3648 358391
rect 3974 345400 4030 345409
rect 3974 345335 4030 345344
rect 3988 312866 4016 345335
rect 3976 312860 4028 312866
rect 3976 312802 4028 312808
rect 3608 312792 3660 312798
rect 3608 312734 3660 312740
rect 3332 312520 3384 312526
rect 3332 312462 3384 312468
rect 2964 306264 3016 306270
rect 2962 306232 2964 306241
rect 3016 306232 3018 306241
rect 2962 306167 3018 306176
rect 2780 293276 2832 293282
rect 2780 293218 2832 293224
rect 2792 293185 2820 293218
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2780 267232 2832 267238
rect 2778 267200 2780 267209
rect 2832 267200 2834 267209
rect 2778 267135 2834 267144
rect 3148 255196 3200 255202
rect 3148 255138 3200 255144
rect 3160 254153 3188 255138
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 2780 241120 2832 241126
rect 2778 241088 2780 241097
rect 2832 241088 2834 241097
rect 2778 241023 2834 241032
rect 2780 215008 2832 215014
rect 2778 214976 2780 214985
rect 2832 214976 2834 214985
rect 2778 214911 2834 214920
rect 3344 201929 3372 312462
rect 3884 312452 3936 312458
rect 3884 312394 3936 312400
rect 3792 312180 3844 312186
rect 3792 312122 3844 312128
rect 3700 311976 3752 311982
rect 3514 311944 3570 311953
rect 3700 311918 3752 311924
rect 3514 311879 3570 311888
rect 3424 309664 3476 309670
rect 3424 309606 3476 309612
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3148 150272 3200 150278
rect 3148 150214 3200 150220
rect 3160 149841 3188 150214
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 2780 123888 2832 123894
rect 2780 123830 2832 123836
rect 2792 123729 2820 123830
rect 2778 123720 2834 123729
rect 2778 123655 2834 123664
rect 2780 111512 2832 111518
rect 2780 111454 2832 111460
rect 2792 110673 2820 111454
rect 2778 110664 2834 110673
rect 2778 110599 2834 110608
rect 2780 85196 2832 85202
rect 2780 85138 2832 85144
rect 2792 84697 2820 85138
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 2780 71664 2832 71670
rect 2778 71632 2780 71641
rect 2832 71632 2834 71641
rect 2778 71567 2834 71576
rect 2780 45552 2832 45558
rect 2778 45520 2780 45529
rect 2832 45520 2834 45529
rect 2778 45455 2834 45464
rect 3436 6497 3464 309606
rect 3528 19417 3556 311879
rect 3608 309732 3660 309738
rect 3608 309674 3660 309680
rect 3620 32473 3648 309674
rect 3712 58585 3740 311918
rect 3804 97617 3832 312122
rect 3896 136785 3924 312394
rect 4712 310140 4764 310146
rect 4712 310082 4764 310088
rect 4068 309868 4120 309874
rect 4068 309810 4120 309816
rect 3976 309800 4028 309806
rect 3976 309742 4028 309748
rect 3988 162897 4016 309742
rect 4080 188873 4108 309810
rect 4724 293282 4752 310082
rect 4712 293276 4764 293282
rect 4712 293218 4764 293224
rect 4066 188864 4122 188873
rect 4066 188799 4122 188808
rect 3974 162888 4030 162897
rect 3974 162823 4030 162832
rect 3882 136776 3938 136785
rect 3882 136711 3938 136720
rect 4816 123894 4844 645866
rect 90822 639976 90878 639985
rect 90822 639911 90824 639920
rect 90876 639911 90878 639920
rect 96342 639976 96398 639985
rect 96342 639911 96344 639920
rect 90824 639882 90876 639888
rect 96396 639911 96398 639920
rect 96344 639882 96396 639888
rect 90824 634976 90876 634982
rect 90822 634944 90824 634953
rect 96988 634976 97040 634982
rect 90876 634944 90878 634953
rect 90822 634879 90878 634888
rect 96986 634944 96988 634953
rect 97040 634944 97042 634953
rect 96986 634879 97042 634888
rect 97908 633412 97960 633418
rect 97908 633354 97960 633360
rect 97920 633321 97948 633354
rect 97906 633312 97962 633321
rect 97906 633247 97962 633256
rect 31758 622160 31814 622169
rect 31758 622095 31814 622104
rect 31772 621042 31800 622095
rect 31760 621036 31812 621042
rect 31760 620978 31812 620984
rect 31758 619712 31814 619721
rect 31758 619647 31760 619656
rect 31812 619647 31814 619656
rect 31760 619618 31812 619624
rect 79244 618594 79824 618610
rect 79232 618588 79836 618594
rect 79284 618582 79784 618588
rect 79232 618530 79284 618536
rect 79784 618530 79836 618536
rect 98656 611354 98684 700266
rect 105464 699990 105492 703520
rect 137848 702434 137876 703520
rect 154132 702434 154160 703520
rect 137848 702406 137968 702434
rect 154132 702406 154436 702434
rect 137100 700324 137152 700330
rect 137100 700266 137152 700272
rect 105452 699984 105504 699990
rect 105452 699926 105504 699932
rect 133604 696992 133656 696998
rect 133604 696934 133656 696940
rect 132788 643346 133184 643362
rect 124772 643340 124824 643346
rect 124772 643282 124824 643288
rect 128912 643340 128964 643346
rect 129280 643340 129332 643346
rect 128964 643300 129280 643328
rect 128912 643282 128964 643288
rect 129280 643282 129332 643288
rect 132776 643340 133196 643346
rect 132828 643334 133144 643340
rect 132776 643282 132828 643288
rect 133144 643282 133196 643288
rect 120262 634944 120318 634953
rect 120262 634879 120264 634888
rect 120316 634879 120318 634888
rect 120264 634850 120316 634856
rect 99746 633312 99802 633321
rect 99746 633247 99802 633256
rect 99760 632738 99788 633247
rect 99748 632732 99800 632738
rect 99748 632674 99800 632680
rect 124128 618044 124180 618050
rect 124128 617986 124180 617992
rect 98472 611326 98684 611354
rect 31758 602304 31814 602313
rect 31758 602239 31814 602248
rect 31772 540938 31800 602239
rect 98472 602041 98500 611326
rect 98458 602032 98514 602041
rect 124140 602002 124168 617986
rect 124784 602002 124812 643282
rect 126794 634944 126850 634953
rect 126794 634879 126796 634888
rect 126848 634879 126850 634888
rect 126796 634850 126848 634856
rect 126888 632732 126940 632738
rect 126888 632674 126940 632680
rect 126900 632369 126928 632674
rect 126886 632360 126942 632369
rect 126886 632295 126942 632304
rect 128268 631440 128320 631446
rect 128268 631382 128320 631388
rect 128912 631440 128964 631446
rect 129280 631440 129332 631446
rect 128964 631400 129280 631428
rect 128912 631382 128964 631388
rect 129280 631382 129332 631388
rect 132776 631440 132828 631446
rect 133144 631440 133196 631446
rect 132828 631388 133144 631394
rect 132776 631382 133196 631388
rect 128280 621926 128308 631382
rect 132788 631366 133184 631382
rect 128268 621920 128320 621926
rect 128268 621862 128320 621868
rect 128268 621376 128320 621382
rect 128268 621318 128320 621324
rect 128280 602002 128308 621318
rect 131488 618044 131540 618050
rect 131488 617986 131540 617992
rect 131500 617114 131528 617986
rect 131500 617098 132080 617114
rect 131500 617092 132092 617098
rect 131500 617086 132040 617092
rect 132040 617034 132092 617040
rect 133616 602002 133644 696934
rect 136652 643346 137048 643362
rect 136640 643340 137060 643346
rect 136692 643334 137008 643340
rect 136640 643282 136692 643288
rect 137008 643282 137060 643288
rect 136640 631440 136692 631446
rect 137008 631440 137060 631446
rect 136692 631388 137008 631394
rect 136640 631382 137060 631388
rect 136652 631366 137048 631382
rect 137112 618934 137140 700266
rect 137100 618928 137152 618934
rect 137100 618870 137152 618876
rect 137100 618316 137152 618322
rect 137100 618258 137152 618264
rect 98458 601967 98514 601976
rect 124128 601996 124180 602002
rect 124128 601938 124180 601944
rect 124772 601996 124824 602002
rect 124772 601938 124824 601944
rect 128268 601996 128320 602002
rect 128268 601938 128320 601944
rect 133604 601996 133656 602002
rect 133604 601938 133656 601944
rect 98642 601624 98698 601633
rect 98642 601559 98698 601568
rect 124128 601588 124180 601594
rect 31850 578368 31906 578377
rect 31850 578303 31906 578312
rect 31864 578270 31892 578303
rect 31852 578264 31904 578270
rect 31852 578206 31904 578212
rect 98656 577998 98684 601559
rect 124128 601530 124180 601536
rect 124772 601588 124824 601594
rect 124772 601530 124824 601536
rect 128268 601588 128320 601594
rect 128268 601530 128320 601536
rect 133604 601588 133656 601594
rect 133604 601530 133656 601536
rect 118606 590744 118662 590753
rect 118606 590679 118662 590688
rect 98644 577992 98696 577998
rect 98644 577934 98696 577940
rect 98644 577584 98696 577590
rect 98644 577526 98696 577532
rect 92388 558952 92440 558958
rect 92388 558894 92440 558900
rect 31760 540932 31812 540938
rect 31760 540874 31812 540880
rect 89628 378208 89680 378214
rect 89628 378150 89680 378156
rect 88248 351960 88300 351966
rect 88248 351902 88300 351908
rect 82544 324352 82596 324358
rect 82544 324294 82596 324300
rect 77668 312996 77720 313002
rect 77668 312938 77720 312944
rect 75276 312928 75328 312934
rect 75276 312870 75328 312876
rect 6368 312724 6420 312730
rect 6368 312666 6420 312672
rect 5356 312656 5408 312662
rect 5356 312598 5408 312604
rect 5172 312316 5224 312322
rect 5172 312258 5224 312264
rect 5080 312248 5132 312254
rect 5080 312190 5132 312196
rect 4988 312112 5040 312118
rect 4988 312054 5040 312060
rect 4896 312044 4948 312050
rect 4896 311986 4948 311992
rect 4804 123888 4856 123894
rect 4804 123830 4856 123836
rect 3790 97608 3846 97617
rect 3790 97543 3846 97552
rect 3698 58576 3754 58585
rect 3698 58511 3754 58520
rect 4908 45558 4936 311986
rect 5000 71670 5028 312054
rect 5092 85202 5120 312190
rect 5184 111518 5212 312258
rect 5264 310004 5316 310010
rect 5264 309946 5316 309952
rect 5276 215014 5304 309946
rect 5368 241126 5396 312598
rect 6276 312588 6328 312594
rect 6276 312530 6328 312536
rect 6184 312384 6236 312390
rect 6184 312326 6236 312332
rect 5448 310072 5500 310078
rect 5448 310014 5500 310020
rect 5460 267238 5488 310014
rect 5448 267232 5500 267238
rect 5448 267174 5500 267180
rect 5356 241120 5408 241126
rect 5356 241062 5408 241068
rect 5264 215008 5316 215014
rect 5264 214950 5316 214956
rect 6196 150278 6224 312326
rect 6288 255202 6316 312530
rect 6380 306270 6408 312666
rect 68006 312352 68062 312361
rect 68006 312287 68062 312296
rect 50986 312216 51042 312225
rect 50986 312151 51042 312160
rect 43994 312080 44050 312089
rect 43994 312015 44050 312024
rect 44008 310706 44036 312015
rect 51000 310706 51028 312151
rect 68020 310706 68048 312287
rect 75288 310706 75316 312870
rect 77680 310706 77708 312938
rect 82556 310706 82584 324294
rect 88260 313070 88288 351902
rect 87328 313064 87380 313070
rect 87328 313006 87380 313012
rect 88248 313064 88300 313070
rect 88248 313006 88300 313012
rect 84936 311908 84988 311914
rect 84936 311850 84988 311856
rect 84948 310706 84976 311850
rect 87340 310706 87368 313006
rect 89640 310706 89668 378150
rect 92400 316034 92428 558894
rect 96528 430636 96580 430642
rect 96528 430578 96580 430584
rect 95148 404388 95200 404394
rect 95148 404330 95200 404336
rect 92216 316006 92428 316034
rect 92216 310706 92244 316006
rect 95160 313070 95188 404330
rect 94504 313064 94556 313070
rect 94504 313006 94556 313012
rect 95148 313064 95200 313070
rect 95148 313006 95200 313012
rect 94516 310706 94544 313006
rect 43700 310678 44036 310706
rect 50876 310678 51028 310706
rect 67712 310678 68048 310706
rect 74980 310678 75316 310706
rect 77372 310678 77708 310706
rect 82156 310678 82584 310706
rect 84640 310678 84976 310706
rect 87032 310678 87368 310706
rect 89424 310678 89668 310706
rect 91816 310678 92244 310706
rect 94208 310678 94544 310706
rect 96540 310706 96568 430578
rect 98656 314226 98684 577526
rect 99288 542428 99340 542434
rect 99288 542370 99340 542376
rect 98644 314220 98696 314226
rect 98644 314162 98696 314168
rect 99300 310706 99328 542370
rect 111708 536852 111760 536858
rect 111708 536794 111760 536800
rect 108948 510672 109000 510678
rect 108948 510614 109000 510620
rect 104808 484424 104860 484430
rect 104808 484366 104860 484372
rect 100760 457496 100812 457502
rect 100760 457438 100812 457444
rect 100772 325694 100800 457438
rect 100772 325666 101076 325694
rect 96540 310678 96600 310706
rect 99084 310678 99328 310706
rect 101048 310706 101076 325666
rect 104820 313070 104848 484366
rect 106188 470620 106240 470626
rect 106188 470562 106240 470568
rect 104164 313064 104216 313070
rect 104164 313006 104216 313012
rect 104808 313064 104860 313070
rect 104808 313006 104860 313012
rect 104176 310706 104204 313006
rect 101048 310678 101476 310706
rect 103868 310678 104204 310706
rect 106200 310706 106228 470562
rect 108960 310706 108988 510614
rect 111720 316034 111748 536794
rect 115848 533384 115900 533390
rect 115848 533326 115900 533332
rect 114468 524476 114520 524482
rect 114468 524418 114520 524424
rect 111444 316006 111748 316034
rect 111444 310706 111472 316006
rect 114480 313070 114508 524418
rect 113824 313064 113876 313070
rect 113824 313006 113876 313012
rect 114468 313064 114520 313070
rect 114468 313006 114520 313012
rect 113836 310706 113864 313006
rect 106200 310678 106260 310706
rect 108652 310678 108988 310706
rect 111044 310678 111472 310706
rect 113528 310678 113864 310706
rect 115860 310706 115888 533326
rect 118620 310706 118648 590679
rect 121366 576872 121422 576881
rect 121366 576807 121422 576816
rect 121380 316034 121408 576807
rect 121104 316006 121408 316034
rect 121104 310706 121132 316006
rect 124140 313070 124168 601530
rect 124784 313070 124812 601530
rect 123392 313064 123444 313070
rect 123392 313006 123444 313012
rect 124128 313064 124180 313070
rect 124128 313006 124180 313012
rect 124772 313064 124824 313070
rect 124772 313006 124824 313012
rect 125232 313064 125284 313070
rect 125232 313006 125284 313012
rect 123404 310706 123432 313006
rect 115860 310678 115920 310706
rect 118312 310678 118648 310706
rect 120704 310678 121132 310706
rect 123096 310678 123432 310706
rect 125244 310706 125272 313006
rect 128280 310706 128308 601530
rect 130660 313948 130712 313954
rect 130660 313890 130712 313896
rect 130672 310706 130700 313890
rect 133616 313070 133644 601530
rect 135076 314016 135128 314022
rect 135076 313958 135128 313964
rect 133052 313064 133104 313070
rect 133052 313006 133104 313012
rect 133604 313064 133656 313070
rect 133604 313006 133656 313012
rect 133064 310706 133092 313006
rect 125244 310678 125580 310706
rect 127972 310678 128308 310706
rect 130364 310678 130700 310706
rect 132756 310678 133092 310706
rect 135088 310570 135116 313958
rect 137112 310706 137140 618258
rect 137940 313070 137968 702406
rect 148324 700596 148376 700602
rect 148324 700538 148376 700544
rect 144828 700460 144880 700466
rect 144828 700402 144880 700408
rect 140688 700392 140740 700398
rect 140688 700334 140740 700340
rect 139492 577516 139544 577522
rect 139492 577458 139544 577464
rect 139504 576881 139532 577458
rect 139490 576872 139546 576881
rect 139490 576807 139546 576816
rect 140700 316034 140728 700334
rect 143448 533452 143500 533458
rect 143448 533394 143500 533400
rect 140424 316006 140728 316034
rect 137928 313064 137980 313070
rect 137928 313006 137980 313012
rect 140424 310706 140452 316006
rect 143460 313138 143488 533394
rect 142712 313132 142764 313138
rect 142712 313074 142764 313080
rect 143448 313132 143500 313138
rect 143448 313074 143500 313080
rect 142724 310706 142752 313074
rect 144840 310978 144868 700402
rect 148336 313138 148364 700538
rect 150348 700528 150400 700534
rect 150348 700470 150400 700476
rect 150360 313138 150388 700470
rect 153106 639840 153162 639849
rect 153106 639775 153162 639784
rect 153120 313138 153148 639775
rect 154408 313206 154436 702406
rect 164148 700868 164200 700874
rect 164148 700810 164200 700816
rect 154488 700732 154540 700738
rect 154488 700674 154540 700680
rect 154396 313200 154448 313206
rect 154396 313142 154448 313148
rect 147496 313132 147548 313138
rect 147496 313074 147548 313080
rect 148324 313132 148376 313138
rect 148324 313074 148376 313080
rect 149888 313132 149940 313138
rect 149888 313074 149940 313080
rect 150348 313132 150400 313138
rect 150348 313074 150400 313080
rect 152280 313132 152332 313138
rect 152280 313074 152332 313080
rect 153108 313132 153160 313138
rect 153108 313074 153160 313080
rect 137112 310678 137540 310706
rect 140024 310678 140452 310706
rect 142416 310678 142752 310706
rect 144794 310950 144868 310978
rect 144794 310692 144822 310950
rect 147508 310706 147536 313074
rect 149900 310706 149928 313074
rect 152292 310706 152320 313074
rect 154500 310978 154528 700674
rect 157248 700664 157300 700670
rect 157248 700606 157300 700612
rect 147200 310678 147536 310706
rect 149592 310678 149928 310706
rect 151984 310678 152320 310706
rect 154454 310950 154528 310978
rect 154454 310692 154482 310950
rect 157260 310706 157288 700606
rect 162768 700256 162820 700262
rect 162768 700198 162820 700204
rect 160006 640112 160062 640121
rect 160006 640047 160062 640056
rect 159548 591320 159600 591326
rect 159548 591262 159600 591268
rect 159560 590753 159588 591262
rect 159546 590744 159602 590753
rect 159546 590679 159602 590688
rect 160020 313138 160048 640047
rect 160098 607200 160154 607209
rect 160098 607135 160100 607144
rect 160152 607135 160154 607144
rect 160926 607200 160982 607209
rect 160926 607135 160928 607144
rect 160100 607106 160152 607112
rect 160980 607135 160982 607144
rect 160928 607106 160980 607112
rect 162780 313206 162808 700198
rect 161940 313200 161992 313206
rect 161940 313142 161992 313148
rect 162768 313200 162820 313206
rect 162768 313142 162820 313148
rect 159548 313132 159600 313138
rect 159548 313074 159600 313080
rect 160008 313132 160060 313138
rect 160008 313074 160060 313080
rect 159560 310706 159588 313074
rect 161952 310706 161980 313142
rect 164160 310706 164188 700810
rect 169668 700052 169720 700058
rect 169668 699994 169720 700000
rect 166816 314152 166868 314158
rect 166816 314094 166868 314100
rect 166828 310706 166856 314094
rect 169680 313206 169708 699994
rect 170324 699718 170352 703520
rect 196348 701004 196400 701010
rect 196348 700946 196400 700952
rect 188988 700936 189040 700942
rect 188988 700878 189040 700884
rect 188344 700188 188396 700194
rect 188344 700130 188396 700136
rect 188436 700188 188488 700194
rect 188436 700130 188488 700136
rect 172428 700120 172480 700126
rect 172428 700062 172480 700068
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 171060 314294 171088 699654
rect 171048 314288 171100 314294
rect 171048 314230 171100 314236
rect 172440 313206 172468 700062
rect 187976 699984 188028 699990
rect 187976 699926 188028 699932
rect 173808 699916 173860 699922
rect 173808 699858 173860 699864
rect 169208 313200 169260 313206
rect 169208 313142 169260 313148
rect 169668 313200 169720 313206
rect 169668 313142 169720 313148
rect 171600 313200 171652 313206
rect 171600 313142 171652 313148
rect 172428 313200 172480 313206
rect 172428 313142 172480 313148
rect 169220 310706 169248 313142
rect 171612 310706 171640 313142
rect 173820 310706 173848 699858
rect 175924 699848 175976 699854
rect 175924 699790 175976 699796
rect 156860 310678 157288 310706
rect 159252 310678 159588 310706
rect 161644 310678 161980 310706
rect 164036 310678 164188 310706
rect 166520 310678 166856 310706
rect 168912 310678 169248 310706
rect 171304 310678 171640 310706
rect 173696 310678 173848 310706
rect 175936 310706 175964 699790
rect 187988 654134 188016 699926
rect 187988 654106 188108 654134
rect 188080 645658 188108 654106
rect 188356 645658 188384 700130
rect 188448 645658 188476 700130
rect 188528 670744 188580 670750
rect 188528 670686 188580 670692
rect 188540 645930 188568 670686
rect 188528 645924 188580 645930
rect 188528 645866 188580 645872
rect 188068 645652 188120 645658
rect 188068 645594 188120 645600
rect 188344 645652 188396 645658
rect 188344 645594 188396 645600
rect 188436 645652 188488 645658
rect 188436 645594 188488 645600
rect 187976 645380 188028 645386
rect 187976 645322 188028 645328
rect 188436 645380 188488 645386
rect 188436 645322 188488 645328
rect 182914 639296 182970 639305
rect 182914 639231 182970 639240
rect 182928 639130 182956 639231
rect 184018 639160 184074 639169
rect 182916 639124 182968 639130
rect 184018 639095 184074 639104
rect 182916 639066 182968 639072
rect 184032 639062 184060 639095
rect 184020 639056 184072 639062
rect 182546 639024 182602 639033
rect 184020 638998 184072 639004
rect 182546 638959 182548 638968
rect 182600 638959 182602 638968
rect 182548 638930 182600 638936
rect 187988 638858 188016 645322
rect 188448 638858 188476 645322
rect 189000 638858 189028 700878
rect 196360 645590 196388 700946
rect 202800 699854 202828 703520
rect 218992 700194 219020 703520
rect 227720 700800 227772 700806
rect 227720 700742 227772 700748
rect 218980 700188 219032 700194
rect 218980 700130 219032 700136
rect 202788 699848 202840 699854
rect 202788 699790 202840 699796
rect 197820 657552 197872 657558
rect 197820 657494 197872 657500
rect 197832 652754 197860 657494
rect 197832 652726 198228 652754
rect 198200 645930 198228 652726
rect 227732 647154 227760 700742
rect 235184 699922 235212 703520
rect 235172 699916 235224 699922
rect 235172 699858 235224 699864
rect 251468 699718 251496 703520
rect 267660 700058 267688 703520
rect 283852 700126 283880 703520
rect 283840 700120 283892 700126
rect 283840 700062 283892 700068
rect 267648 700052 267700 700058
rect 267648 699994 267700 700000
rect 251456 699712 251508 699718
rect 251456 699654 251508 699660
rect 252468 699712 252520 699718
rect 252468 699654 252520 699660
rect 252480 669361 252508 699654
rect 252466 669352 252522 669361
rect 252466 669287 252522 669296
rect 227720 647148 227772 647154
rect 227720 647090 227772 647096
rect 226156 646400 226208 646406
rect 226156 646342 226208 646348
rect 226168 646066 226196 646342
rect 226156 646060 226208 646066
rect 226156 646002 226208 646008
rect 198188 645924 198240 645930
rect 198188 645866 198240 645872
rect 196348 645584 196400 645590
rect 196348 645526 196400 645532
rect 197912 645176 197964 645182
rect 197912 645118 197964 645124
rect 196900 642388 196952 642394
rect 196900 642330 196952 642336
rect 196912 640914 196940 642330
rect 196912 640886 197124 640914
rect 196992 640756 197044 640762
rect 196992 640698 197044 640704
rect 194692 639532 194744 639538
rect 194692 639474 194744 639480
rect 194600 639464 194652 639470
rect 194600 639406 194652 639412
rect 194612 639169 194640 639406
rect 194704 639305 194732 639474
rect 194690 639296 194746 639305
rect 194690 639231 194746 639240
rect 194598 639160 194654 639169
rect 194598 639095 194654 639104
rect 196348 639124 196400 639130
rect 196348 639066 196400 639072
rect 187976 638852 188028 638858
rect 187976 638794 188028 638800
rect 188436 638852 188488 638858
rect 188436 638794 188488 638800
rect 188988 638852 189040 638858
rect 188988 638794 189040 638800
rect 188988 638580 189040 638586
rect 188988 638522 189040 638528
rect 187976 638512 188028 638518
rect 187976 638454 188028 638460
rect 188344 638512 188396 638518
rect 188344 638454 188396 638460
rect 188436 638512 188488 638518
rect 188436 638454 188488 638460
rect 176198 635216 176254 635225
rect 176254 635174 176424 635202
rect 176198 635151 176254 635160
rect 176396 634930 176424 635174
rect 176566 634944 176622 634953
rect 176396 634902 176566 634930
rect 176566 634879 176622 634888
rect 184202 634944 184258 634953
rect 184754 634944 184810 634953
rect 184258 634902 184754 634930
rect 184202 634879 184258 634888
rect 184754 634879 184810 634888
rect 184202 632496 184258 632505
rect 184754 632496 184810 632505
rect 184258 632454 184754 632482
rect 184202 632431 184258 632440
rect 184754 632431 184810 632440
rect 187988 624714 188016 638454
rect 188356 624714 188384 638454
rect 188448 624714 188476 638454
rect 188528 638376 188580 638382
rect 188528 638318 188580 638324
rect 188540 624714 188568 638318
rect 189000 624714 189028 638522
rect 196256 638444 196308 638450
rect 196256 638386 196308 638392
rect 196268 635662 196296 638386
rect 196360 635662 196388 639066
rect 197004 638450 197032 640698
rect 197096 639130 197124 640886
rect 197452 639600 197504 639606
rect 197452 639542 197504 639548
rect 197084 639124 197136 639130
rect 197084 639066 197136 639072
rect 197464 639033 197492 639542
rect 197450 639024 197506 639033
rect 197450 638959 197506 638968
rect 196992 638444 197044 638450
rect 196992 638386 197044 638392
rect 197924 636194 197952 645118
rect 199568 641028 199620 641034
rect 199568 640970 199620 640976
rect 214564 641028 214616 641034
rect 214564 640970 214616 640976
rect 197832 636166 197952 636194
rect 197832 636018 197860 636166
rect 197832 635990 198504 636018
rect 196256 635656 196308 635662
rect 196256 635598 196308 635604
rect 196348 635656 196400 635662
rect 196348 635598 196400 635604
rect 196164 635384 196216 635390
rect 196164 635326 196216 635332
rect 189262 634944 189318 634953
rect 189262 634879 189264 634888
rect 189316 634879 189318 634888
rect 191562 634944 191618 634953
rect 191562 634879 191564 634888
rect 189264 634850 189316 634856
rect 191616 634879 191618 634888
rect 191564 634850 191616 634856
rect 196176 634001 196204 635326
rect 196348 635180 196400 635186
rect 196348 635122 196400 635128
rect 196360 634001 196388 635122
rect 198476 634030 198504 635990
rect 199580 634030 199608 640970
rect 205362 639024 205418 639033
rect 205362 638959 205418 638968
rect 205376 636820 205404 638959
rect 214576 637906 214604 640970
rect 233884 639600 233936 639606
rect 233884 639542 233936 639548
rect 233896 639305 233924 639542
rect 233882 639296 233938 639305
rect 233882 639231 233938 639240
rect 218886 639024 218942 639033
rect 218886 638959 218942 638968
rect 218900 637906 218928 638959
rect 214564 637900 214616 637906
rect 214564 637842 214616 637848
rect 218888 637900 218940 637906
rect 218888 637842 218940 637848
rect 214564 637628 214616 637634
rect 214564 637570 214616 637576
rect 218888 637628 218940 637634
rect 218888 637570 218940 637576
rect 201866 634944 201922 634953
rect 201866 634879 201922 634888
rect 201880 634250 201908 634879
rect 201880 634236 202233 634250
rect 201880 634222 202247 634236
rect 198464 634024 198516 634030
rect 196162 633992 196218 634001
rect 196162 633927 196218 633936
rect 196346 633992 196402 634001
rect 198464 633966 198516 633972
rect 199568 634024 199620 634030
rect 199568 633966 199620 633972
rect 196346 633927 196402 633936
rect 202219 633758 202247 634222
rect 202207 633752 202259 633758
rect 196346 633720 196402 633729
rect 202207 633694 202259 633700
rect 196346 633655 196402 633664
rect 196254 633584 196310 633593
rect 196254 633519 196310 633528
rect 189814 632496 189870 632505
rect 189814 632431 189816 632440
rect 189868 632431 189870 632440
rect 191564 632460 191616 632466
rect 189816 632402 189868 632408
rect 191564 632402 191616 632408
rect 191576 632369 191604 632402
rect 191562 632360 191618 632369
rect 191562 632295 191618 632304
rect 191564 631440 191616 631446
rect 191562 631408 191564 631417
rect 191616 631408 191618 631417
rect 191562 631343 191618 631352
rect 192942 631408 192998 631417
rect 192942 631343 192998 631352
rect 192956 631174 192984 631343
rect 192944 631168 192996 631174
rect 192944 631110 192996 631116
rect 187976 624708 188028 624714
rect 187976 624650 188028 624656
rect 188344 624708 188396 624714
rect 188344 624650 188396 624656
rect 188436 624708 188488 624714
rect 188436 624650 188488 624656
rect 188528 624708 188580 624714
rect 188528 624650 188580 624656
rect 188988 624708 189040 624714
rect 188988 624650 189040 624656
rect 187976 624368 188028 624374
rect 187976 624310 188028 624316
rect 188344 624368 188396 624374
rect 188344 624310 188396 624316
rect 188436 624368 188488 624374
rect 188436 624310 188488 624316
rect 188528 624368 188580 624374
rect 188528 624310 188580 624316
rect 188988 624368 189040 624374
rect 188988 624310 189040 624316
rect 180892 314288 180944 314294
rect 180892 314230 180944 314236
rect 178776 313200 178828 313206
rect 178776 313142 178828 313148
rect 178788 310706 178816 313142
rect 175936 310678 176088 310706
rect 178480 310678 178816 310706
rect 180904 310706 180932 314230
rect 185400 313132 185452 313138
rect 185400 313074 185452 313080
rect 183008 313064 183060 313070
rect 183008 313006 183060 313012
rect 183020 310706 183048 313006
rect 185412 310706 185440 313074
rect 187988 310706 188016 624310
rect 188356 313274 188384 624310
rect 188344 313268 188396 313274
rect 188344 313210 188396 313216
rect 188448 313206 188476 624310
rect 188436 313200 188488 313206
rect 188436 313142 188488 313148
rect 188540 313138 188568 624310
rect 188528 313132 188580 313138
rect 188528 313074 188580 313080
rect 189000 313070 189028 624310
rect 192576 314220 192628 314226
rect 192576 314162 192628 314168
rect 190460 313268 190512 313274
rect 190460 313210 190512 313216
rect 188988 313064 189040 313070
rect 188988 313006 189040 313012
rect 190472 310706 190500 313210
rect 192588 310706 192616 314162
rect 196268 313070 196296 633519
rect 196360 313274 196388 633655
rect 214576 632806 214604 637570
rect 218900 636002 218928 637570
rect 218888 635996 218940 636002
rect 218888 635938 218940 635944
rect 214564 632800 214616 632806
rect 214564 632742 214616 632748
rect 198464 632528 198516 632534
rect 198464 632470 198516 632476
rect 199568 632528 199620 632534
rect 199568 632470 199620 632476
rect 198476 628318 198504 632470
rect 199580 628318 199608 632470
rect 201960 632256 202012 632262
rect 201960 632198 202012 632204
rect 210238 632224 210294 632233
rect 198464 628312 198516 628318
rect 198464 628254 198516 628260
rect 199568 628312 199620 628318
rect 199568 628254 199620 628260
rect 201972 628250 202000 632198
rect 210238 632159 210294 632168
rect 210252 628250 210280 632159
rect 215392 631780 215444 631786
rect 215392 631722 215444 631728
rect 215404 631281 215432 631722
rect 215390 631272 215446 631281
rect 215390 631207 215446 631216
rect 221094 631272 221150 631281
rect 221094 631207 221150 631216
rect 221108 630698 221136 631207
rect 221096 630692 221148 630698
rect 221096 630634 221148 630640
rect 218888 629128 218940 629134
rect 218888 629070 218940 629076
rect 201960 628244 202012 628250
rect 201960 628186 202012 628192
rect 210240 628244 210292 628250
rect 210240 628186 210292 628192
rect 214564 628244 214616 628250
rect 214564 628186 214616 628192
rect 210976 628040 211028 628046
rect 210976 627982 211028 627988
rect 197360 627972 197412 627978
rect 197360 627914 197412 627920
rect 197820 627972 197872 627978
rect 197820 627914 197872 627920
rect 199568 627972 199620 627978
rect 199568 627914 199620 627920
rect 197372 515438 197400 627914
rect 197360 515432 197412 515438
rect 197360 515374 197412 515380
rect 197372 514826 197400 515374
rect 197360 514820 197412 514826
rect 197360 514762 197412 514768
rect 196348 313268 196400 313274
rect 196348 313210 196400 313216
rect 197832 313206 197860 627914
rect 199580 618594 199608 627914
rect 201960 627904 202012 627910
rect 201960 627846 202012 627852
rect 199568 618588 199620 618594
rect 199568 618530 199620 618536
rect 198004 514820 198056 514826
rect 198004 514762 198056 514768
rect 198016 314226 198044 514762
rect 200764 462392 200816 462398
rect 200764 462334 200816 462340
rect 198004 314220 198056 314226
rect 198004 314162 198056 314168
rect 200120 313268 200172 313274
rect 200120 313210 200172 313216
rect 197452 313200 197504 313206
rect 197452 313142 197504 313148
rect 197820 313200 197872 313206
rect 197820 313142 197872 313148
rect 195704 313064 195756 313070
rect 195704 313006 195756 313012
rect 196256 313064 196308 313070
rect 196256 313006 196308 313012
rect 195716 310706 195744 313006
rect 180904 310678 180964 310706
rect 183020 310678 183356 310706
rect 185412 310678 185748 310706
rect 187988 310678 188140 310706
rect 190472 310678 190532 310706
rect 192588 310678 192924 310706
rect 195408 310678 195744 310706
rect 197464 310706 197492 313142
rect 200132 310706 200160 313210
rect 200776 313070 200804 462334
rect 201972 325694 202000 627846
rect 204902 607200 204958 607209
rect 204902 607135 204958 607144
rect 201972 325666 202184 325694
rect 200764 313064 200816 313070
rect 200764 313006 200816 313012
rect 202156 310706 202184 325666
rect 204916 313274 204944 607135
rect 210988 316034 211016 627982
rect 214576 626822 214604 628186
rect 218900 627774 218928 629070
rect 218888 627768 218940 627774
rect 218888 627710 218940 627716
rect 214564 626816 214616 626822
rect 214564 626758 214616 626764
rect 214564 626612 214616 626618
rect 214564 626554 214616 626560
rect 211804 553444 211856 553450
rect 211804 553386 211856 553392
rect 210252 316006 211016 316034
rect 204904 313268 204956 313274
rect 204904 313210 204956 313216
rect 204628 313200 204680 313206
rect 204628 313142 204680 313148
rect 204640 310706 204668 313142
rect 207020 313132 207072 313138
rect 207020 313074 207072 313080
rect 207032 310706 207060 313074
rect 210252 310706 210280 316006
rect 211816 313138 211844 553386
rect 211896 313268 211948 313274
rect 211896 313210 211948 313216
rect 211804 313132 211856 313138
rect 211804 313074 211856 313080
rect 197464 310678 197800 310706
rect 200132 310678 200192 310706
rect 202156 310678 202584 310706
rect 204640 310678 204976 310706
rect 207032 310678 207368 310706
rect 209852 310678 210280 310706
rect 211908 310706 211936 313210
rect 214576 310706 214604 626554
rect 218888 620016 218940 620022
rect 218888 619958 218940 619964
rect 218704 501016 218756 501022
rect 218704 500958 218756 500964
rect 216680 314084 216732 314090
rect 216680 314026 216732 314032
rect 216692 310706 216720 314026
rect 218716 313206 218744 500958
rect 218900 313274 218928 619958
rect 223580 527196 223632 527202
rect 223580 527138 223632 527144
rect 221464 409896 221516 409902
rect 221464 409838 221516 409844
rect 218888 313268 218940 313274
rect 218888 313210 218940 313216
rect 218704 313200 218756 313206
rect 218704 313142 218756 313148
rect 221476 313138 221504 409838
rect 223592 325694 223620 527138
rect 230480 474768 230532 474774
rect 230480 474710 230532 474716
rect 226984 448588 227036 448594
rect 226984 448530 227036 448536
rect 223592 325666 223896 325694
rect 221556 313268 221608 313274
rect 221556 313210 221608 313216
rect 219072 313132 219124 313138
rect 219072 313074 219124 313080
rect 221464 313132 221516 313138
rect 221464 313074 221516 313080
rect 219084 310706 219112 313074
rect 221568 310706 221596 313210
rect 223868 310706 223896 325666
rect 226996 313206 227024 448530
rect 230492 325694 230520 474710
rect 237380 422340 237432 422346
rect 237380 422282 237432 422288
rect 233884 397520 233936 397526
rect 233884 397462 233936 397468
rect 230492 325666 231072 325694
rect 228732 314220 228784 314226
rect 228732 314162 228784 314168
rect 226340 313200 226392 313206
rect 226340 313142 226392 313148
rect 226984 313200 227036 313206
rect 226984 313142 227036 313148
rect 226352 310706 226380 313142
rect 228744 310706 228772 314162
rect 231044 310706 231072 325666
rect 233896 313274 233924 397462
rect 237392 325694 237420 422282
rect 245660 371272 245712 371278
rect 245660 371214 245712 371220
rect 237392 325666 238340 325694
rect 233884 313268 233936 313274
rect 233884 313210 233936 313216
rect 233516 313200 233568 313206
rect 233516 313142 233568 313148
rect 233528 310706 233556 313142
rect 236000 313064 236052 313070
rect 236000 313006 236052 313012
rect 236012 310706 236040 313006
rect 238312 310706 238340 325666
rect 240784 313268 240836 313274
rect 240784 313210 240836 313216
rect 240796 310706 240824 313210
rect 243176 313132 243228 313138
rect 243176 313074 243228 313080
rect 243188 310706 243216 313074
rect 245672 310706 245700 371214
rect 252744 318844 252796 318850
rect 252744 318786 252796 318792
rect 247960 312860 248012 312866
rect 247960 312802 248012 312808
rect 247972 310706 248000 312802
rect 250444 312792 250496 312798
rect 250444 312734 250496 312740
rect 250456 310706 250484 312734
rect 252756 310706 252784 318786
rect 299492 314158 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700262 332548 703520
rect 348804 700874 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700868 348844 700874
rect 348792 700810 348844 700816
rect 332508 700256 332560 700262
rect 332508 700198 332560 700204
rect 364352 639169 364380 702406
rect 381188 699718 381216 703520
rect 397472 700738 397500 703520
rect 397460 700732 397512 700738
rect 397460 700674 397512 700680
rect 413664 700670 413692 703520
rect 413652 700664 413704 700670
rect 413652 700606 413704 700612
rect 381176 699712 381228 699718
rect 381176 699654 381228 699660
rect 382188 699712 382240 699718
rect 382188 699654 382240 699660
rect 364338 639160 364394 639169
rect 364338 639095 364394 639104
rect 382200 619682 382228 699654
rect 410616 692844 410668 692850
rect 410616 692786 410668 692792
rect 404266 632088 404322 632097
rect 404266 632023 404322 632032
rect 382188 619676 382240 619682
rect 382188 619618 382240 619624
rect 404280 566914 404308 632023
rect 410628 569974 410656 692786
rect 429212 648378 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700602 462360 703520
rect 462320 700596 462372 700602
rect 462320 700538 462372 700544
rect 478524 700534 478552 703520
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 527192 700398 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 463330 692880 463386 692889
rect 463330 692815 463332 692824
rect 463384 692815 463386 692824
rect 465538 692880 465594 692889
rect 465594 692838 465750 692866
rect 465538 692815 465594 692824
rect 463332 692786 463384 692792
rect 542372 670410 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580354 683904 580410 683913
rect 580354 683839 580410 683848
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 542360 670404 542412 670410
rect 542360 670346 542412 670352
rect 542360 668432 542412 668438
rect 542360 668374 542412 668380
rect 429200 648372 429252 648378
rect 429200 648314 429252 648320
rect 429200 648100 429252 648106
rect 429200 648042 429252 648048
rect 429212 640257 429240 648042
rect 471888 644904 471940 644910
rect 471888 644846 471940 644852
rect 471900 644609 471928 644846
rect 459558 644600 459614 644609
rect 459558 644535 459614 644544
rect 468666 644600 468722 644609
rect 469034 644600 469090 644609
rect 468722 644558 469034 644586
rect 468666 644535 468722 644544
rect 469034 644535 469090 644544
rect 471886 644600 471942 644609
rect 471886 644535 471942 644544
rect 459572 644502 459600 644535
rect 459560 644496 459612 644502
rect 459560 644438 459612 644444
rect 443644 643204 443696 643210
rect 443644 643146 443696 643152
rect 415306 640248 415362 640257
rect 415306 640183 415362 640192
rect 423586 640248 423642 640257
rect 424230 640248 424286 640257
rect 423642 640206 424230 640234
rect 423586 640183 423642 640192
rect 424230 640183 424286 640192
rect 429198 640248 429254 640257
rect 429198 640183 429254 640192
rect 415320 639606 415348 640183
rect 415308 639600 415360 639606
rect 415308 639542 415360 639548
rect 436744 631848 436796 631854
rect 436744 631790 436796 631796
rect 436756 631281 436784 631790
rect 414662 631272 414718 631281
rect 414662 631207 414718 631216
rect 422666 631272 422722 631281
rect 423402 631272 423458 631281
rect 422722 631230 423402 631258
rect 422666 631207 422722 631216
rect 423402 631207 423458 631216
rect 436742 631272 436798 631281
rect 436742 631207 436798 631216
rect 414676 628998 414704 631207
rect 414664 628992 414716 628998
rect 414664 628934 414716 628940
rect 410340 569968 410392 569974
rect 410340 569910 410392 569916
rect 410616 569968 410668 569974
rect 410616 569910 410668 569916
rect 410352 567610 410380 569910
rect 410044 567582 410380 567610
rect 404268 566908 404320 566914
rect 404268 566850 404320 566856
rect 427820 566500 427872 566506
rect 427820 566442 427872 566448
rect 391846 559464 391902 559473
rect 391846 559399 391902 559408
rect 391860 558958 391888 559399
rect 391848 558952 391900 558958
rect 391848 558894 391900 558900
rect 391386 543552 391442 543561
rect 391386 543487 391442 543496
rect 391400 542434 391428 543487
rect 391388 542428 391440 542434
rect 391388 542370 391440 542376
rect 391756 542428 391808 542434
rect 391756 542370 391808 542376
rect 391768 419490 391796 542370
rect 391756 419484 391808 419490
rect 391756 419426 391808 419432
rect 391860 365702 391888 558894
rect 427832 551585 427860 566442
rect 427818 551576 427874 551585
rect 427818 551511 427874 551520
rect 402040 535758 402100 535786
rect 402072 534002 402100 535758
rect 417712 535622 418048 535650
rect 417712 534070 417740 535622
rect 417700 534064 417752 534070
rect 417700 534006 417752 534012
rect 401600 533996 401652 534002
rect 401600 533938 401652 533944
rect 402060 533996 402112 534002
rect 402060 533938 402112 533944
rect 401612 533458 401640 533938
rect 401600 533452 401652 533458
rect 401600 533394 401652 533400
rect 417712 533390 417740 534006
rect 417700 533384 417752 533390
rect 417700 533326 417752 533332
rect 391848 365696 391900 365702
rect 391848 365638 391900 365644
rect 299480 314152 299532 314158
rect 299480 314094 299532 314100
rect 443656 314022 443684 643146
rect 506664 631236 506716 631242
rect 506664 631178 506716 631184
rect 506676 631145 506704 631178
rect 496082 631136 496138 631145
rect 496082 631071 496138 631080
rect 506662 631136 506718 631145
rect 506662 631071 506718 631080
rect 496096 630834 496124 631071
rect 496084 630828 496136 630834
rect 496084 630770 496136 630776
rect 542372 623082 542400 668374
rect 579618 644056 579674 644065
rect 579618 643991 579674 644000
rect 579632 643346 579660 643991
rect 579620 643340 579672 643346
rect 579620 643282 579672 643288
rect 579804 631372 579856 631378
rect 579804 631314 579856 631320
rect 579816 630873 579844 631314
rect 579802 630864 579858 630873
rect 579802 630799 579858 630808
rect 542360 623076 542412 623082
rect 542360 623018 542412 623024
rect 542452 619880 542504 619886
rect 542452 619822 542504 619828
rect 542464 611354 542492 619822
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 617098 580212 617471
rect 580172 617092 580224 617098
rect 580172 617034 580224 617040
rect 542372 611326 542492 611354
rect 542372 534002 542400 611326
rect 580172 591320 580224 591326
rect 580172 591262 580224 591268
rect 580184 591025 580212 591262
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 579986 577688 580042 577697
rect 579986 577623 580042 577632
rect 580000 577522 580028 577623
rect 579988 577516 580040 577522
rect 579988 577458 580040 577464
rect 579620 569968 579672 569974
rect 579620 569910 579672 569916
rect 542360 533996 542412 534002
rect 542360 533938 542412 533944
rect 579632 458153 579660 569910
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 579986 484664 580042 484673
rect 579986 484599 580042 484608
rect 580000 484430 580028 484599
rect 579988 484424 580040 484430
rect 579988 484366 580040 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 579618 458144 579674 458153
rect 579618 458079 579674 458088
rect 579632 457502 579660 458079
rect 579620 457496 579672 457502
rect 579620 457438 579672 457444
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 579908 430642 579936 431559
rect 579896 430636 579948 430642
rect 579896 430578 579948 430584
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 443644 314016 443696 314022
rect 443644 313958 443696 313964
rect 580276 313954 580304 670647
rect 580368 645862 580396 683839
rect 580356 645856 580408 645862
rect 580356 645798 580408 645804
rect 580354 564360 580410 564369
rect 580354 564295 580410 564304
rect 580368 534070 580396 564295
rect 580356 534064 580408 534070
rect 580356 534006 580408 534012
rect 580264 313948 580316 313954
rect 580264 313890 580316 313896
rect 303436 312996 303488 313002
rect 303436 312938 303488 312944
rect 257620 312724 257672 312730
rect 257620 312666 257672 312672
rect 257632 310706 257660 312666
rect 262496 312656 262548 312662
rect 262496 312598 262548 312604
rect 262508 310706 262536 312598
rect 264980 312588 265032 312594
rect 264980 312530 265032 312536
rect 264992 310706 265020 312530
rect 272064 312520 272116 312526
rect 272064 312462 272116 312468
rect 272076 310706 272104 312462
rect 276940 312452 276992 312458
rect 276940 312394 276992 312400
rect 276952 310706 276980 312394
rect 279332 312384 279384 312390
rect 279332 312326 279384 312332
rect 279344 310706 279372 312326
rect 281724 312316 281776 312322
rect 281724 312258 281776 312264
rect 281736 310706 281764 312258
rect 284300 312248 284352 312254
rect 284300 312190 284352 312196
rect 303250 312216 303306 312225
rect 284312 310706 284340 312190
rect 286508 312180 286560 312186
rect 303250 312151 303306 312160
rect 286508 312122 286560 312128
rect 286520 310706 286548 312122
rect 288900 312112 288952 312118
rect 288900 312054 288952 312060
rect 303066 312080 303122 312089
rect 288912 310706 288940 312054
rect 291384 312044 291436 312050
rect 303066 312015 303122 312024
rect 291384 311986 291436 311992
rect 291396 310706 291424 311986
rect 293960 311976 294012 311982
rect 293960 311918 294012 311924
rect 300950 311944 301006 311953
rect 293972 310706 294000 311918
rect 300950 311879 301006 311888
rect 300964 310706 300992 311879
rect 211908 310678 212244 310706
rect 214576 310678 214636 310706
rect 216692 310678 217028 310706
rect 219084 310678 219420 310706
rect 221568 310678 221904 310706
rect 223868 310678 224296 310706
rect 226352 310678 226688 310706
rect 228744 310678 229080 310706
rect 231044 310678 231472 310706
rect 233528 310678 233864 310706
rect 236012 310678 236348 310706
rect 238312 310678 238740 310706
rect 240796 310678 241132 310706
rect 243188 310678 243524 310706
rect 245672 310678 245916 310706
rect 247972 310678 248308 310706
rect 250456 310678 250792 310706
rect 252756 310678 253184 310706
rect 257632 310678 257968 310706
rect 262508 310678 262844 310706
rect 264992 310678 265236 310706
rect 272076 310678 272412 310706
rect 276952 310678 277288 310706
rect 279344 310678 279680 310706
rect 281736 310678 282072 310706
rect 284312 310678 284464 310706
rect 286520 310678 286856 310706
rect 288912 310678 289248 310706
rect 291396 310678 291732 310706
rect 293972 310678 294124 310706
rect 300964 310678 301300 310706
rect 31648 310554 31800 310570
rect 31648 310548 31812 310554
rect 31648 310542 31760 310548
rect 135088 310542 135148 310570
rect 302884 310548 302936 310554
rect 31760 310490 31812 310496
rect 302884 310490 302936 310496
rect 79968 310480 80020 310486
rect 65320 310418 65656 310434
rect 72588 310418 72924 310434
rect 79764 310428 79968 310434
rect 79764 310422 80020 310428
rect 65320 310412 65668 310418
rect 65320 310406 65616 310412
rect 72588 310412 72936 310418
rect 72588 310406 72884 310412
rect 65616 310354 65668 310360
rect 79764 310406 80008 310422
rect 72884 310354 72936 310360
rect 60648 310344 60700 310350
rect 55660 310282 55996 310298
rect 58144 310282 58480 310298
rect 60536 310292 60648 310298
rect 63224 310344 63276 310350
rect 60536 310286 60700 310292
rect 62928 310292 63224 310298
rect 70308 310344 70360 310350
rect 62928 310286 63276 310292
rect 70104 310292 70308 310298
rect 70104 310286 70360 310292
rect 55660 310276 56008 310282
rect 55660 310270 55956 310276
rect 58144 310276 58492 310282
rect 58144 310270 58440 310276
rect 55956 310218 56008 310224
rect 60536 310270 60688 310286
rect 62928 310270 63264 310286
rect 70104 310270 70348 310286
rect 58440 310218 58492 310224
rect 39120 310208 39172 310214
rect 29550 310176 29606 310185
rect 29256 310134 29550 310162
rect 38824 310156 39120 310162
rect 41328 310208 41380 310214
rect 38824 310150 39172 310156
rect 41216 310156 41328 310162
rect 46388 310208 46440 310214
rect 41216 310150 41380 310156
rect 46092 310156 46388 310162
rect 48780 310208 48832 310214
rect 46092 310150 46440 310156
rect 48484 310156 48780 310162
rect 53564 310208 53616 310214
rect 48484 310150 48832 310156
rect 53268 310156 53564 310162
rect 53268 310150 53616 310156
rect 38824 310134 39160 310150
rect 41216 310134 41368 310150
rect 46092 310134 46428 310150
rect 48484 310134 48820 310150
rect 53268 310134 53604 310150
rect 255332 310146 255576 310162
rect 255320 310140 255576 310146
rect 29550 310111 29606 310120
rect 255372 310134 255576 310140
rect 255320 310082 255372 310088
rect 260012 310072 260064 310078
rect 34334 310040 34390 310049
rect 34040 309998 34334 310026
rect 36726 310040 36782 310049
rect 36432 309998 36726 310026
rect 34334 309975 34390 309984
rect 260064 310020 260360 310026
rect 260012 310014 260360 310020
rect 260024 309998 260360 310014
rect 267292 310010 267628 310026
rect 269684 310010 270020 310026
rect 274652 310010 274804 310026
rect 296180 310010 296516 310026
rect 298572 310010 298908 310026
rect 267280 310004 267628 310010
rect 36726 309975 36782 309984
rect 267332 309998 267628 310004
rect 269672 310004 270020 310010
rect 267280 309946 267332 309952
rect 269724 309998 270020 310004
rect 274640 310004 274804 310010
rect 269672 309946 269724 309952
rect 274692 309998 274804 310004
rect 296168 310004 296516 310010
rect 274640 309946 274692 309952
rect 296220 309998 296516 310004
rect 298560 310004 298908 310010
rect 296168 309946 296220 309952
rect 298612 309998 298908 310004
rect 298560 309946 298612 309952
rect 6368 306264 6420 306270
rect 6368 306206 6420 306212
rect 6276 255196 6328 255202
rect 6276 255138 6328 255144
rect 6184 150272 6236 150278
rect 6184 150214 6236 150220
rect 5172 111512 5224 111518
rect 5172 111454 5224 111460
rect 5080 85196 5132 85202
rect 5080 85138 5132 85144
rect 4988 71664 5040 71670
rect 4988 71606 5040 71612
rect 4896 45552 4948 45558
rect 4896 45494 4948 45500
rect 27632 34054 28336 34082
rect 28552 34054 28888 34082
rect 29104 34054 29440 34082
rect 29656 34054 29992 34082
rect 30392 34054 30544 34082
rect 30760 34054 31096 34082
rect 31312 34054 31648 34082
rect 31864 34054 32200 34082
rect 32416 34054 32752 34082
rect 33152 34054 33304 34082
rect 33520 34054 33856 34082
rect 34072 34054 34408 34082
rect 34624 34054 34960 34082
rect 35176 34054 35512 34082
rect 3606 32464 3662 32473
rect 3606 32399 3662 32408
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 19248 31680 19300 31686
rect 19248 31622 19300 31628
rect 16488 31612 16540 31618
rect 16488 31554 16540 31560
rect 13728 31544 13780 31550
rect 13728 31486 13780 31492
rect 10968 31408 11020 31414
rect 10968 31350 11020 31356
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 6828 31204 6880 31210
rect 6828 31146 6880 31152
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 2884 480 2912 3538
rect 4080 480 4108 31078
rect 5448 31068 5500 31074
rect 5448 31010 5500 31016
rect 5460 6914 5488 31010
rect 6840 6914 6868 31146
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7668 480 7696 3606
rect 9600 3398 9628 31214
rect 10980 3398 11008 31350
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 8772 480 8800 3334
rect 9968 480 9996 3334
rect 11164 480 11192 3334
rect 12268 1850 12296 3674
rect 12360 3398 12388 31282
rect 13740 6914 13768 31486
rect 15108 31476 15160 31482
rect 15108 31418 15160 31424
rect 15120 6914 15148 31418
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12268 1822 12388 1850
rect 12360 480 12388 1822
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3398 16528 31554
rect 17040 3868 17092 3874
rect 17040 3810 17092 3816
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 15948 480 15976 3334
rect 17052 480 17080 3810
rect 19260 3398 19288 31622
rect 20548 16574 20576 31690
rect 23388 31000 23440 31006
rect 23388 30942 23440 30948
rect 20628 30932 20680 30938
rect 20628 30874 20680 30880
rect 20456 16546 20576 16574
rect 19432 3800 19484 3806
rect 19432 3742 19484 3748
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 18248 480 18276 3334
rect 19444 480 19472 3742
rect 20456 3482 20484 16546
rect 20640 6914 20668 30874
rect 22008 30864 22060 30870
rect 22008 30806 22060 30812
rect 22020 6914 22048 30806
rect 23400 6914 23428 30942
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 20548 6886 20668 6914
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20548 3806 20576 6886
rect 20536 3800 20588 3806
rect 20536 3742 20588 3748
rect 20456 3454 20668 3482
rect 20640 480 20668 3454
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3398 24808 30738
rect 27528 30660 27580 30666
rect 27528 30602 27580 30608
rect 26148 30592 26200 30598
rect 26148 30534 26200 30540
rect 26160 3398 26188 30534
rect 27540 3534 27568 30602
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 24228 480 24256 3334
rect 25332 480 25360 3334
rect 26528 480 26556 3470
rect 27632 3466 27660 34054
rect 28552 26234 28580 34054
rect 28908 30728 28960 30734
rect 28908 30670 28960 30676
rect 28816 30524 28868 30530
rect 28816 30466 28868 30472
rect 27816 26206 28580 26234
rect 27816 3874 27844 26206
rect 27804 3868 27856 3874
rect 27804 3810 27856 3816
rect 28828 3534 28856 30466
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 27620 3460 27672 3466
rect 27620 3402 27672 3408
rect 27724 480 27752 3470
rect 28920 480 28948 30670
rect 29104 3670 29132 34054
rect 29656 31142 29684 34054
rect 29644 31136 29696 31142
rect 29644 31078 29696 31084
rect 30288 31136 30340 31142
rect 30288 31078 30340 31084
rect 30300 6914 30328 31078
rect 30392 31074 30420 34054
rect 30760 31210 30788 34054
rect 30748 31204 30800 31210
rect 30748 31146 30800 31152
rect 30380 31068 30432 31074
rect 30380 31010 30432 31016
rect 31312 26234 31340 34054
rect 31864 31278 31892 34054
rect 32416 31414 32444 34054
rect 32404 31408 32456 31414
rect 32404 31350 32456 31356
rect 33152 31346 33180 34054
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 31852 31272 31904 31278
rect 31852 31214 31904 31220
rect 33048 31204 33100 31210
rect 33048 31146 33100 31152
rect 31668 31068 31720 31074
rect 31668 31010 31720 31016
rect 30116 6886 30328 6914
rect 30576 26206 31340 26234
rect 29092 3664 29144 3670
rect 29092 3606 29144 3612
rect 30116 480 30144 6886
rect 30576 3738 30604 26206
rect 31680 6914 31708 31010
rect 31312 6886 31708 6914
rect 30564 3732 30616 3738
rect 30564 3674 30616 3680
rect 31312 480 31340 6886
rect 33060 3534 33088 31146
rect 33520 26234 33548 34054
rect 34072 31550 34100 34054
rect 34060 31544 34112 31550
rect 34060 31486 34112 31492
rect 34624 31482 34652 34054
rect 35176 31618 35204 34054
rect 36050 33810 36078 34068
rect 36280 34054 36616 34082
rect 36832 34054 37168 34082
rect 37384 34054 37720 34082
rect 37936 34054 38272 34082
rect 38672 34054 38916 34082
rect 39132 34054 39468 34082
rect 39684 34054 40020 34082
rect 40236 34054 40572 34082
rect 40788 34054 41124 34082
rect 41432 34054 41676 34082
rect 41892 34054 42228 34082
rect 42444 34054 42780 34082
rect 42996 34054 43332 34082
rect 43548 34054 43884 34082
rect 44192 34054 44436 34082
rect 44652 34054 44988 34082
rect 45204 34054 45540 34082
rect 45756 34054 46092 34082
rect 46308 34054 46644 34082
rect 46952 34054 47196 34082
rect 47412 34054 47748 34082
rect 47964 34054 48300 34082
rect 48516 34054 48852 34082
rect 49160 34054 49496 34082
rect 49712 34054 50048 34082
rect 50264 34054 50600 34082
rect 51092 34054 51152 34082
rect 51276 34054 51704 34082
rect 51828 34054 52256 34082
rect 52564 34054 52808 34082
rect 53024 34054 53360 34082
rect 53912 34054 54064 34082
rect 54464 34054 54892 34082
rect 55016 34054 55168 34082
rect 55568 34054 55904 34082
rect 56120 34054 56456 34082
rect 56672 34054 57008 34082
rect 57224 34054 57560 34082
rect 36050 33782 36124 33810
rect 35164 31612 35216 31618
rect 35164 31554 35216 31560
rect 34612 31476 34664 31482
rect 34612 31418 34664 31424
rect 34428 31340 34480 31346
rect 34428 31282 34480 31288
rect 33336 26206 33548 26234
rect 33336 3942 33364 26206
rect 33324 3936 33376 3942
rect 33324 3878 33376 3884
rect 34440 3534 34468 31282
rect 35808 31272 35860 31278
rect 35808 31214 35860 31220
rect 35820 3534 35848 31214
rect 36096 3806 36124 33782
rect 36280 31686 36308 34054
rect 36268 31680 36320 31686
rect 36268 31622 36320 31628
rect 36832 30938 36860 34054
rect 37384 31754 37412 34054
rect 37372 31748 37424 31754
rect 37372 31690 37424 31696
rect 36820 30932 36872 30938
rect 36820 30874 36872 30880
rect 37936 30870 37964 34054
rect 38568 31476 38620 31482
rect 38568 31418 38620 31424
rect 37924 30864 37976 30870
rect 37924 30806 37976 30812
rect 37096 30456 37148 30462
rect 37096 30398 37148 30404
rect 37108 16574 37136 30398
rect 37188 30388 37240 30394
rect 37188 30330 37240 30336
rect 37016 16546 37136 16574
rect 36084 3800 36136 3806
rect 36084 3742 36136 3748
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34808 480 34836 3470
rect 36004 480 36032 3538
rect 37016 3482 37044 16546
rect 37200 6914 37228 30330
rect 38580 6914 38608 31418
rect 38672 31006 38700 34054
rect 38660 31000 38712 31006
rect 38660 30942 38712 30948
rect 39132 30802 39160 34054
rect 39120 30796 39172 30802
rect 39120 30738 39172 30744
rect 39684 30598 39712 34054
rect 39948 31000 40000 31006
rect 39948 30942 40000 30948
rect 39672 30592 39724 30598
rect 39672 30534 39724 30540
rect 39960 6914 39988 30942
rect 40236 30666 40264 34054
rect 40224 30660 40276 30666
rect 40224 30602 40276 30608
rect 40788 30530 40816 34054
rect 41328 31748 41380 31754
rect 41328 31690 41380 31696
rect 40776 30524 40828 30530
rect 40776 30466 40828 30472
rect 37108 6886 37228 6914
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 37108 3602 37136 6886
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 37016 3454 37228 3482
rect 37200 480 37228 3454
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3534 41368 31690
rect 41432 30734 41460 34054
rect 41892 31142 41920 34054
rect 41880 31136 41932 31142
rect 41880 31078 41932 31084
rect 42444 31074 42472 34054
rect 42708 31612 42760 31618
rect 42708 31554 42760 31560
rect 42432 31068 42484 31074
rect 42432 31010 42484 31016
rect 41420 30728 41472 30734
rect 41420 30670 41472 30676
rect 42720 3534 42748 31554
rect 42996 31210 43024 34054
rect 43548 31346 43576 34054
rect 44088 31680 44140 31686
rect 44088 31622 44140 31628
rect 43536 31340 43588 31346
rect 43536 31282 43588 31288
rect 42984 31204 43036 31210
rect 42984 31146 43036 31152
rect 44100 3534 44128 31622
rect 44192 31278 44220 34054
rect 44180 31272 44232 31278
rect 44180 31214 44232 31220
rect 44652 30394 44680 34054
rect 45204 30462 45232 34054
rect 45756 31482 45784 34054
rect 45744 31476 45796 31482
rect 45744 31418 45796 31424
rect 45468 31272 45520 31278
rect 45468 31214 45520 31220
rect 45376 31136 45428 31142
rect 45376 31078 45428 31084
rect 45192 30456 45244 30462
rect 45192 30398 45244 30404
rect 44640 30388 44692 30394
rect 44640 30330 44692 30336
rect 45388 16574 45416 31078
rect 45296 16546 45416 16574
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3538
rect 45296 3482 45324 16546
rect 45480 6914 45508 31214
rect 46308 31006 46336 34054
rect 46952 31754 46980 34054
rect 46940 31748 46992 31754
rect 46940 31690 46992 31696
rect 47412 31618 47440 34054
rect 47964 31686 47992 34054
rect 47952 31680 48004 31686
rect 47952 31622 48004 31628
rect 47400 31612 47452 31618
rect 47400 31554 47452 31560
rect 48516 31278 48544 34054
rect 48504 31272 48556 31278
rect 48504 31214 48556 31220
rect 49160 31142 49188 34054
rect 49148 31136 49200 31142
rect 49148 31078 49200 31084
rect 46296 31000 46348 31006
rect 46296 30942 46348 30948
rect 49608 30524 49660 30530
rect 49608 30466 49660 30472
rect 46848 30456 46900 30462
rect 46848 30398 46900 30404
rect 46860 6914 46888 30398
rect 48228 30388 48280 30394
rect 48228 30330 48280 30336
rect 48240 6914 48268 30330
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 45388 3602 45416 6886
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45296 3454 45508 3482
rect 45480 480 45508 3454
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3534 49648 30466
rect 49712 30462 49740 34054
rect 49700 30456 49752 30462
rect 49700 30398 49752 30404
rect 50264 30394 50292 34054
rect 51092 30530 51120 34054
rect 51080 30524 51132 30530
rect 51080 30466 51132 30472
rect 51276 30410 51304 34054
rect 50252 30388 50304 30394
rect 50252 30330 50304 30336
rect 51000 30382 51304 30410
rect 51000 3534 51028 30382
rect 51828 26234 51856 34054
rect 52460 30388 52512 30394
rect 52460 30330 52512 30336
rect 51276 26206 51856 26234
rect 51276 16574 51304 26206
rect 51276 16546 51396 16574
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51368 480 51396 16546
rect 52472 3534 52500 30330
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 34054
rect 53024 30394 53052 34054
rect 53012 30388 53064 30394
rect 53012 30330 53064 30336
rect 54036 3534 54064 34054
rect 54864 26234 54892 34054
rect 54864 26206 55076 26234
rect 55048 4146 55076 26206
rect 55036 4140 55088 4146
rect 55036 4082 55088 4088
rect 55140 4078 55168 34054
rect 55876 30394 55904 34054
rect 55864 30388 55916 30394
rect 55864 30330 55916 30336
rect 56048 4140 56100 4146
rect 56048 4082 56100 4088
rect 55128 4072 55180 4078
rect 55128 4014 55180 4020
rect 53748 3528 53800 3534
rect 53748 3470 53800 3476
rect 54024 3528 54076 3534
rect 54024 3470 54076 3476
rect 54944 3528 54996 3534
rect 54944 3470 54996 3476
rect 53760 480 53788 3470
rect 54956 480 54984 3470
rect 56060 480 56088 4082
rect 56428 3194 56456 34054
rect 56980 30462 57008 34054
rect 56968 30456 57020 30462
rect 56968 30398 57020 30404
rect 57532 30394 57560 34054
rect 57716 34054 57776 34082
rect 58328 34054 58664 34082
rect 58880 34054 59216 34082
rect 59432 34054 59768 34082
rect 60076 34054 60412 34082
rect 56508 30388 56560 30394
rect 56508 30330 56560 30336
rect 57520 30388 57572 30394
rect 57520 30330 57572 30336
rect 56416 3188 56468 3194
rect 56416 3130 56468 3136
rect 56520 2990 56548 30330
rect 57244 4072 57296 4078
rect 57244 4014 57296 4020
rect 56508 2984 56560 2990
rect 56508 2926 56560 2932
rect 57256 480 57284 4014
rect 57716 3670 57744 34054
rect 57888 30456 57940 30462
rect 57888 30398 57940 30404
rect 57796 30388 57848 30394
rect 57796 30330 57848 30336
rect 57704 3664 57756 3670
rect 57704 3606 57756 3612
rect 57808 3466 57836 30330
rect 57900 3534 57928 30398
rect 58636 30394 58664 34054
rect 58624 30388 58676 30394
rect 58624 30330 58676 30336
rect 59188 3942 59216 34054
rect 59740 30462 59768 34054
rect 59728 30456 59780 30462
rect 59728 30398 59780 30404
rect 60384 30394 60412 34054
rect 60476 34054 60628 34082
rect 61180 34054 61516 34082
rect 61732 34054 62068 34082
rect 62284 34054 62620 34082
rect 62836 34054 63264 34082
rect 59268 30388 59320 30394
rect 59268 30330 59320 30336
rect 60372 30388 60424 30394
rect 60372 30330 60424 30336
rect 59176 3936 59228 3942
rect 59176 3878 59228 3884
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 57796 3460 57848 3466
rect 57796 3402 57848 3408
rect 59280 3398 59308 30330
rect 60476 3806 60504 34054
rect 60648 30456 60700 30462
rect 60648 30398 60700 30404
rect 60556 30388 60608 30394
rect 60556 30330 60608 30336
rect 60464 3800 60516 3806
rect 60464 3742 60516 3748
rect 60568 3602 60596 30330
rect 60556 3596 60608 3602
rect 60556 3538 60608 3544
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 60660 3194 60688 30398
rect 61488 30394 61516 34054
rect 61476 30388 61528 30394
rect 61476 30330 61528 30336
rect 61936 30388 61988 30394
rect 61936 30330 61988 30336
rect 61948 3738 61976 30330
rect 61936 3732 61988 3738
rect 61936 3674 61988 3680
rect 62040 3602 62068 34054
rect 62592 30394 62620 34054
rect 62580 30388 62632 30394
rect 62580 30330 62632 30336
rect 63236 6914 63264 34054
rect 63144 6886 63264 6914
rect 63328 34054 63388 34082
rect 63940 34054 64276 34082
rect 64492 34054 64828 34082
rect 65044 34054 65380 34082
rect 65596 34054 66024 34082
rect 62028 3596 62080 3602
rect 62028 3538 62080 3544
rect 60832 3528 60884 3534
rect 60832 3470 60884 3476
rect 59636 3188 59688 3194
rect 59636 3130 59688 3136
rect 60648 3188 60700 3194
rect 60648 3130 60700 3136
rect 58440 2984 58492 2990
rect 58440 2926 58492 2932
rect 58452 480 58480 2926
rect 59648 480 59676 3130
rect 60844 480 60872 3470
rect 62028 3460 62080 3466
rect 62028 3402 62080 3408
rect 62040 480 62068 3402
rect 63144 3330 63172 6886
rect 63328 4078 63356 34054
rect 64248 30394 64276 34054
rect 63408 30388 63460 30394
rect 63408 30330 63460 30336
rect 64236 30388 64288 30394
rect 64236 30330 64288 30336
rect 64696 30388 64748 30394
rect 64696 30330 64748 30336
rect 63316 4072 63368 4078
rect 63316 4014 63368 4020
rect 63224 3664 63276 3670
rect 63224 3606 63276 3612
rect 63132 3324 63184 3330
rect 63132 3266 63184 3272
rect 63236 480 63264 3606
rect 63420 3262 63448 30330
rect 64708 4146 64736 30330
rect 64696 4140 64748 4146
rect 64696 4082 64748 4088
rect 64800 4010 64828 34054
rect 65352 30394 65380 34054
rect 65340 30388 65392 30394
rect 65340 30330 65392 30336
rect 65892 30388 65944 30394
rect 65892 30330 65944 30336
rect 65904 26234 65932 30330
rect 65996 30138 66024 34054
rect 66134 33810 66162 34068
rect 66700 34054 67036 34082
rect 67252 34054 67588 34082
rect 67804 34054 68140 34082
rect 68356 34054 68784 34082
rect 66134 33782 66208 33810
rect 65996 30110 66116 30138
rect 65904 26206 66024 26234
rect 64788 4004 64840 4010
rect 64788 3946 64840 3952
rect 65524 3936 65576 3942
rect 65524 3878 65576 3884
rect 64328 3392 64380 3398
rect 64328 3334 64380 3340
rect 63408 3256 63460 3262
rect 63408 3198 63460 3204
rect 64340 480 64368 3334
rect 65536 480 65564 3878
rect 65996 3126 66024 26206
rect 66088 3942 66116 30110
rect 66076 3936 66128 3942
rect 66076 3878 66128 3884
rect 66180 3398 66208 33782
rect 67008 30394 67036 34054
rect 67560 31074 67588 34054
rect 67548 31068 67600 31074
rect 67548 31010 67600 31016
rect 68112 30394 68140 34054
rect 66996 30388 67048 30394
rect 66996 30330 67048 30336
rect 67548 30388 67600 30394
rect 67548 30330 67600 30336
rect 68100 30388 68152 30394
rect 68100 30330 68152 30336
rect 67560 3874 67588 30330
rect 68756 26234 68784 34054
rect 68848 34054 68908 34082
rect 69460 34054 69796 34082
rect 70012 34054 70256 34082
rect 70656 34054 70992 34082
rect 71208 34054 71636 34082
rect 68848 31686 68876 34054
rect 68836 31680 68888 31686
rect 68836 31622 68888 31628
rect 69768 30394 69796 34054
rect 68928 30388 68980 30394
rect 68928 30330 68980 30336
rect 69756 30388 69808 30394
rect 69756 30330 69808 30336
rect 68756 26206 68876 26234
rect 67548 3868 67600 3874
rect 67548 3810 67600 3816
rect 68848 3534 68876 26206
rect 68940 3670 68968 30330
rect 70228 3806 70256 34054
rect 70964 31414 70992 34054
rect 70952 31408 71004 31414
rect 70952 31350 71004 31356
rect 70308 30388 70360 30394
rect 70308 30330 70360 30336
rect 70320 3890 70348 30330
rect 70320 3862 70440 3890
rect 70216 3800 70268 3806
rect 70216 3742 70268 3748
rect 70308 3732 70360 3738
rect 70308 3674 70360 3680
rect 68928 3664 68980 3670
rect 68928 3606 68980 3612
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68836 3528 68888 3534
rect 68836 3470 68888 3476
rect 66168 3392 66220 3398
rect 66168 3334 66220 3340
rect 66720 3188 66772 3194
rect 66720 3130 66772 3136
rect 65984 3120 66036 3126
rect 65984 3062 66036 3068
rect 66732 480 66760 3130
rect 67928 480 67956 3470
rect 69112 3460 69164 3466
rect 69112 3402 69164 3408
rect 69124 480 69152 3402
rect 70320 480 70348 3674
rect 70412 3058 70440 3862
rect 71504 3596 71556 3602
rect 71504 3538 71556 3544
rect 70400 3052 70452 3058
rect 70400 2994 70452 3000
rect 71516 480 71544 3538
rect 71608 3466 71636 34054
rect 71700 34054 71760 34082
rect 72312 34054 72648 34082
rect 72864 34054 73108 34082
rect 73416 34054 73752 34082
rect 73968 34054 74304 34082
rect 71700 3602 71728 34054
rect 72620 31550 72648 34054
rect 72608 31544 72660 31550
rect 72608 31486 72660 31492
rect 71688 3596 71740 3602
rect 71688 3538 71740 3544
rect 71596 3460 71648 3466
rect 71596 3402 71648 3408
rect 72608 3256 72660 3262
rect 72608 3198 72660 3204
rect 72620 480 72648 3198
rect 73080 2922 73108 34054
rect 73724 30394 73752 34054
rect 73712 30388 73764 30394
rect 73712 30330 73764 30336
rect 73804 3324 73856 3330
rect 73804 3266 73856 3272
rect 73068 2916 73120 2922
rect 73068 2858 73120 2864
rect 73816 480 73844 3266
rect 74276 2990 74304 34054
rect 74368 34054 74520 34082
rect 75072 34054 75408 34082
rect 75624 34054 75776 34082
rect 76176 34054 76512 34082
rect 76728 34054 77064 34082
rect 74368 3126 74396 34054
rect 75380 30394 75408 34054
rect 74448 30388 74500 30394
rect 74448 30330 74500 30336
rect 75368 30388 75420 30394
rect 75368 30330 75420 30336
rect 74356 3120 74408 3126
rect 74356 3062 74408 3068
rect 74264 2984 74316 2990
rect 74264 2926 74316 2932
rect 74460 2854 74488 30330
rect 75000 4072 75052 4078
rect 75000 4014 75052 4020
rect 74448 2848 74500 2854
rect 74448 2790 74500 2796
rect 75012 480 75040 4014
rect 75748 3262 75776 34054
rect 76484 30394 76512 34054
rect 77036 31278 77064 34054
rect 77128 34054 77280 34082
rect 77832 34054 78168 34082
rect 78384 34054 78628 34082
rect 78936 34054 79272 34082
rect 79488 34054 79732 34082
rect 77024 31272 77076 31278
rect 77024 31214 77076 31220
rect 75828 30388 75880 30394
rect 75828 30330 75880 30336
rect 76472 30388 76524 30394
rect 76472 30330 76524 30336
rect 75736 3256 75788 3262
rect 75736 3198 75788 3204
rect 75840 3058 75868 30330
rect 77128 4146 77156 34054
rect 78140 30394 78168 34054
rect 78600 31210 78628 34054
rect 78588 31204 78640 31210
rect 78588 31146 78640 31152
rect 79244 30462 79272 34054
rect 79232 30456 79284 30462
rect 79232 30398 79284 30404
rect 79704 30394 79732 34054
rect 79796 34054 80040 34082
rect 80592 34054 81112 34082
rect 81236 34054 81388 34082
rect 81788 34054 82124 34082
rect 82340 34054 82768 34082
rect 82892 34054 83228 34082
rect 83444 34054 83872 34082
rect 83996 34054 84148 34082
rect 84548 34054 84884 34082
rect 85100 34054 85436 34082
rect 85652 34054 85988 34082
rect 86204 34054 86540 34082
rect 86756 34054 86908 34082
rect 87308 34054 87644 34082
rect 87860 34054 88196 34082
rect 88412 34054 88748 34082
rect 88964 34054 89300 34082
rect 89516 34054 89668 34082
rect 90068 34054 90404 34082
rect 90620 34054 90956 34082
rect 91172 34054 91508 34082
rect 91816 34054 92244 34082
rect 77208 30388 77260 30394
rect 77208 30330 77260 30336
rect 78128 30388 78180 30394
rect 78128 30330 78180 30336
rect 78588 30388 78640 30394
rect 78588 30330 78640 30336
rect 79692 30388 79744 30394
rect 79692 30330 79744 30336
rect 76196 4140 76248 4146
rect 76196 4082 76248 4088
rect 77116 4140 77168 4146
rect 77116 4082 77168 4088
rect 75828 3052 75880 3058
rect 75828 2994 75880 3000
rect 76208 480 76236 4082
rect 77220 3194 77248 30330
rect 77392 4004 77444 4010
rect 77392 3946 77444 3952
rect 77208 3188 77260 3194
rect 77208 3130 77260 3136
rect 77404 480 77432 3946
rect 78600 3482 78628 30330
rect 79692 3936 79744 3942
rect 79692 3878 79744 3884
rect 78600 3454 78720 3482
rect 78692 3398 78720 3454
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 78680 3392 78732 3398
rect 78680 3334 78732 3340
rect 78600 480 78628 3334
rect 79704 480 79732 3878
rect 79796 3641 79824 34054
rect 79876 30456 79928 30462
rect 79876 30398 79928 30404
rect 79888 4078 79916 30398
rect 79968 30388 80020 30394
rect 79968 30330 80020 30336
rect 79876 4072 79928 4078
rect 79876 4014 79928 4020
rect 79980 4010 80008 30330
rect 81084 26234 81112 34054
rect 81084 26206 81296 26234
rect 79968 4004 80020 4010
rect 79968 3946 80020 3952
rect 81268 3942 81296 26206
rect 81256 3936 81308 3942
rect 81256 3878 81308 3884
rect 81360 3874 81388 34054
rect 82096 31142 82124 34054
rect 82084 31136 82136 31142
rect 82084 31078 82136 31084
rect 80888 3868 80940 3874
rect 80888 3810 80940 3816
rect 81348 3868 81400 3874
rect 81348 3810 81400 3816
rect 79782 3632 79838 3641
rect 79782 3567 79838 3576
rect 80900 480 80928 3810
rect 82740 3806 82768 34054
rect 83200 31686 83228 34054
rect 83188 31680 83240 31686
rect 83188 31622 83240 31628
rect 83004 31068 83056 31074
rect 83004 31010 83056 31016
rect 83016 16574 83044 31010
rect 83844 26234 83872 34054
rect 83844 26206 84056 26234
rect 83016 16546 83320 16574
rect 82084 3800 82136 3806
rect 82084 3742 82136 3748
rect 82728 3800 82780 3806
rect 82728 3742 82780 3748
rect 82096 480 82124 3742
rect 83292 480 83320 16546
rect 84028 3505 84056 26206
rect 84014 3496 84070 3505
rect 84014 3431 84070 3440
rect 84120 3369 84148 34054
rect 84856 31346 84884 34054
rect 84844 31340 84896 31346
rect 84844 31282 84896 31288
rect 85408 31074 85436 34054
rect 85764 31612 85816 31618
rect 85764 31554 85816 31560
rect 85396 31068 85448 31074
rect 85396 31010 85448 31016
rect 85776 16574 85804 31554
rect 85960 30394 85988 34054
rect 86512 31482 86540 34054
rect 86500 31476 86552 31482
rect 86500 31418 86552 31424
rect 85948 30388 86000 30394
rect 85948 30330 86000 30336
rect 86776 30388 86828 30394
rect 86776 30330 86828 30336
rect 85776 16546 86448 16574
rect 84476 3664 84528 3670
rect 84476 3606 84528 3612
rect 84106 3360 84162 3369
rect 84106 3295 84162 3304
rect 84488 480 84516 3606
rect 85672 3528 85724 3534
rect 85672 3470 85724 3476
rect 85684 480 85712 3470
rect 86420 490 86448 16546
rect 86788 3534 86816 30330
rect 86880 3670 86908 34054
rect 87512 31544 87564 31550
rect 87512 31486 87564 31492
rect 87524 26234 87552 31486
rect 87616 30394 87644 34054
rect 88168 31754 88196 34054
rect 88156 31748 88208 31754
rect 88156 31690 88208 31696
rect 88720 30462 88748 34054
rect 88984 31408 89036 31414
rect 88984 31350 89036 31356
rect 88708 30456 88760 30462
rect 88708 30398 88760 30404
rect 87604 30388 87656 30394
rect 87604 30330 87656 30336
rect 88248 30388 88300 30394
rect 88248 30330 88300 30336
rect 87524 26206 87644 26234
rect 87616 3670 87644 26206
rect 88260 4622 88288 30330
rect 88248 4616 88300 4622
rect 88248 4558 88300 4564
rect 86868 3664 86920 3670
rect 86868 3606 86920 3612
rect 87604 3664 87656 3670
rect 87604 3606 87656 3612
rect 88996 3534 89024 31350
rect 89272 26234 89300 34054
rect 89640 30734 89668 34054
rect 90376 31686 90404 34054
rect 90272 31680 90324 31686
rect 90272 31622 90324 31628
rect 90364 31680 90416 31686
rect 90364 31622 90416 31628
rect 89628 30728 89680 30734
rect 89628 30670 89680 30676
rect 90284 26234 90312 31622
rect 90928 30870 90956 34054
rect 90916 30864 90968 30870
rect 90916 30806 90968 30812
rect 91480 30394 91508 34054
rect 92216 30546 92244 34054
rect 92308 34054 92368 34082
rect 92920 34054 93256 34082
rect 93472 34054 93716 34082
rect 94024 34054 94360 34082
rect 94576 34054 95004 34082
rect 92308 30938 92336 34054
rect 92296 30932 92348 30938
rect 92296 30874 92348 30880
rect 92216 30518 92428 30546
rect 91468 30388 91520 30394
rect 91468 30330 91520 30336
rect 92296 30388 92348 30394
rect 92296 30330 92348 30336
rect 89272 26206 89668 26234
rect 90284 26206 90404 26234
rect 89640 4690 89668 26206
rect 90376 16574 90404 26206
rect 90376 16546 90496 16574
rect 89628 4684 89680 4690
rect 89628 4626 89680 4632
rect 89168 3732 89220 3738
rect 89168 3674 89220 3680
rect 86776 3528 86828 3534
rect 86776 3470 86828 3476
rect 88984 3528 89036 3534
rect 88984 3470 89036 3476
rect 87972 3324 88024 3330
rect 87972 3266 88024 3272
rect 86696 598 86908 626
rect 86696 490 86724 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 462 86724 490
rect 86880 480 86908 598
rect 87984 480 88012 3266
rect 89180 480 89208 3674
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 90376 480 90404 3470
rect 90468 3330 90496 16546
rect 92308 4758 92336 30330
rect 92296 4752 92348 4758
rect 92296 4694 92348 4700
rect 92400 3466 92428 30518
rect 93124 30456 93176 30462
rect 93124 30398 93176 30404
rect 93136 3738 93164 30398
rect 93228 30394 93256 34054
rect 93688 31618 93716 34054
rect 93676 31612 93728 31618
rect 93676 31554 93728 31560
rect 94332 30394 94360 34054
rect 94504 31680 94556 31686
rect 94504 31622 94556 31628
rect 93216 30388 93268 30394
rect 93216 30330 93268 30336
rect 93768 30388 93820 30394
rect 93768 30330 93820 30336
rect 94320 30388 94372 30394
rect 94320 30330 94372 30336
rect 93780 5506 93808 30330
rect 93768 5500 93820 5506
rect 93768 5442 93820 5448
rect 93124 3732 93176 3738
rect 93124 3674 93176 3680
rect 94516 3602 94544 31622
rect 94872 30388 94924 30394
rect 94872 30330 94924 30336
rect 94884 26234 94912 30330
rect 94976 30138 95004 34054
rect 95114 33810 95142 34068
rect 95680 34054 96016 34082
rect 96232 34054 96476 34082
rect 96784 34054 97120 34082
rect 97336 34054 97672 34082
rect 95114 33782 95188 33810
rect 94976 30110 95096 30138
rect 94884 26206 95004 26234
rect 94976 5438 95004 26206
rect 94964 5432 95016 5438
rect 94964 5374 95016 5380
rect 95068 5370 95096 30110
rect 95056 5364 95108 5370
rect 95056 5306 95108 5312
rect 92756 3596 92808 3602
rect 92756 3538 92808 3544
rect 93952 3596 94004 3602
rect 93952 3538 94004 3544
rect 94504 3596 94556 3602
rect 94504 3538 94556 3544
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 92388 3460 92440 3466
rect 92388 3402 92440 3408
rect 90456 3324 90508 3330
rect 90456 3266 90508 3272
rect 91572 480 91600 3402
rect 92768 480 92796 3538
rect 93964 480 93992 3538
rect 95160 3074 95188 33782
rect 95884 31612 95936 31618
rect 95884 31554 95936 31560
rect 95160 3046 95280 3074
rect 95148 2916 95200 2922
rect 95148 2858 95200 2864
rect 95160 480 95188 2858
rect 95252 2786 95280 3046
rect 95896 2922 95924 31554
rect 95988 30394 96016 34054
rect 95976 30388 96028 30394
rect 95976 30330 96028 30336
rect 96448 5234 96476 34054
rect 97092 30462 97120 34054
rect 97080 30456 97132 30462
rect 97080 30398 97132 30404
rect 97644 30394 97672 34054
rect 97736 34054 97888 34082
rect 98440 34054 98776 34082
rect 98992 34054 99236 34082
rect 99544 34054 99880 34082
rect 100096 34054 100340 34082
rect 96528 30388 96580 30394
rect 96528 30330 96580 30336
rect 97632 30388 97684 30394
rect 97632 30330 97684 30336
rect 96540 5302 96568 30330
rect 96528 5296 96580 5302
rect 96528 5238 96580 5244
rect 96436 5228 96488 5234
rect 96436 5170 96488 5176
rect 97736 5098 97764 34054
rect 97908 30456 97960 30462
rect 97908 30398 97960 30404
rect 97816 30388 97868 30394
rect 97816 30330 97868 30336
rect 97828 5166 97856 30330
rect 97816 5160 97868 5166
rect 97816 5102 97868 5108
rect 97724 5092 97776 5098
rect 97724 5034 97776 5040
rect 97920 2990 97948 30398
rect 98748 30394 98776 34054
rect 98736 30388 98788 30394
rect 98736 30330 98788 30336
rect 99208 6322 99236 34054
rect 99852 30394 99880 34054
rect 100312 30462 100340 34054
rect 100496 34054 100648 34082
rect 101200 34054 101536 34082
rect 101752 34054 102088 34082
rect 102396 34054 102732 34082
rect 102948 34054 103376 34082
rect 100300 30456 100352 30462
rect 100300 30398 100352 30404
rect 99288 30388 99340 30394
rect 99288 30330 99340 30336
rect 99840 30388 99892 30394
rect 99840 30330 99892 30336
rect 99196 6316 99248 6322
rect 99196 6258 99248 6264
rect 98644 3120 98696 3126
rect 98644 3062 98696 3068
rect 97448 2984 97500 2990
rect 96356 2922 96568 2938
rect 97448 2926 97500 2932
rect 97908 2984 97960 2990
rect 97908 2926 97960 2932
rect 95884 2916 95936 2922
rect 95884 2858 95936 2864
rect 96344 2916 96568 2922
rect 96396 2910 96568 2916
rect 96344 2858 96396 2864
rect 96540 2854 96568 2910
rect 96252 2848 96304 2854
rect 96252 2790 96304 2796
rect 96528 2848 96580 2854
rect 96528 2790 96580 2796
rect 95240 2780 95292 2786
rect 95240 2722 95292 2728
rect 96264 480 96292 2790
rect 97460 480 97488 2926
rect 98656 480 98684 3062
rect 99300 2922 99328 30330
rect 100496 6254 100524 34054
rect 101404 31476 101456 31482
rect 101404 31418 101456 31424
rect 100668 30456 100720 30462
rect 100668 30398 100720 30404
rect 100576 30388 100628 30394
rect 100576 30330 100628 30336
rect 100484 6248 100536 6254
rect 100484 6190 100536 6196
rect 100588 5030 100616 30330
rect 100576 5024 100628 5030
rect 100576 4966 100628 4972
rect 100680 3058 100708 30398
rect 101416 3262 101444 31418
rect 101508 30394 101536 34054
rect 102060 30802 102088 34054
rect 102324 31272 102376 31278
rect 102324 31214 102376 31220
rect 102048 30796 102100 30802
rect 102048 30738 102100 30744
rect 101496 30388 101548 30394
rect 101496 30330 101548 30336
rect 102048 30388 102100 30394
rect 102048 30330 102100 30336
rect 102060 4962 102088 30330
rect 102336 16574 102364 31214
rect 102704 30394 102732 34054
rect 102692 30388 102744 30394
rect 102692 30330 102744 30336
rect 103244 30388 103296 30394
rect 103244 30330 103296 30336
rect 102336 16546 103192 16574
rect 102048 4956 102100 4962
rect 102048 4898 102100 4904
rect 103164 3482 103192 16546
rect 103256 5574 103284 30330
rect 103244 5568 103296 5574
rect 103244 5510 103296 5516
rect 103348 4894 103376 34054
rect 103440 34054 103500 34082
rect 104052 34054 104388 34082
rect 104604 34054 104848 34082
rect 105156 34054 105492 34082
rect 105708 34054 106044 34082
rect 103336 4888 103388 4894
rect 103336 4830 103388 4836
rect 103164 3454 103376 3482
rect 101036 3256 101088 3262
rect 101036 3198 101088 3204
rect 101404 3256 101456 3262
rect 101404 3198 101456 3204
rect 99840 3052 99892 3058
rect 99840 2994 99892 3000
rect 100668 3052 100720 3058
rect 100668 2994 100720 3000
rect 99288 2916 99340 2922
rect 99288 2858 99340 2864
rect 99852 480 99880 2994
rect 101048 480 101076 3198
rect 102232 3188 102284 3194
rect 102232 3130 102284 3136
rect 102244 480 102272 3130
rect 103348 480 103376 3454
rect 103440 3126 103468 34054
rect 104360 31550 104388 34054
rect 104348 31544 104400 31550
rect 104348 31486 104400 31492
rect 104164 31000 104216 31006
rect 104164 30942 104216 30948
rect 104176 3398 104204 30942
rect 104820 5642 104848 34054
rect 105464 30394 105492 34054
rect 106016 31482 106044 34054
rect 106108 34054 106260 34082
rect 106812 34054 107148 34082
rect 107364 34054 107608 34082
rect 107916 34054 108252 34082
rect 108468 34054 108896 34082
rect 106004 31476 106056 31482
rect 106004 31418 106056 31424
rect 105544 31340 105596 31346
rect 105544 31282 105596 31288
rect 105452 30388 105504 30394
rect 105452 30330 105504 30336
rect 105556 16574 105584 31282
rect 105556 16546 105860 16574
rect 104808 5636 104860 5642
rect 104808 5578 104860 5584
rect 104532 4140 104584 4146
rect 104532 4082 104584 4088
rect 104164 3392 104216 3398
rect 104164 3334 104216 3340
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 104544 480 104572 4082
rect 105832 3806 105860 16546
rect 106108 5778 106136 34054
rect 107120 30394 107148 34054
rect 107580 31414 107608 34054
rect 107568 31408 107620 31414
rect 107568 31350 107620 31356
rect 108224 30394 108252 34054
rect 108304 31136 108356 31142
rect 108304 31078 108356 31084
rect 106188 30388 106240 30394
rect 106188 30330 106240 30336
rect 107108 30388 107160 30394
rect 107108 30330 107160 30336
rect 107568 30388 107620 30394
rect 107568 30330 107620 30336
rect 108212 30388 108264 30394
rect 108212 30330 108264 30336
rect 106096 5772 106148 5778
rect 106096 5714 106148 5720
rect 106200 4826 106228 30330
rect 106188 4820 106240 4826
rect 106188 4762 106240 4768
rect 105728 3800 105780 3806
rect 105728 3742 105780 3748
rect 105820 3800 105872 3806
rect 105820 3742 105872 3748
rect 105740 480 105768 3742
rect 107580 3398 107608 30330
rect 108316 16574 108344 31078
rect 108316 16546 108436 16574
rect 108120 4072 108172 4078
rect 108120 4014 108172 4020
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 107568 3392 107620 3398
rect 107568 3334 107620 3340
rect 106936 480 106964 3334
rect 108132 480 108160 4014
rect 108408 3874 108436 16546
rect 108868 5846 108896 34054
rect 108960 34054 109020 34082
rect 109572 34054 110000 34082
rect 110124 34054 110368 34082
rect 110676 34054 111012 34082
rect 111228 34054 111656 34082
rect 108960 31686 108988 34054
rect 108948 31680 109000 31686
rect 108948 31622 109000 31628
rect 108948 30388 109000 30394
rect 108948 30330 109000 30336
rect 108856 5840 108908 5846
rect 108856 5782 108908 5788
rect 108960 5710 108988 30330
rect 109972 26234 110000 34054
rect 109972 26206 110276 26234
rect 110248 5914 110276 26206
rect 110236 5908 110288 5914
rect 110236 5850 110288 5856
rect 108948 5704 109000 5710
rect 108948 5646 109000 5652
rect 110340 4078 110368 34054
rect 110984 31006 111012 34054
rect 110972 31000 111024 31006
rect 110972 30942 111024 30948
rect 111628 6186 111656 34054
rect 111720 34054 111780 34082
rect 112332 34054 112668 34082
rect 112976 34054 113128 34082
rect 113528 34054 113864 34082
rect 114080 34054 114416 34082
rect 114632 34054 114968 34082
rect 115184 34054 115612 34082
rect 115736 34054 115888 34082
rect 116288 34054 116624 34082
rect 116840 34054 117268 34082
rect 117392 34054 117728 34082
rect 117944 34054 118280 34082
rect 118496 34054 118648 34082
rect 119048 34054 119384 34082
rect 119600 34054 120028 34082
rect 120152 34054 120488 34082
rect 120704 34054 121040 34082
rect 111616 6180 111668 6186
rect 111616 6122 111668 6128
rect 110328 4072 110380 4078
rect 110328 4014 110380 4020
rect 109316 4004 109368 4010
rect 109316 3946 109368 3952
rect 108396 3868 108448 3874
rect 108396 3810 108448 3816
rect 108212 3392 108264 3398
rect 108264 3340 108436 3346
rect 108212 3334 108436 3340
rect 108224 3318 108436 3334
rect 108408 3262 108436 3318
rect 108396 3256 108448 3262
rect 108396 3198 108448 3204
rect 109328 480 109356 3946
rect 111616 3936 111668 3942
rect 111616 3878 111668 3884
rect 110510 3632 110566 3641
rect 110510 3567 110566 3576
rect 110524 480 110552 3567
rect 111628 480 111656 3878
rect 111720 3346 111748 34054
rect 112640 31210 112668 34054
rect 112628 31204 112680 31210
rect 112628 31146 112680 31152
rect 113100 5982 113128 34054
rect 113836 30394 113864 34054
rect 114388 31278 114416 34054
rect 114376 31272 114428 31278
rect 114376 31214 114428 31220
rect 114940 30394 114968 34054
rect 113824 30388 113876 30394
rect 113824 30330 113876 30336
rect 114468 30388 114520 30394
rect 114468 30330 114520 30336
rect 114928 30388 114980 30394
rect 114928 30330 114980 30336
rect 115480 30388 115532 30394
rect 115480 30330 115532 30336
rect 114480 6050 114508 30330
rect 115492 26234 115520 30330
rect 115584 30138 115612 34054
rect 115860 31142 115888 34054
rect 115848 31136 115900 31142
rect 115848 31078 115900 31084
rect 116596 30394 116624 34054
rect 116584 30388 116636 30394
rect 116584 30330 116636 30336
rect 117136 30388 117188 30394
rect 117136 30330 117188 30336
rect 115584 30110 115888 30138
rect 115492 26206 115796 26234
rect 115768 6118 115796 26206
rect 115756 6112 115808 6118
rect 115756 6054 115808 6060
rect 114468 6044 114520 6050
rect 114468 5986 114520 5992
rect 113088 5976 113140 5982
rect 113088 5918 113140 5924
rect 112812 4140 112864 4146
rect 112812 4082 112864 4088
rect 111720 3318 112116 3346
rect 112088 3262 112116 3318
rect 112076 3256 112128 3262
rect 112076 3198 112128 3204
rect 112824 480 112852 4082
rect 115860 4078 115888 30110
rect 117148 6798 117176 30330
rect 117136 6792 117188 6798
rect 117136 6734 117188 6740
rect 117240 4214 117268 34054
rect 117700 30666 117728 34054
rect 117688 30660 117740 30666
rect 117688 30602 117740 30608
rect 118252 26234 118280 34054
rect 118252 26206 118556 26234
rect 118528 6730 118556 26206
rect 118516 6724 118568 6730
rect 118516 6666 118568 6672
rect 117228 4208 117280 4214
rect 117228 4150 117280 4156
rect 114008 4072 114060 4078
rect 114008 4014 114060 4020
rect 115848 4072 115900 4078
rect 115848 4014 115900 4020
rect 114020 480 114048 4014
rect 118620 3874 118648 34054
rect 119356 31346 119384 34054
rect 119344 31340 119396 31346
rect 119344 31282 119396 31288
rect 119344 31068 119396 31074
rect 119344 31010 119396 31016
rect 118608 3868 118660 3874
rect 118608 3810 118660 3816
rect 119356 3534 119384 31010
rect 120000 6662 120028 34054
rect 120460 30394 120488 34054
rect 121012 31074 121040 34054
rect 121242 33810 121270 34068
rect 121808 34054 122144 34082
rect 122360 34054 122696 34082
rect 122912 34054 123248 34082
rect 123556 34054 123892 34082
rect 121242 33782 121316 33810
rect 121000 31068 121052 31074
rect 121000 31010 121052 31016
rect 120448 30388 120500 30394
rect 120448 30330 120500 30336
rect 119988 6656 120040 6662
rect 119988 6598 120040 6604
rect 121288 6594 121316 33782
rect 122116 30394 122144 34054
rect 121368 30388 121420 30394
rect 121368 30330 121420 30336
rect 122104 30388 122156 30394
rect 122104 30330 122156 30336
rect 121276 6588 121328 6594
rect 121276 6530 121328 6536
rect 119896 4140 119948 4146
rect 119896 4082 119948 4088
rect 119344 3528 119396 3534
rect 117594 3496 117650 3505
rect 119344 3470 119396 3476
rect 117594 3431 117650 3440
rect 115204 3392 115256 3398
rect 115204 3334 115256 3340
rect 115216 480 115244 3334
rect 116400 3324 116452 3330
rect 116400 3266 116452 3272
rect 116412 480 116440 3266
rect 117608 480 117636 3431
rect 118790 3360 118846 3369
rect 118790 3295 118846 3304
rect 118804 480 118832 3295
rect 119908 480 119936 4082
rect 121380 4078 121408 30330
rect 122668 4282 122696 34054
rect 123220 30394 123248 34054
rect 123864 30462 123892 34054
rect 124048 34054 124108 34082
rect 124660 34054 124996 34082
rect 125212 34054 125548 34082
rect 125764 34054 126100 34082
rect 126316 34054 126744 34082
rect 123852 30456 123904 30462
rect 123852 30398 123904 30404
rect 122748 30388 122800 30394
rect 122748 30330 122800 30336
rect 123208 30388 123260 30394
rect 123208 30330 123260 30336
rect 123944 30388 123996 30394
rect 123944 30330 123996 30336
rect 122656 4276 122708 4282
rect 122656 4218 122708 4224
rect 121368 4072 121420 4078
rect 121368 4014 121420 4020
rect 122760 4010 122788 30330
rect 123956 8226 123984 30330
rect 123944 8220 123996 8226
rect 123944 8162 123996 8168
rect 124048 4486 124076 34054
rect 124128 30456 124180 30462
rect 124128 30398 124180 30404
rect 124036 4480 124088 4486
rect 124036 4422 124088 4428
rect 122748 4004 122800 4010
rect 122748 3946 122800 3952
rect 124140 3942 124168 30398
rect 124968 30394 124996 34054
rect 124956 30388 125008 30394
rect 124956 30330 125008 30336
rect 125416 30388 125468 30394
rect 125416 30330 125468 30336
rect 125428 8158 125456 30330
rect 125416 8152 125468 8158
rect 125416 8094 125468 8100
rect 123484 3936 123536 3942
rect 123484 3878 123536 3884
rect 124128 3936 124180 3942
rect 124128 3878 124180 3884
rect 122288 3664 122340 3670
rect 122288 3606 122340 3612
rect 121092 3528 121144 3534
rect 121092 3470 121144 3476
rect 121104 480 121132 3470
rect 122300 480 122328 3606
rect 123496 480 123524 3878
rect 125520 3806 125548 34054
rect 126072 30394 126100 34054
rect 126060 30388 126112 30394
rect 126060 30330 126112 30336
rect 126716 8090 126744 34054
rect 126854 33810 126882 34068
rect 127420 34054 127756 34082
rect 127972 34054 128308 34082
rect 128524 34054 128860 34082
rect 129076 34054 129412 34082
rect 126854 33782 126928 33810
rect 126796 30388 126848 30394
rect 126796 30330 126848 30336
rect 126704 8084 126756 8090
rect 126704 8026 126756 8032
rect 125876 4616 125928 4622
rect 125876 4558 125928 4564
rect 124680 3800 124732 3806
rect 124680 3742 124732 3748
rect 125508 3800 125560 3806
rect 125508 3742 125560 3748
rect 124692 480 124720 3742
rect 125888 480 125916 4558
rect 126808 4418 126836 30330
rect 126796 4412 126848 4418
rect 126796 4354 126848 4360
rect 126900 3670 126928 33782
rect 127164 31748 127216 31754
rect 127164 31690 127216 31696
rect 127176 6914 127204 31690
rect 127728 30394 127756 34054
rect 128280 30666 128308 34054
rect 128268 30660 128320 30666
rect 128268 30602 128320 30608
rect 128832 30462 128860 34054
rect 128820 30456 128872 30462
rect 128820 30398 128872 30404
rect 129384 30394 129412 34054
rect 129476 34054 129628 34082
rect 130180 34054 130516 34082
rect 130732 34054 130976 34082
rect 131284 34054 131620 34082
rect 131836 34054 132172 34082
rect 127716 30388 127768 30394
rect 127716 30330 127768 30336
rect 128268 30388 128320 30394
rect 128268 30330 128320 30336
rect 129372 30388 129424 30394
rect 129372 30330 129424 30336
rect 126992 6886 127204 6914
rect 126888 3664 126940 3670
rect 126888 3606 126940 3612
rect 126992 480 127020 6886
rect 128280 4214 128308 30330
rect 129476 7954 129504 34054
rect 129740 30728 129792 30734
rect 129740 30670 129792 30676
rect 129648 30456 129700 30462
rect 129648 30398 129700 30404
rect 129556 30388 129608 30394
rect 129556 30330 129608 30336
rect 129464 7948 129516 7954
rect 129464 7890 129516 7896
rect 129372 4684 129424 4690
rect 129372 4626 129424 4632
rect 128268 4208 128320 4214
rect 128268 4150 128320 4156
rect 127440 3936 127492 3942
rect 127492 3884 127848 3890
rect 127440 3878 127848 3884
rect 127452 3862 127848 3878
rect 127820 3806 127848 3862
rect 127808 3800 127860 3806
rect 127808 3742 127860 3748
rect 128176 3732 128228 3738
rect 128176 3674 128228 3680
rect 128188 480 128216 3674
rect 129384 480 129412 4626
rect 129568 4350 129596 30330
rect 129556 4344 129608 4350
rect 129556 4286 129608 4292
rect 129660 3670 129688 30398
rect 129752 16574 129780 30670
rect 130488 30394 130516 34054
rect 130476 30388 130528 30394
rect 130476 30330 130528 30336
rect 129752 16546 130608 16574
rect 129648 3664 129700 3670
rect 129648 3606 129700 3612
rect 130580 480 130608 16546
rect 130948 4554 130976 34054
rect 131592 30394 131620 34054
rect 132144 30462 132172 34054
rect 132328 34054 132388 34082
rect 132940 34054 133276 34082
rect 133492 34054 133828 34082
rect 134136 34054 134472 34082
rect 134688 34054 135024 34082
rect 132132 30456 132184 30462
rect 132132 30398 132184 30404
rect 131028 30388 131080 30394
rect 131028 30330 131080 30336
rect 131580 30388 131632 30394
rect 131580 30330 131632 30336
rect 132224 30388 132276 30394
rect 132224 30330 132276 30336
rect 130936 4548 130988 4554
rect 130936 4490 130988 4496
rect 131040 3777 131068 30330
rect 132236 8022 132264 30330
rect 132224 8016 132276 8022
rect 132224 7958 132276 7964
rect 132328 4622 132356 34054
rect 132500 30864 132552 30870
rect 132500 30806 132552 30812
rect 132408 30456 132460 30462
rect 132408 30398 132460 30404
rect 132316 4616 132368 4622
rect 132316 4558 132368 4564
rect 131026 3768 131082 3777
rect 131026 3703 131082 3712
rect 131764 3596 131816 3602
rect 131764 3538 131816 3544
rect 131776 480 131804 3538
rect 132420 3534 132448 30398
rect 132512 16574 132540 30806
rect 133248 30394 133276 34054
rect 133236 30388 133288 30394
rect 133236 30330 133288 30336
rect 133696 30388 133748 30394
rect 133696 30330 133748 30336
rect 132512 16546 133000 16574
rect 132408 3528 132460 3534
rect 132408 3470 132460 3476
rect 132972 480 133000 16546
rect 133708 7886 133736 30330
rect 133696 7880 133748 7886
rect 133696 7822 133748 7828
rect 133800 3641 133828 34054
rect 134444 30394 134472 34054
rect 134432 30388 134484 30394
rect 134432 30330 134484 30336
rect 134996 7818 135024 34054
rect 135180 34054 135240 34082
rect 135792 34054 136128 34082
rect 136344 34054 136588 34082
rect 136896 34054 137232 34082
rect 137448 34054 137876 34082
rect 135076 30388 135128 30394
rect 135076 30330 135128 30336
rect 134984 7812 135036 7818
rect 134984 7754 135036 7760
rect 134156 4752 134208 4758
rect 134156 4694 134208 4700
rect 133786 3632 133842 3641
rect 133786 3567 133842 3576
rect 134168 480 134196 4694
rect 135088 4690 135116 30330
rect 135076 4684 135128 4690
rect 135076 4626 135128 4632
rect 135180 3505 135208 34054
rect 135444 30932 135496 30938
rect 135444 30874 135496 30880
rect 135456 16574 135484 30874
rect 136100 30394 136128 34054
rect 136560 30734 136588 34054
rect 136548 30728 136600 30734
rect 136548 30670 136600 30676
rect 137204 30394 137232 34054
rect 136088 30388 136140 30394
rect 136088 30330 136140 30336
rect 136548 30388 136600 30394
rect 136548 30330 136600 30336
rect 137192 30388 137244 30394
rect 137192 30330 137244 30336
rect 135456 16546 136496 16574
rect 135166 3496 135222 3505
rect 135166 3431 135222 3440
rect 135260 3460 135312 3466
rect 135260 3402 135312 3408
rect 135272 480 135300 3402
rect 136468 480 136496 16546
rect 136560 4758 136588 30330
rect 137848 5506 137876 34054
rect 137940 34054 138000 34082
rect 138552 34054 138980 34082
rect 139104 34054 139348 34082
rect 139656 34054 139992 34082
rect 140208 34054 140544 34082
rect 137940 30870 137968 34054
rect 137928 30864 137980 30870
rect 137928 30806 137980 30812
rect 137928 30388 137980 30394
rect 137928 30330 137980 30336
rect 137652 5500 137704 5506
rect 137652 5442 137704 5448
rect 137836 5500 137888 5506
rect 137836 5442 137888 5448
rect 136548 4752 136600 4758
rect 136548 4694 136600 4700
rect 137664 480 137692 5442
rect 137940 3466 137968 30330
rect 138952 26234 138980 34054
rect 138952 26206 139256 26234
rect 139228 7750 139256 26206
rect 139216 7744 139268 7750
rect 139216 7686 139268 7692
rect 139320 5137 139348 34054
rect 139964 30598 139992 34054
rect 139952 30592 140004 30598
rect 139952 30534 140004 30540
rect 140516 30394 140544 34054
rect 140608 34054 140760 34082
rect 141312 34054 141648 34082
rect 141864 34054 142016 34082
rect 142416 34054 142752 34082
rect 142968 34054 143396 34082
rect 140504 30388 140556 30394
rect 140504 30330 140556 30336
rect 140608 5438 140636 34054
rect 141620 30394 141648 34054
rect 140688 30388 140740 30394
rect 140688 30330 140740 30336
rect 141608 30388 141660 30394
rect 141608 30330 141660 30336
rect 140044 5432 140096 5438
rect 140044 5374 140096 5380
rect 140596 5432 140648 5438
rect 140596 5374 140648 5380
rect 139306 5128 139362 5137
rect 139306 5063 139362 5072
rect 137928 3460 137980 3466
rect 137928 3402 137980 3408
rect 138848 2848 138900 2854
rect 138848 2790 138900 2796
rect 138860 480 138888 2790
rect 140056 480 140084 5374
rect 140700 3369 140728 30330
rect 141988 7682 142016 34054
rect 142724 30394 142752 34054
rect 142804 30796 142856 30802
rect 142804 30738 142856 30744
rect 142068 30388 142120 30394
rect 142068 30330 142120 30336
rect 142712 30388 142764 30394
rect 142712 30330 142764 30336
rect 141976 7676 142028 7682
rect 141976 7618 142028 7624
rect 142080 6866 142108 30330
rect 142068 6860 142120 6866
rect 142068 6802 142120 6808
rect 141240 5364 141292 5370
rect 141240 5306 141292 5312
rect 140686 3360 140742 3369
rect 140686 3295 140742 3304
rect 141252 480 141280 5306
rect 142816 2922 142844 30738
rect 143264 30388 143316 30394
rect 143264 30330 143316 30336
rect 143276 7614 143304 30330
rect 143264 7608 143316 7614
rect 143264 7550 143316 7556
rect 143368 6526 143396 34054
rect 143460 34054 143520 34082
rect 144072 34054 144408 34082
rect 143460 30394 143488 34054
rect 144380 30394 144408 34054
rect 144702 33810 144730 34068
rect 145268 34054 145604 34082
rect 145820 34054 146248 34082
rect 146372 34054 146708 34082
rect 146924 34054 147352 34082
rect 147476 34054 147628 34082
rect 148028 34054 148364 34082
rect 148580 34054 148916 34082
rect 149132 34054 149468 34082
rect 149684 34054 150020 34082
rect 144702 33782 144776 33810
rect 143448 30388 143500 30394
rect 143448 30330 143500 30336
rect 144368 30388 144420 30394
rect 144368 30330 144420 30336
rect 143448 30252 143500 30258
rect 143448 30194 143500 30200
rect 143356 6520 143408 6526
rect 143356 6462 143408 6468
rect 143460 5370 143488 30194
rect 144748 6458 144776 33782
rect 145576 30394 145604 34054
rect 144828 30388 144880 30394
rect 144828 30330 144880 30336
rect 145564 30388 145616 30394
rect 145564 30330 145616 30336
rect 146116 30388 146168 30394
rect 146116 30330 146168 30336
rect 144736 6452 144788 6458
rect 144736 6394 144788 6400
rect 143448 5364 143500 5370
rect 143448 5306 143500 5312
rect 144840 5302 144868 30330
rect 146128 8498 146156 30330
rect 146116 8492 146168 8498
rect 146116 8434 146168 8440
rect 143540 5296 143592 5302
rect 143540 5238 143592 5244
rect 144828 5296 144880 5302
rect 144828 5238 144880 5244
rect 142436 2916 142488 2922
rect 142436 2858 142488 2864
rect 142804 2916 142856 2922
rect 142804 2858 142856 2864
rect 142448 480 142476 2858
rect 143552 480 143580 5238
rect 146220 5234 146248 34054
rect 146680 30394 146708 34054
rect 146668 30388 146720 30394
rect 146668 30330 146720 30336
rect 147324 26234 147352 34054
rect 147496 30388 147548 30394
rect 147496 30330 147548 30336
rect 147324 26206 147444 26234
rect 147416 8566 147444 26206
rect 147404 8560 147456 8566
rect 147404 8502 147456 8508
rect 147508 6390 147536 30330
rect 147496 6384 147548 6390
rect 147496 6326 147548 6332
rect 144736 5228 144788 5234
rect 144736 5170 144788 5176
rect 146208 5228 146260 5234
rect 146208 5170 146260 5176
rect 144748 480 144776 5170
rect 147600 5166 147628 34054
rect 148336 30394 148364 34054
rect 148324 30388 148376 30394
rect 148324 30330 148376 30336
rect 148888 8634 148916 34054
rect 149440 30462 149468 34054
rect 149428 30456 149480 30462
rect 149428 30398 149480 30404
rect 149992 30394 150020 34054
rect 150176 34054 150236 34082
rect 150788 34054 151124 34082
rect 151340 34054 151676 34082
rect 151892 34054 152228 34082
rect 152444 34054 152780 34082
rect 148968 30388 149020 30394
rect 148968 30330 149020 30336
rect 149980 30388 150032 30394
rect 149980 30330 150032 30336
rect 148876 8628 148928 8634
rect 148876 8570 148928 8576
rect 148980 6633 149008 30330
rect 150176 8702 150204 34054
rect 150348 30456 150400 30462
rect 150348 30398 150400 30404
rect 150256 30388 150308 30394
rect 150256 30330 150308 30336
rect 150164 8696 150216 8702
rect 150164 8638 150216 8644
rect 148966 6624 149022 6633
rect 148966 6559 149022 6568
rect 150268 6497 150296 30330
rect 150254 6488 150310 6497
rect 150254 6423 150310 6432
rect 147128 5160 147180 5166
rect 147128 5102 147180 5108
rect 147588 5160 147640 5166
rect 147588 5102 147640 5108
rect 145932 2984 145984 2990
rect 145932 2926 145984 2932
rect 145944 480 145972 2926
rect 147140 480 147168 5102
rect 150360 5098 150388 30398
rect 151096 30394 151124 34054
rect 151084 30388 151136 30394
rect 151084 30330 151136 30336
rect 151648 6322 151676 34054
rect 152200 30394 152228 34054
rect 152752 30462 152780 34054
rect 152982 33810 153010 34068
rect 153548 34054 153884 34082
rect 154100 34054 154528 34082
rect 154652 34054 154988 34082
rect 155296 34054 155724 34082
rect 152982 33782 153056 33810
rect 152740 30456 152792 30462
rect 152740 30398 152792 30404
rect 151728 30388 151780 30394
rect 151728 30330 151780 30336
rect 152188 30388 152240 30394
rect 152188 30330 152240 30336
rect 152924 30388 152976 30394
rect 152924 30330 152976 30336
rect 150624 6316 150676 6322
rect 150624 6258 150676 6264
rect 151636 6316 151688 6322
rect 151636 6258 151688 6264
rect 148324 5092 148376 5098
rect 148324 5034 148376 5040
rect 150348 5092 150400 5098
rect 150348 5034 150400 5040
rect 148336 480 148364 5034
rect 149520 3052 149572 3058
rect 149520 2994 149572 3000
rect 149532 480 149560 2994
rect 150636 480 150664 6258
rect 151740 5001 151768 30330
rect 152936 8770 152964 30330
rect 152924 8764 152976 8770
rect 152924 8706 152976 8712
rect 153028 6361 153056 33782
rect 153108 30456 153160 30462
rect 153108 30398 153160 30404
rect 153014 6352 153070 6361
rect 153014 6287 153070 6296
rect 153120 5030 153148 30398
rect 153856 30394 153884 34054
rect 153844 30388 153896 30394
rect 153844 30330 153896 30336
rect 154396 30388 154448 30394
rect 154396 30330 154448 30336
rect 154408 8838 154436 30330
rect 154396 8832 154448 8838
rect 154396 8774 154448 8780
rect 154212 6248 154264 6254
rect 154212 6190 154264 6196
rect 151820 5024 151872 5030
rect 151726 4992 151782 5001
rect 151820 4966 151872 4972
rect 153108 5024 153160 5030
rect 153108 4966 153160 4972
rect 151726 4927 151782 4936
rect 151832 480 151860 4966
rect 153016 3120 153068 3126
rect 153016 3062 153068 3068
rect 153028 480 153056 3062
rect 154224 480 154252 6190
rect 154500 4865 154528 34054
rect 154960 30394 154988 34054
rect 155224 31544 155276 31550
rect 155224 31486 155276 31492
rect 154948 30388 155000 30394
rect 154948 30330 155000 30336
rect 154486 4856 154542 4865
rect 154486 4791 154542 4800
rect 155236 3126 155264 31486
rect 155696 8906 155724 34054
rect 155834 33810 155862 34068
rect 156400 34054 156736 34082
rect 156952 34054 157196 34082
rect 157504 34054 157840 34082
rect 158056 34054 158392 34082
rect 155834 33782 155908 33810
rect 155776 30388 155828 30394
rect 155776 30330 155828 30336
rect 155684 8900 155736 8906
rect 155684 8842 155736 8848
rect 155788 6254 155816 30330
rect 155776 6248 155828 6254
rect 155776 6190 155828 6196
rect 155880 4962 155908 33782
rect 156604 31476 156656 31482
rect 156604 31418 156656 31424
rect 155408 4956 155460 4962
rect 155408 4898 155460 4904
rect 155868 4956 155920 4962
rect 155868 4898 155920 4904
rect 155224 3120 155276 3126
rect 155224 3062 155276 3068
rect 155420 480 155448 4898
rect 156616 3058 156644 31418
rect 156708 30394 156736 34054
rect 156696 30388 156748 30394
rect 156696 30330 156748 30336
rect 157168 9654 157196 34054
rect 157812 30394 157840 34054
rect 157984 31612 158036 31618
rect 157984 31554 158036 31560
rect 157248 30388 157300 30394
rect 157248 30330 157300 30336
rect 157800 30388 157852 30394
rect 157800 30330 157852 30336
rect 157156 9648 157208 9654
rect 157156 9590 157208 9596
rect 157260 6225 157288 30330
rect 157246 6216 157302 6225
rect 157246 6151 157302 6160
rect 157800 5568 157852 5574
rect 157800 5510 157852 5516
rect 156604 3052 156656 3058
rect 156604 2994 156656 3000
rect 156604 2916 156656 2922
rect 156604 2858 156656 2864
rect 156616 480 156644 2858
rect 157812 480 157840 5510
rect 157996 2922 158024 31554
rect 158364 30462 158392 34054
rect 158548 34054 158608 34082
rect 159160 34054 159496 34082
rect 159712 34054 160048 34082
rect 160264 34054 160600 34082
rect 160816 34054 161152 34082
rect 158352 30456 158404 30462
rect 158352 30398 158404 30404
rect 158444 30388 158496 30394
rect 158444 30330 158496 30336
rect 158456 13462 158484 30330
rect 158444 13456 158496 13462
rect 158444 13398 158496 13404
rect 158548 9586 158576 34054
rect 159364 31680 159416 31686
rect 159364 31622 159416 31628
rect 158628 30456 158680 30462
rect 158628 30398 158680 30404
rect 158536 9580 158588 9586
rect 158536 9522 158588 9528
rect 158640 7002 158668 30398
rect 158628 6996 158680 7002
rect 158628 6938 158680 6944
rect 158904 4888 158956 4894
rect 158904 4830 158956 4836
rect 157984 2916 158036 2922
rect 157984 2858 158036 2864
rect 158916 480 158944 4830
rect 159376 2854 159404 31622
rect 159468 30394 159496 34054
rect 159456 30388 159508 30394
rect 159456 30330 159508 30336
rect 159916 30388 159968 30394
rect 159916 30330 159968 30336
rect 159928 13394 159956 30330
rect 159916 13388 159968 13394
rect 159916 13330 159968 13336
rect 160020 9518 160048 34054
rect 160572 30394 160600 34054
rect 160744 31000 160796 31006
rect 160744 30942 160796 30948
rect 160560 30388 160612 30394
rect 160560 30330 160612 30336
rect 160008 9512 160060 9518
rect 160008 9454 160060 9460
rect 160756 3194 160784 30942
rect 161124 30462 161152 34054
rect 161308 34054 161368 34082
rect 161920 34054 162256 34082
rect 162472 34054 162808 34082
rect 163024 34054 163360 34082
rect 163576 34054 163912 34082
rect 161112 30456 161164 30462
rect 161112 30398 161164 30404
rect 161204 30388 161256 30394
rect 161204 30330 161256 30336
rect 161216 9450 161244 30330
rect 161204 9444 161256 9450
rect 161204 9386 161256 9392
rect 161308 9314 161336 34054
rect 162228 31686 162256 34054
rect 162216 31680 162268 31686
rect 162216 31622 162268 31628
rect 161388 30456 161440 30462
rect 161388 30398 161440 30404
rect 161296 9308 161348 9314
rect 161296 9250 161348 9256
rect 161400 4894 161428 30398
rect 162780 13326 162808 34054
rect 163332 30462 163360 34054
rect 163320 30456 163372 30462
rect 163320 30398 163372 30404
rect 163884 30394 163912 34054
rect 163976 34054 164128 34082
rect 164680 34054 165016 34082
rect 165232 34054 165476 34082
rect 165876 34054 166212 34082
rect 166428 34054 166856 34082
rect 163872 30388 163924 30394
rect 163872 30330 163924 30336
rect 162768 13320 162820 13326
rect 162768 13262 162820 13268
rect 163976 13258 164004 34054
rect 164148 30456 164200 30462
rect 164148 30398 164200 30404
rect 164056 30388 164108 30394
rect 164056 30330 164108 30336
rect 163964 13252 164016 13258
rect 163964 13194 164016 13200
rect 164068 11150 164096 30330
rect 164056 11144 164108 11150
rect 164056 11086 164108 11092
rect 164160 9382 164188 30398
rect 164988 30394 165016 34054
rect 165448 30462 165476 34054
rect 165436 30456 165488 30462
rect 165436 30398 165488 30404
rect 166184 30394 166212 34054
rect 166264 31204 166316 31210
rect 166264 31146 166316 31152
rect 164976 30388 165028 30394
rect 164976 30330 165028 30336
rect 165528 30388 165580 30394
rect 165528 30330 165580 30336
rect 166172 30388 166224 30394
rect 166172 30330 166224 30336
rect 164148 9376 164200 9382
rect 164148 9318 164200 9324
rect 165540 9246 165568 30330
rect 165528 9240 165580 9246
rect 165528 9182 165580 9188
rect 166080 5772 166132 5778
rect 166080 5714 166132 5720
rect 162492 5636 162544 5642
rect 162492 5578 162544 5584
rect 161388 4888 161440 4894
rect 161388 4830 161440 4836
rect 160100 3188 160152 3194
rect 160100 3130 160152 3136
rect 160744 3188 160796 3194
rect 160744 3130 160796 3136
rect 159364 2848 159416 2854
rect 159364 2790 159416 2796
rect 160112 480 160140 3130
rect 161296 3120 161348 3126
rect 161296 3062 161348 3068
rect 161308 480 161336 3062
rect 162504 480 162532 5578
rect 163688 4820 163740 4826
rect 163688 4762 163740 4768
rect 163700 480 163728 4762
rect 164884 3052 164936 3058
rect 164884 2994 164936 3000
rect 164896 480 164924 2994
rect 166092 480 166120 5714
rect 166276 2990 166304 31146
rect 166828 9178 166856 34054
rect 166920 34054 166980 34082
rect 167532 34054 167960 34082
rect 168084 34054 168328 34082
rect 168636 34054 168972 34082
rect 169188 34054 169616 34082
rect 166920 31550 166948 34054
rect 166908 31544 166960 31550
rect 166908 31486 166960 31492
rect 167644 31272 167696 31278
rect 167644 31214 167696 31220
rect 166908 30388 166960 30394
rect 166908 30330 166960 30336
rect 166816 9172 166868 9178
rect 166816 9114 166868 9120
rect 166920 4826 166948 30330
rect 166908 4820 166960 4826
rect 166908 4762 166960 4768
rect 167184 3256 167236 3262
rect 167184 3198 167236 3204
rect 166264 2984 166316 2990
rect 166264 2926 166316 2932
rect 167196 480 167224 3198
rect 167656 3058 167684 31214
rect 167932 26234 167960 34054
rect 167932 26206 168236 26234
rect 168208 12510 168236 26206
rect 168196 12504 168248 12510
rect 168196 12446 168248 12452
rect 168300 9042 168328 34054
rect 168944 31482 168972 34054
rect 168932 31476 168984 31482
rect 168932 31418 168984 31424
rect 169024 31136 169076 31142
rect 169024 31078 169076 31084
rect 168288 9036 168340 9042
rect 168288 8978 168340 8984
rect 167644 3052 167696 3058
rect 167644 2994 167696 3000
rect 169036 2922 169064 31078
rect 169588 13190 169616 34054
rect 169680 34054 169740 34082
rect 170292 34054 170628 34082
rect 170844 34054 171088 34082
rect 171396 34054 171732 34082
rect 171948 34054 172284 34082
rect 169576 13184 169628 13190
rect 169576 13126 169628 13132
rect 169680 8974 169708 34054
rect 170404 31408 170456 31414
rect 170404 31350 170456 31356
rect 169668 8968 169720 8974
rect 169668 8910 169720 8916
rect 169576 5704 169628 5710
rect 169576 5646 169628 5652
rect 168380 2916 168432 2922
rect 168380 2858 168432 2864
rect 169024 2916 169076 2922
rect 169024 2858 169076 2864
rect 168392 480 168420 2858
rect 169588 480 169616 5646
rect 170416 3194 170444 31350
rect 170600 30462 170628 34054
rect 170588 30456 170640 30462
rect 170588 30398 170640 30404
rect 171060 13122 171088 34054
rect 171704 30530 171732 34054
rect 172256 30802 172284 34054
rect 172348 34054 172500 34082
rect 173052 34054 173388 34082
rect 173604 34054 173756 34082
rect 174156 34054 174492 34082
rect 174708 34054 175136 34082
rect 172244 30796 172296 30802
rect 172244 30738 172296 30744
rect 171692 30524 171744 30530
rect 171692 30466 171744 30472
rect 171048 13116 171100 13122
rect 171048 13058 171100 13064
rect 172348 12646 172376 34054
rect 173164 31340 173216 31346
rect 173164 31282 173216 31288
rect 172428 30524 172480 30530
rect 172428 30466 172480 30472
rect 172336 12640 172388 12646
rect 172336 12582 172388 12588
rect 172440 8362 172468 30466
rect 173176 16574 173204 31282
rect 173360 30530 173388 34054
rect 173348 30524 173400 30530
rect 173348 30466 173400 30472
rect 173176 16546 173296 16574
rect 172428 8356 172480 8362
rect 172428 8298 172480 8304
rect 173164 5908 173216 5914
rect 173164 5850 173216 5856
rect 170772 5840 170824 5846
rect 170772 5782 170824 5788
rect 170404 3188 170456 3194
rect 170404 3130 170456 3136
rect 170784 480 170812 5782
rect 171968 2848 172020 2854
rect 171968 2790 172020 2796
rect 171980 480 172008 2790
rect 173176 480 173204 5850
rect 173268 2854 173296 16546
rect 173728 13870 173756 34054
rect 174464 30530 174492 34054
rect 173808 30524 173860 30530
rect 173808 30466 173860 30472
rect 174452 30524 174504 30530
rect 174452 30466 174504 30472
rect 175004 30524 175056 30530
rect 175004 30466 175056 30472
rect 173716 13864 173768 13870
rect 173716 13806 173768 13812
rect 173820 9110 173848 30466
rect 175016 26234 175044 30466
rect 175108 30138 175136 34054
rect 175200 34054 175260 34082
rect 175812 34054 176148 34082
rect 176456 34054 176608 34082
rect 177008 34054 177344 34082
rect 177560 34054 177988 34082
rect 178112 34054 178448 34082
rect 178664 34054 179000 34082
rect 179216 34054 179368 34082
rect 179768 34054 180104 34082
rect 180320 34054 180564 34082
rect 180872 34054 181208 34082
rect 181424 34054 181760 34082
rect 175200 30734 175228 34054
rect 175924 31068 175976 31074
rect 175924 31010 175976 31016
rect 175188 30728 175240 30734
rect 175188 30670 175240 30676
rect 175108 30110 175228 30138
rect 175016 26206 175136 26234
rect 175108 12578 175136 26206
rect 175096 12572 175148 12578
rect 175096 12514 175148 12520
rect 173808 9104 173860 9110
rect 173808 9046 173860 9052
rect 175200 8430 175228 30110
rect 175188 8424 175240 8430
rect 175188 8366 175240 8372
rect 175936 3330 175964 31010
rect 176120 26234 176148 34054
rect 176120 26206 176516 26234
rect 176488 12714 176516 26206
rect 176476 12708 176528 12714
rect 176476 12650 176528 12656
rect 176580 9353 176608 34054
rect 177212 30660 177264 30666
rect 177212 30602 177264 30608
rect 177224 26234 177252 30602
rect 177316 30530 177344 34054
rect 177396 30864 177448 30870
rect 177396 30806 177448 30812
rect 177304 30524 177356 30530
rect 177304 30466 177356 30472
rect 177224 26206 177344 26234
rect 176566 9344 176622 9353
rect 176566 9279 176622 9288
rect 176660 6180 176712 6186
rect 176660 6122 176712 6128
rect 174268 3324 174320 3330
rect 174268 3266 174320 3272
rect 175924 3324 175976 3330
rect 175924 3266 175976 3272
rect 173256 2848 173308 2854
rect 173256 2790 173308 2796
rect 174280 480 174308 3266
rect 175464 3120 175516 3126
rect 175464 3062 175516 3068
rect 175476 480 175504 3062
rect 176672 480 176700 6122
rect 177316 3262 177344 26206
rect 177304 3256 177356 3262
rect 177304 3198 177356 3204
rect 177408 3126 177436 30806
rect 177856 30524 177908 30530
rect 177856 30466 177908 30472
rect 177868 13938 177896 30466
rect 177856 13932 177908 13938
rect 177856 13874 177908 13880
rect 177960 12782 177988 34054
rect 178420 30530 178448 34054
rect 178972 30666 179000 34054
rect 178960 30660 179012 30666
rect 178960 30602 179012 30608
rect 178408 30524 178460 30530
rect 178408 30466 178460 30472
rect 179236 30524 179288 30530
rect 179236 30466 179288 30472
rect 177948 12776 178000 12782
rect 177948 12718 178000 12724
rect 179248 9217 179276 30466
rect 179234 9208 179290 9217
rect 179234 9143 179290 9152
rect 179340 6186 179368 34054
rect 179972 30932 180024 30938
rect 179972 30874 180024 30880
rect 179984 26234 180012 30874
rect 180076 30802 180104 34054
rect 180536 31074 180564 34054
rect 180524 31068 180576 31074
rect 180524 31010 180576 31016
rect 181180 30802 181208 34054
rect 180064 30796 180116 30802
rect 180064 30738 180116 30744
rect 180708 30796 180760 30802
rect 180708 30738 180760 30744
rect 181168 30796 181220 30802
rect 181168 30738 181220 30744
rect 179984 26206 180104 26234
rect 179328 6180 179380 6186
rect 179328 6122 179380 6128
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 177396 3120 177448 3126
rect 177396 3062 177448 3068
rect 177868 480 177896 3334
rect 180076 2990 180104 26206
rect 180720 9081 180748 30738
rect 181444 30592 181496 30598
rect 181444 30534 181496 30540
rect 181456 16574 181484 30534
rect 181732 26234 181760 34054
rect 181962 33810 181990 34068
rect 182528 34054 182864 34082
rect 183080 34054 183416 34082
rect 183632 34054 183968 34082
rect 184184 34054 184520 34082
rect 181962 33782 182036 33810
rect 181732 26206 181944 26234
rect 181456 16546 181576 16574
rect 180706 9072 180762 9081
rect 180706 9007 180762 9016
rect 181444 6044 181496 6050
rect 181444 5986 181496 5992
rect 180248 5976 180300 5982
rect 180248 5918 180300 5924
rect 179052 2984 179104 2990
rect 179052 2926 179104 2932
rect 180064 2984 180116 2990
rect 180064 2926 180116 2932
rect 179064 480 179092 2926
rect 180260 480 180288 5918
rect 181456 480 181484 5986
rect 181548 3126 181576 16546
rect 181916 14006 181944 26206
rect 182008 14074 182036 33782
rect 182088 30796 182140 30802
rect 182088 30738 182140 30744
rect 181996 14068 182048 14074
rect 181996 14010 182048 14016
rect 181904 14000 181956 14006
rect 181904 13942 181956 13948
rect 182100 5574 182128 30738
rect 182836 30598 182864 34054
rect 182824 30592 182876 30598
rect 182824 30534 182876 30540
rect 183388 14142 183416 34054
rect 183940 30802 183968 34054
rect 183928 30796 183980 30802
rect 183928 30738 183980 30744
rect 184492 30598 184520 34054
rect 184676 34054 184736 34082
rect 185288 34054 185624 34082
rect 185840 34054 186268 34082
rect 186392 34054 186728 34082
rect 187036 34054 187372 34082
rect 183468 30592 183520 30598
rect 183468 30534 183520 30540
rect 184480 30592 184532 30598
rect 184480 30534 184532 30540
rect 183376 14136 183428 14142
rect 183376 14078 183428 14084
rect 183480 5642 183508 30534
rect 184676 14210 184704 34054
rect 185492 31068 185544 31074
rect 185492 31010 185544 31016
rect 184848 30796 184900 30802
rect 184848 30738 184900 30744
rect 184756 30592 184808 30598
rect 184756 30534 184808 30540
rect 184664 14204 184716 14210
rect 184664 14146 184716 14152
rect 183744 6112 183796 6118
rect 183744 6054 183796 6060
rect 183468 5636 183520 5642
rect 183468 5578 183520 5584
rect 182088 5568 182140 5574
rect 182088 5510 182140 5516
rect 181536 3120 181588 3126
rect 181536 3062 181588 3068
rect 182548 3052 182600 3058
rect 182548 2994 182600 3000
rect 182560 480 182588 2994
rect 183756 480 183784 6054
rect 184768 5710 184796 30534
rect 184756 5704 184808 5710
rect 184756 5646 184808 5652
rect 184860 3058 184888 30738
rect 185504 26234 185532 31010
rect 185596 30870 185624 34054
rect 185584 30864 185636 30870
rect 185584 30806 185636 30812
rect 185504 26206 185624 26234
rect 185596 4146 185624 26206
rect 186240 5778 186268 34054
rect 186700 30598 186728 34054
rect 187344 30870 187372 34054
rect 187528 34054 187588 34082
rect 188140 34054 188476 34082
rect 188692 34054 189028 34082
rect 189244 34054 189580 34082
rect 189796 34054 190224 34082
rect 187332 30864 187384 30870
rect 187332 30806 187384 30812
rect 186688 30592 186740 30598
rect 186688 30534 186740 30540
rect 187424 30592 187476 30598
rect 187424 30534 187476 30540
rect 187436 14278 187464 30534
rect 187424 14272 187476 14278
rect 187424 14214 187476 14220
rect 187332 6792 187384 6798
rect 187332 6734 187384 6740
rect 186228 5772 186280 5778
rect 186228 5714 186280 5720
rect 184940 4140 184992 4146
rect 184940 4082 184992 4088
rect 185584 4140 185636 4146
rect 185584 4082 185636 4088
rect 184848 3052 184900 3058
rect 184848 2994 184900 3000
rect 184952 480 184980 4082
rect 186136 2916 186188 2922
rect 186136 2858 186188 2864
rect 186148 480 186176 2858
rect 187344 480 187372 6734
rect 187528 5846 187556 34054
rect 187608 30864 187660 30870
rect 187608 30806 187660 30812
rect 187516 5840 187568 5846
rect 187516 5782 187568 5788
rect 187620 3058 187648 30806
rect 188448 30598 188476 34054
rect 189000 31618 189028 34054
rect 188988 31612 189040 31618
rect 188988 31554 189040 31560
rect 189552 30870 189580 34054
rect 189540 30864 189592 30870
rect 189540 30806 189592 30812
rect 188436 30592 188488 30598
rect 188436 30534 188488 30540
rect 188988 30592 189040 30598
rect 188988 30534 189040 30540
rect 189000 9790 189028 30534
rect 190196 9858 190224 34054
rect 190334 33810 190362 34068
rect 190900 34054 191236 34082
rect 191452 34054 191696 34082
rect 192004 34054 192340 34082
rect 192556 34054 192892 34082
rect 190334 33782 190408 33810
rect 190276 30864 190328 30870
rect 190276 30806 190328 30812
rect 190184 9852 190236 9858
rect 190184 9794 190236 9800
rect 188988 9784 189040 9790
rect 188988 9726 189040 9732
rect 190288 5914 190316 30806
rect 190276 5908 190328 5914
rect 190276 5850 190328 5856
rect 188528 4072 188580 4078
rect 188528 4014 188580 4020
rect 187608 3052 187660 3058
rect 187608 2994 187660 3000
rect 188540 480 188568 4014
rect 190380 3194 190408 33782
rect 191208 30870 191236 34054
rect 191196 30864 191248 30870
rect 191196 30806 191248 30812
rect 191668 9926 191696 34054
rect 192312 30938 192340 34054
rect 192300 30932 192352 30938
rect 192300 30874 192352 30880
rect 191748 30864 191800 30870
rect 191748 30806 191800 30812
rect 191656 9920 191708 9926
rect 191656 9862 191708 9868
rect 190828 6724 190880 6730
rect 190828 6666 190880 6672
rect 189724 3188 189776 3194
rect 189724 3130 189776 3136
rect 190368 3188 190420 3194
rect 190368 3130 190420 3136
rect 189736 480 189764 3130
rect 190840 480 190868 6666
rect 191760 5982 191788 30806
rect 192864 30598 192892 34054
rect 193048 34054 193108 34082
rect 193660 34054 193996 34082
rect 194212 34054 194456 34082
rect 194764 34054 195100 34082
rect 195316 34054 195652 34082
rect 192852 30592 192904 30598
rect 192852 30534 192904 30540
rect 193048 9994 193076 34054
rect 193968 30870 193996 34054
rect 193956 30864 194008 30870
rect 193956 30806 194008 30812
rect 193128 30592 193180 30598
rect 193128 30534 193180 30540
rect 193036 9988 193088 9994
rect 193036 9930 193088 9936
rect 193140 6050 193168 30534
rect 194324 6656 194376 6662
rect 194324 6598 194376 6604
rect 193128 6044 193180 6050
rect 193128 5986 193180 5992
rect 191748 5976 191800 5982
rect 191748 5918 191800 5924
rect 192024 3936 192076 3942
rect 192024 3878 192076 3884
rect 192036 480 192064 3878
rect 194336 3346 194364 6598
rect 194428 6118 194456 34054
rect 194508 30864 194560 30870
rect 194508 30806 194560 30812
rect 194416 6112 194468 6118
rect 194416 6054 194468 6060
rect 194520 3942 194548 30806
rect 195072 30598 195100 34054
rect 195624 31006 195652 34054
rect 195854 33810 195882 34068
rect 196420 34054 196756 34082
rect 196972 34054 197308 34082
rect 197616 34054 197952 34082
rect 198168 34054 198596 34082
rect 195854 33782 195928 33810
rect 195612 31000 195664 31006
rect 195612 30942 195664 30948
rect 195060 30592 195112 30598
rect 195060 30534 195112 30540
rect 195796 30592 195848 30598
rect 195796 30534 195848 30540
rect 195808 10062 195836 30534
rect 195796 10056 195848 10062
rect 195796 9998 195848 10004
rect 195900 5273 195928 33782
rect 196728 30598 196756 34054
rect 196716 30592 196768 30598
rect 196716 30534 196768 30540
rect 197176 30592 197228 30598
rect 197176 30534 197228 30540
rect 197188 10130 197216 30534
rect 197176 10124 197228 10130
rect 197176 10066 197228 10072
rect 195886 5264 195942 5273
rect 195886 5199 195942 5208
rect 195612 4004 195664 4010
rect 195612 3946 195664 3952
rect 194508 3936 194560 3942
rect 194508 3878 194560 3884
rect 194336 3318 194456 3346
rect 193220 3256 193272 3262
rect 193220 3198 193272 3204
rect 193232 480 193260 3198
rect 194428 480 194456 3318
rect 195624 480 195652 3946
rect 197280 3330 197308 34054
rect 197924 30598 197952 34054
rect 197912 30592 197964 30598
rect 197912 30534 197964 30540
rect 198568 10198 198596 34054
rect 198660 34054 198720 34082
rect 199272 34054 199608 34082
rect 199824 34054 199976 34082
rect 200376 34054 200712 34082
rect 200928 34054 201356 34082
rect 198660 31210 198688 34054
rect 198648 31204 198700 31210
rect 198648 31146 198700 31152
rect 199580 30598 199608 34054
rect 198648 30592 198700 30598
rect 198648 30534 198700 30540
rect 199568 30592 199620 30598
rect 199568 30534 199620 30540
rect 198556 10192 198608 10198
rect 198556 10134 198608 10140
rect 198660 6798 198688 30534
rect 199948 10266 199976 34054
rect 200028 30592 200080 30598
rect 200028 30534 200080 30540
rect 199936 10260 199988 10266
rect 199936 10202 199988 10208
rect 198648 6792 198700 6798
rect 198648 6734 198700 6740
rect 200040 6730 200068 30534
rect 200684 30394 200712 34054
rect 200764 31748 200816 31754
rect 200764 31690 200816 31696
rect 200672 30388 200724 30394
rect 200672 30330 200724 30336
rect 200028 6724 200080 6730
rect 200028 6666 200080 6672
rect 197912 6588 197964 6594
rect 197912 6530 197964 6536
rect 197268 3324 197320 3330
rect 197268 3266 197320 3272
rect 196808 2916 196860 2922
rect 196808 2858 196860 2864
rect 196820 480 196848 2858
rect 197924 480 197952 6530
rect 200776 4282 200804 31690
rect 201224 30388 201276 30394
rect 201224 30330 201276 30336
rect 201236 11014 201264 30330
rect 201224 11008 201276 11014
rect 201224 10950 201276 10956
rect 201328 6662 201356 34054
rect 201420 34054 201480 34082
rect 202032 34054 202368 34082
rect 202584 34054 202828 34082
rect 203136 34054 203472 34082
rect 203688 34054 203932 34082
rect 201420 30394 201448 34054
rect 202340 31686 202368 34054
rect 202328 31680 202380 31686
rect 202328 31622 202380 31628
rect 201408 30388 201460 30394
rect 201408 30330 201460 30336
rect 201408 30252 201460 30258
rect 201408 30194 201460 30200
rect 201316 6656 201368 6662
rect 201316 6598 201368 6604
rect 200304 4276 200356 4282
rect 200304 4218 200356 4224
rect 200764 4276 200816 4282
rect 200764 4218 200816 4224
rect 199108 3868 199160 3874
rect 199108 3810 199160 3816
rect 199120 480 199148 3810
rect 200316 480 200344 4218
rect 201420 4146 201448 30194
rect 202800 12850 202828 34054
rect 203444 30598 203472 34054
rect 203432 30592 203484 30598
rect 203432 30534 203484 30540
rect 203904 30394 203932 34054
rect 203996 34054 204240 34082
rect 204792 34054 205128 34082
rect 205344 34054 205588 34082
rect 205896 34054 206232 34082
rect 206448 34054 206876 34082
rect 203892 30388 203944 30394
rect 203892 30330 203944 30336
rect 203996 12918 204024 34054
rect 204904 30932 204956 30938
rect 204904 30874 204956 30880
rect 204076 30592 204128 30598
rect 204076 30534 204128 30540
rect 203984 12912 204036 12918
rect 203984 12854 204036 12860
rect 202788 12844 202840 12850
rect 202788 12786 202840 12792
rect 204088 10946 204116 30534
rect 204168 30388 204220 30394
rect 204168 30330 204220 30336
rect 204076 10940 204128 10946
rect 204076 10882 204128 10888
rect 201500 8220 201552 8226
rect 201500 8162 201552 8168
rect 201408 4140 201460 4146
rect 201408 4082 201460 4088
rect 201512 480 201540 8162
rect 203892 4480 203944 4486
rect 203892 4422 203944 4428
rect 202696 3868 202748 3874
rect 202696 3810 202748 3816
rect 202708 480 202736 3810
rect 203904 480 203932 4422
rect 204180 4078 204208 30330
rect 204916 4486 204944 30874
rect 205100 30394 205128 34054
rect 205560 31278 205588 34054
rect 205548 31272 205600 31278
rect 205548 31214 205600 31220
rect 206204 30394 206232 34054
rect 205088 30388 205140 30394
rect 205088 30330 205140 30336
rect 205548 30388 205600 30394
rect 205548 30330 205600 30336
rect 206192 30388 206244 30394
rect 206192 30330 206244 30336
rect 206744 30388 206796 30394
rect 206744 30330 206796 30336
rect 205560 10878 205588 30330
rect 206756 14346 206784 30330
rect 206744 14340 206796 14346
rect 206744 14282 206796 14288
rect 205548 10872 205600 10878
rect 205548 10814 205600 10820
rect 206848 10810 206876 34054
rect 206940 34054 207000 34082
rect 207552 34054 208072 34082
rect 208196 34054 208348 34082
rect 208748 34054 209084 34082
rect 209300 34054 209728 34082
rect 209852 34054 210188 34082
rect 210404 34054 210740 34082
rect 206836 10804 206888 10810
rect 206836 10746 206888 10752
rect 205088 8152 205140 8158
rect 205088 8094 205140 8100
rect 204904 4480 204956 4486
rect 204904 4422 204956 4428
rect 204168 4072 204220 4078
rect 204168 4014 204220 4020
rect 205100 480 205128 8094
rect 206940 4010 206968 34054
rect 208044 26234 208072 34054
rect 208044 26206 208256 26234
rect 208228 14414 208256 26206
rect 208216 14408 208268 14414
rect 208216 14350 208268 14356
rect 208320 10742 208348 34054
rect 208952 31544 209004 31550
rect 208952 31486 209004 31492
rect 208964 26234 208992 31486
rect 209056 30938 209084 34054
rect 209044 30932 209096 30938
rect 209044 30874 209096 30880
rect 208964 26206 209084 26234
rect 208308 10736 208360 10742
rect 208308 10678 208360 10684
rect 208584 8084 208636 8090
rect 208584 8026 208636 8032
rect 207388 4412 207440 4418
rect 207388 4354 207440 4360
rect 206192 4004 206244 4010
rect 206192 3946 206244 3952
rect 206928 4004 206980 4010
rect 206928 3946 206980 3952
rect 206204 480 206232 3946
rect 207400 480 207428 4354
rect 208596 480 208624 8026
rect 209056 4418 209084 26206
rect 209700 7070 209728 34054
rect 210160 30394 210188 34054
rect 210712 30598 210740 34054
rect 210942 33810 210970 34068
rect 211508 34054 211844 34082
rect 212060 34054 212396 34082
rect 212612 34054 212948 34082
rect 213164 34054 213592 34082
rect 213716 34054 213868 34082
rect 214268 34054 214604 34082
rect 214820 34054 215156 34082
rect 215372 34054 215708 34082
rect 215924 34054 216260 34082
rect 210942 33782 211016 33810
rect 210700 30592 210752 30598
rect 210700 30534 210752 30540
rect 210148 30388 210200 30394
rect 210148 30330 210200 30336
rect 210884 30388 210936 30394
rect 210884 30330 210936 30336
rect 210896 10674 210924 30330
rect 210884 10668 210936 10674
rect 210884 10610 210936 10616
rect 210988 7138 211016 33782
rect 211068 30592 211120 30598
rect 211068 30534 211120 30540
rect 210976 7132 211028 7138
rect 210976 7074 211028 7080
rect 209688 7064 209740 7070
rect 209688 7006 209740 7012
rect 209044 4412 209096 4418
rect 209044 4354 209096 4360
rect 210976 4208 211028 4214
rect 210976 4150 211028 4156
rect 209780 3800 209832 3806
rect 209780 3742 209832 3748
rect 209792 480 209820 3742
rect 210988 480 211016 4150
rect 211080 3942 211108 30534
rect 211816 30394 211844 34054
rect 212368 31346 212396 34054
rect 212356 31340 212408 31346
rect 212356 31282 212408 31288
rect 212920 30394 212948 34054
rect 213184 31476 213236 31482
rect 213184 31418 213236 31424
rect 211804 30388 211856 30394
rect 211804 30330 211856 30336
rect 212448 30388 212500 30394
rect 212448 30330 212500 30336
rect 212908 30388 212960 30394
rect 212908 30330 212960 30336
rect 212460 10606 212488 30330
rect 212448 10600 212500 10606
rect 212448 10542 212500 10548
rect 213196 4214 213224 31418
rect 213564 26234 213592 34054
rect 213736 30388 213788 30394
rect 213736 30330 213788 30336
rect 213564 26206 213684 26234
rect 213656 10538 213684 26206
rect 213644 10532 213696 10538
rect 213644 10474 213696 10480
rect 213748 7206 213776 30330
rect 213736 7200 213788 7206
rect 213736 7142 213788 7148
rect 213184 4208 213236 4214
rect 213184 4150 213236 4156
rect 211068 3936 211120 3942
rect 211068 3878 211120 3884
rect 213840 3874 213868 34054
rect 214576 30394 214604 34054
rect 214564 30388 214616 30394
rect 214564 30330 214616 30336
rect 215128 10470 215156 34054
rect 215680 31754 215708 34054
rect 215668 31748 215720 31754
rect 215668 31690 215720 31696
rect 216232 30394 216260 34054
rect 216462 33810 216490 34068
rect 217028 34054 217364 34082
rect 217580 34054 217916 34082
rect 218132 34054 218468 34082
rect 218776 34054 219112 34082
rect 216462 33782 216536 33810
rect 215208 30388 215260 30394
rect 215208 30330 215260 30336
rect 216220 30388 216272 30394
rect 216220 30330 216272 30336
rect 215116 10464 215168 10470
rect 215116 10406 215168 10412
rect 215220 7274 215248 30330
rect 216508 10402 216536 33782
rect 217336 30394 217364 34054
rect 216588 30388 216640 30394
rect 216588 30330 216640 30336
rect 217324 30388 217376 30394
rect 217324 30330 217376 30336
rect 216496 10396 216548 10402
rect 216496 10338 216548 10344
rect 215668 7948 215720 7954
rect 215668 7890 215720 7896
rect 215208 7268 215260 7274
rect 215208 7210 215260 7216
rect 214472 4344 214524 4350
rect 214472 4286 214524 4292
rect 213828 3868 213880 3874
rect 213828 3810 213880 3816
rect 212172 3664 212224 3670
rect 212172 3606 212224 3612
rect 212184 480 212212 3606
rect 213368 3596 213420 3602
rect 213368 3538 213420 3544
rect 213380 480 213408 3538
rect 214484 480 214512 4286
rect 215680 480 215708 7890
rect 216600 7342 216628 30330
rect 217888 7410 217916 34054
rect 218440 30394 218468 34054
rect 219084 31482 219112 34054
rect 219314 33810 219342 34068
rect 219880 34054 220216 34082
rect 220432 34054 220768 34082
rect 220984 34054 221320 34082
rect 221536 34054 221964 34082
rect 219314 33782 219388 33810
rect 219072 31476 219124 31482
rect 219072 31418 219124 31424
rect 217968 30388 218020 30394
rect 217968 30330 218020 30336
rect 218428 30388 218480 30394
rect 218428 30330 218480 30336
rect 219256 30388 219308 30394
rect 219256 30330 219308 30336
rect 217876 7404 217928 7410
rect 217876 7346 217928 7352
rect 216588 7336 216640 7342
rect 216588 7278 216640 7284
rect 217980 3806 218008 30330
rect 219268 10334 219296 30330
rect 219256 10328 219308 10334
rect 219256 10270 219308 10276
rect 219256 8016 219308 8022
rect 219256 7958 219308 7964
rect 218060 4548 218112 4554
rect 218060 4490 218112 4496
rect 217968 3800 218020 3806
rect 216862 3768 216918 3777
rect 217968 3742 218020 3748
rect 216862 3703 216918 3712
rect 216876 480 216904 3703
rect 218072 480 218100 4490
rect 219268 480 219296 7958
rect 219360 7546 219388 33782
rect 220188 30394 220216 34054
rect 220176 30388 220228 30394
rect 220176 30330 220228 30336
rect 220636 30388 220688 30394
rect 220636 30330 220688 30336
rect 220648 10713 220676 30330
rect 220634 10704 220690 10713
rect 220634 10639 220690 10648
rect 219348 7540 219400 7546
rect 219348 7482 219400 7488
rect 220740 3738 220768 34054
rect 221292 30394 221320 34054
rect 221280 30388 221332 30394
rect 221280 30330 221332 30336
rect 221936 26234 221964 34054
rect 222028 34054 222088 34082
rect 222640 34054 222976 34082
rect 223192 34054 223436 34082
rect 223744 34054 224080 34082
rect 224296 34054 224632 34082
rect 222028 31142 222056 34054
rect 222016 31136 222068 31142
rect 222016 31078 222068 31084
rect 222948 30394 222976 34054
rect 222108 30388 222160 30394
rect 222108 30330 222160 30336
rect 222936 30388 222988 30394
rect 222936 30330 222988 30336
rect 221936 26206 222056 26234
rect 222028 10577 222056 26206
rect 222014 10568 222070 10577
rect 222014 10503 222070 10512
rect 222120 7478 222148 30330
rect 223408 10441 223436 34054
rect 224052 30598 224080 34054
rect 224040 30592 224092 30598
rect 224040 30534 224092 30540
rect 224604 30394 224632 34054
rect 224696 34054 224848 34082
rect 225400 34054 225736 34082
rect 225952 34054 226288 34082
rect 226504 34054 226840 34082
rect 227056 34054 227392 34082
rect 223488 30388 223540 30394
rect 223488 30330 223540 30336
rect 224592 30388 224644 30394
rect 224592 30330 224644 30336
rect 223394 10432 223450 10441
rect 223394 10367 223450 10376
rect 223500 8294 223528 30330
rect 224696 10305 224724 34054
rect 225708 31414 225736 34054
rect 225696 31408 225748 31414
rect 225696 31350 225748 31356
rect 224868 30592 224920 30598
rect 224868 30534 224920 30540
rect 224776 30388 224828 30394
rect 224776 30330 224828 30336
rect 224682 10296 224738 10305
rect 224682 10231 224738 10240
rect 223488 8288 223540 8294
rect 223488 8230 223540 8236
rect 224788 8226 224816 30330
rect 224776 8220 224828 8226
rect 224776 8162 224828 8168
rect 222752 7880 222804 7886
rect 222752 7822 222804 7828
rect 222108 7472 222160 7478
rect 222108 7414 222160 7420
rect 221556 4616 221608 4622
rect 221556 4558 221608 4564
rect 220728 3732 220780 3738
rect 220728 3674 220780 3680
rect 220452 3528 220504 3534
rect 220452 3470 220504 3476
rect 220464 480 220492 3470
rect 221568 480 221596 4558
rect 222764 480 222792 7822
rect 224880 3670 224908 30534
rect 226260 8158 226288 34054
rect 226812 30394 226840 34054
rect 227364 30598 227392 34054
rect 227548 34054 227608 34082
rect 228160 34054 228496 34082
rect 228712 34054 228956 34082
rect 229356 34054 229692 34082
rect 229908 34054 230244 34082
rect 227352 30592 227404 30598
rect 227352 30534 227404 30540
rect 226800 30388 226852 30394
rect 226800 30330 226852 30336
rect 227444 30388 227496 30394
rect 227444 30330 227496 30336
rect 227456 15162 227484 30330
rect 227444 15156 227496 15162
rect 227444 15098 227496 15104
rect 226248 8152 226300 8158
rect 226248 8094 226300 8100
rect 227548 8022 227576 34054
rect 227628 30592 227680 30598
rect 227628 30534 227680 30540
rect 227536 8016 227588 8022
rect 227536 7958 227588 7964
rect 226340 7812 226392 7818
rect 226340 7754 226392 7760
rect 225144 4684 225196 4690
rect 225144 4626 225196 4632
rect 224868 3664 224920 3670
rect 223946 3632 224002 3641
rect 224868 3606 224920 3612
rect 223946 3567 224002 3576
rect 223960 480 223988 3567
rect 225156 480 225184 4626
rect 226352 480 226380 7754
rect 227640 3602 227668 30534
rect 228468 30394 228496 34054
rect 228928 31074 228956 34054
rect 228916 31068 228968 31074
rect 228916 31010 228968 31016
rect 229664 30394 229692 34054
rect 228456 30388 228508 30394
rect 228456 30330 228508 30336
rect 229008 30388 229060 30394
rect 229008 30330 229060 30336
rect 229652 30388 229704 30394
rect 229652 30330 229704 30336
rect 229020 15094 229048 30330
rect 229008 15088 229060 15094
rect 229008 15030 229060 15036
rect 230216 15026 230244 34054
rect 230400 34054 230460 34082
rect 231012 34054 231348 34082
rect 231564 34054 231716 34082
rect 232116 34054 232452 34082
rect 232668 34054 233004 34082
rect 230296 30388 230348 30394
rect 230296 30330 230348 30336
rect 230204 15020 230256 15026
rect 230204 14962 230256 14968
rect 230308 8090 230336 30330
rect 230296 8084 230348 8090
rect 230296 8026 230348 8032
rect 228732 4752 228784 4758
rect 228732 4694 228784 4700
rect 227628 3596 227680 3602
rect 227628 3538 227680 3544
rect 227534 3496 227590 3505
rect 227534 3431 227590 3440
rect 227548 480 227576 3431
rect 228744 480 228772 4694
rect 230400 3534 230428 34054
rect 231320 30394 231348 34054
rect 231308 30388 231360 30394
rect 231308 30330 231360 30336
rect 231688 14958 231716 34054
rect 232424 30598 232452 34054
rect 232412 30592 232464 30598
rect 232412 30534 232464 30540
rect 232976 30394 233004 34054
rect 233068 34054 233220 34082
rect 233772 34054 234200 34082
rect 234324 34054 234568 34082
rect 234876 34054 235212 34082
rect 235428 34054 235764 34082
rect 231768 30388 231820 30394
rect 231768 30330 231820 30336
rect 232964 30388 233016 30394
rect 232964 30330 233016 30336
rect 231676 14952 231728 14958
rect 231676 14894 231728 14900
rect 231780 7954 231808 30330
rect 233068 14890 233096 34054
rect 233148 30388 233200 30394
rect 233148 30330 233200 30336
rect 233056 14884 233108 14890
rect 233056 14826 233108 14832
rect 231768 7948 231820 7954
rect 231768 7890 231820 7896
rect 233160 7886 233188 30330
rect 234172 26234 234200 34054
rect 234172 26206 234476 26234
rect 234448 16114 234476 26206
rect 234436 16108 234488 16114
rect 234436 16050 234488 16056
rect 233148 7880 233200 7886
rect 233148 7822 233200 7828
rect 234540 7818 234568 34054
rect 235184 30394 235212 34054
rect 235172 30388 235224 30394
rect 235172 30330 235224 30336
rect 235736 30326 235764 34054
rect 235920 34054 235980 34082
rect 236532 34054 236960 34082
rect 237084 34054 237328 34082
rect 237636 34054 237972 34082
rect 238188 34054 238616 34082
rect 235816 30388 235868 30394
rect 235816 30330 235868 30336
rect 235724 30320 235776 30326
rect 235724 30262 235776 30268
rect 235828 11218 235856 30330
rect 235816 11212 235868 11218
rect 235816 11154 235868 11160
rect 234528 7812 234580 7818
rect 234528 7754 234580 7760
rect 235920 7750 235948 34054
rect 236932 26234 236960 34054
rect 236932 26206 237236 26234
rect 234620 7744 234672 7750
rect 234620 7686 234672 7692
rect 235908 7744 235960 7750
rect 235908 7686 235960 7692
rect 232228 5500 232280 5506
rect 232228 5442 232280 5448
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 231032 3460 231084 3466
rect 231032 3402 231084 3408
rect 229836 2848 229888 2854
rect 229836 2790 229888 2796
rect 229848 480 229876 2790
rect 231044 480 231072 3402
rect 232240 480 232268 5442
rect 233424 2984 233476 2990
rect 233424 2926 233476 2932
rect 233436 480 233464 2926
rect 234632 480 234660 7686
rect 237208 6594 237236 26206
rect 237196 6588 237248 6594
rect 237196 6530 237248 6536
rect 235814 5128 235870 5137
rect 235814 5063 235870 5072
rect 235828 480 235856 5063
rect 237300 3466 237328 34054
rect 237944 31482 237972 34054
rect 237932 31476 237984 31482
rect 237932 31418 237984 31424
rect 238588 11286 238616 34054
rect 238680 34054 238740 34082
rect 239292 34054 239628 34082
rect 238680 31634 238708 34054
rect 238680 31606 238800 31634
rect 238668 31476 238720 31482
rect 238668 31418 238720 31424
rect 238576 11280 238628 11286
rect 238576 11222 238628 11228
rect 238680 7993 238708 31418
rect 238772 30977 238800 31606
rect 238758 30968 238814 30977
rect 238758 30903 238814 30912
rect 239600 30394 239628 34054
rect 239922 33810 239950 34068
rect 240488 34054 240824 34082
rect 241040 34054 241468 34082
rect 241592 34054 241928 34082
rect 242144 34054 242480 34082
rect 242696 34054 242848 34082
rect 243248 34054 243584 34082
rect 243800 34054 244136 34082
rect 244352 34054 244688 34082
rect 244904 34054 245332 34082
rect 239922 33782 239996 33810
rect 239588 30388 239640 30394
rect 239588 30330 239640 30336
rect 239968 11354 239996 33782
rect 240796 30394 240824 34054
rect 240048 30388 240100 30394
rect 240048 30330 240100 30336
rect 240784 30388 240836 30394
rect 240784 30330 240836 30336
rect 241336 30388 241388 30394
rect 241336 30330 241388 30336
rect 239956 11348 240008 11354
rect 239956 11290 240008 11296
rect 238666 7984 238722 7993
rect 238666 7919 238722 7928
rect 240060 7857 240088 30330
rect 241348 16046 241376 30330
rect 241336 16040 241388 16046
rect 241336 15982 241388 15988
rect 240046 7848 240102 7857
rect 240046 7783 240102 7792
rect 241440 7721 241468 34054
rect 241900 30394 241928 34054
rect 242452 30462 242480 34054
rect 242164 30456 242216 30462
rect 242164 30398 242216 30404
rect 242440 30456 242492 30462
rect 242440 30398 242492 30404
rect 241888 30388 241940 30394
rect 241888 30330 241940 30336
rect 241426 7712 241482 7721
rect 241426 7647 241482 7656
rect 241704 7676 241756 7682
rect 241704 7618 241756 7624
rect 240508 6860 240560 6866
rect 240508 6802 240560 6808
rect 239312 5432 239364 5438
rect 239312 5374 239364 5380
rect 237288 3460 237340 3466
rect 237288 3402 237340 3408
rect 238114 3360 238170 3369
rect 238114 3295 238170 3304
rect 237012 3120 237064 3126
rect 237012 3062 237064 3068
rect 237024 480 237052 3062
rect 238128 480 238156 3295
rect 239324 480 239352 5374
rect 240520 480 240548 6802
rect 241716 480 241744 7618
rect 242176 6866 242204 30398
rect 242716 30388 242768 30394
rect 242716 30330 242768 30336
rect 242728 11422 242756 30330
rect 242716 11416 242768 11422
rect 242716 11358 242768 11364
rect 242820 7682 242848 34054
rect 243556 30394 243584 34054
rect 243544 30388 243596 30394
rect 243544 30330 243596 30336
rect 244108 15978 244136 34054
rect 244660 30394 244688 34054
rect 244924 30524 244976 30530
rect 244924 30466 244976 30472
rect 244188 30388 244240 30394
rect 244188 30330 244240 30336
rect 244648 30388 244700 30394
rect 244648 30330 244700 30336
rect 244096 15972 244148 15978
rect 244096 15914 244148 15920
rect 244200 11490 244228 30330
rect 244188 11484 244240 11490
rect 244188 11426 244240 11432
rect 244936 9722 244964 30466
rect 245304 26234 245332 34054
rect 245442 33810 245470 34068
rect 246008 34054 246344 34082
rect 246560 34054 246896 34082
rect 247112 34054 247448 34082
rect 247664 34054 248092 34082
rect 248216 34054 248368 34082
rect 248768 34054 249104 34082
rect 249320 34054 249748 34082
rect 249872 34054 250208 34082
rect 250516 34054 250852 34082
rect 245442 33782 245516 33810
rect 245488 30462 245516 33782
rect 245476 30456 245528 30462
rect 245476 30398 245528 30404
rect 246316 30394 246344 34054
rect 245568 30388 245620 30394
rect 245568 30330 245620 30336
rect 246304 30388 246356 30394
rect 246304 30330 246356 30336
rect 245304 26206 245516 26234
rect 245488 11558 245516 26206
rect 245476 11552 245528 11558
rect 245476 11494 245528 11500
rect 244924 9716 244976 9722
rect 244924 9658 244976 9664
rect 242808 7676 242860 7682
rect 242808 7618 242860 7624
rect 245580 7614 245608 30330
rect 246868 11626 246896 34054
rect 247420 30394 247448 34054
rect 248064 30546 248092 34054
rect 248064 30518 248276 30546
rect 246948 30388 247000 30394
rect 246948 30330 247000 30336
rect 247408 30388 247460 30394
rect 247408 30330 247460 30336
rect 248144 30388 248196 30394
rect 248144 30330 248196 30336
rect 246856 11620 246908 11626
rect 246856 11562 246908 11568
rect 245200 7608 245252 7614
rect 245200 7550 245252 7556
rect 245568 7608 245620 7614
rect 246960 7585 246988 30330
rect 248156 15910 248184 30330
rect 248144 15904 248196 15910
rect 248144 15846 248196 15852
rect 248248 14822 248276 30518
rect 248236 14816 248288 14822
rect 248236 14758 248288 14764
rect 248340 11694 248368 34054
rect 249076 31249 249104 34054
rect 249062 31240 249118 31249
rect 249062 31175 249118 31184
rect 249720 14754 249748 34054
rect 250180 30530 250208 34054
rect 250824 31822 250852 34054
rect 251008 34054 251068 34082
rect 251620 34054 251956 34082
rect 252172 34054 252508 34082
rect 252724 34054 253060 34082
rect 253276 34054 253704 34082
rect 250812 31816 250864 31822
rect 250812 31758 250864 31764
rect 251008 30818 251036 34054
rect 251088 31816 251140 31822
rect 251088 31758 251140 31764
rect 250916 30790 251036 30818
rect 250168 30524 250220 30530
rect 250168 30466 250220 30472
rect 249708 14748 249760 14754
rect 249708 14690 249760 14696
rect 250916 14618 250944 30790
rect 250996 30524 251048 30530
rect 250996 30466 251048 30472
rect 250904 14612 250956 14618
rect 250904 14554 250956 14560
rect 251008 12442 251036 30466
rect 250996 12436 251048 12442
rect 250996 12378 251048 12384
rect 248328 11688 248380 11694
rect 248328 11630 248380 11636
rect 248788 8492 248840 8498
rect 248788 8434 248840 8440
rect 245568 7550 245620 7556
rect 246946 7576 247002 7585
rect 242164 6860 242216 6866
rect 242164 6802 242216 6808
rect 244096 6520 244148 6526
rect 244096 6462 244148 6468
rect 242900 5364 242952 5370
rect 242900 5306 242952 5312
rect 242912 480 242940 5306
rect 244108 480 244136 6462
rect 245212 480 245240 7550
rect 246946 7511 247002 7520
rect 247592 6452 247644 6458
rect 247592 6394 247644 6400
rect 246396 5296 246448 5302
rect 246396 5238 246448 5244
rect 246408 480 246436 5238
rect 247604 480 247632 6394
rect 248800 480 248828 8434
rect 249984 5228 250036 5234
rect 249984 5170 250036 5176
rect 249996 480 250024 5170
rect 251100 3505 251128 31758
rect 251928 30530 251956 34054
rect 252480 31113 252508 34054
rect 252466 31104 252522 31113
rect 252466 31039 252522 31048
rect 253032 30530 253060 34054
rect 251916 30524 251968 30530
rect 251916 30466 251968 30472
rect 252468 30524 252520 30530
rect 252468 30466 252520 30472
rect 253020 30524 253072 30530
rect 253020 30466 253072 30472
rect 253572 30524 253624 30530
rect 253572 30466 253624 30472
rect 252480 12374 252508 30466
rect 253584 26234 253612 30466
rect 253676 30138 253704 34054
rect 253814 33810 253842 34068
rect 254380 34054 254716 34082
rect 254932 34054 255268 34082
rect 255484 34054 255820 34082
rect 256036 34054 256464 34082
rect 253814 33782 253888 33810
rect 253676 30110 253796 30138
rect 253584 26206 253704 26234
rect 253676 14686 253704 26206
rect 253664 14680 253716 14686
rect 253664 14622 253716 14628
rect 252468 12368 252520 12374
rect 252468 12310 252520 12316
rect 253768 12306 253796 30110
rect 253756 12300 253808 12306
rect 253756 12242 253808 12248
rect 252376 8560 252428 8566
rect 252376 8502 252428 8508
rect 251180 6384 251232 6390
rect 251180 6326 251232 6332
rect 251086 3496 251142 3505
rect 251086 3431 251142 3440
rect 251192 480 251220 6326
rect 252388 480 252416 8502
rect 253480 5160 253532 5166
rect 253480 5102 253532 5108
rect 253492 480 253520 5102
rect 253860 3369 253888 33782
rect 254688 30530 254716 34054
rect 254676 30524 254728 30530
rect 254676 30466 254728 30472
rect 255136 30524 255188 30530
rect 255136 30466 255188 30472
rect 255148 12986 255176 30466
rect 255136 12980 255188 12986
rect 255136 12922 255188 12928
rect 255240 8498 255268 34054
rect 255792 30530 255820 34054
rect 255780 30524 255832 30530
rect 255780 30466 255832 30472
rect 256436 13054 256464 34054
rect 256574 33810 256602 34068
rect 257140 34054 257476 34082
rect 257692 34054 257936 34082
rect 258244 34054 258580 34082
rect 258796 34054 259132 34082
rect 256574 33782 256648 33810
rect 256516 30524 256568 30530
rect 256516 30466 256568 30472
rect 256424 13048 256476 13054
rect 256424 12990 256476 12996
rect 256528 12238 256556 30466
rect 256516 12232 256568 12238
rect 256516 12174 256568 12180
rect 255872 8628 255924 8634
rect 255872 8570 255924 8576
rect 255228 8492 255280 8498
rect 255228 8434 255280 8440
rect 254674 6624 254730 6633
rect 254674 6559 254730 6568
rect 253846 3360 253902 3369
rect 253846 3295 253902 3304
rect 254688 480 254716 6559
rect 255884 480 255912 8570
rect 256620 8566 256648 33782
rect 257448 30530 257476 34054
rect 257436 30524 257488 30530
rect 257436 30466 257488 30472
rect 257908 13802 257936 34054
rect 257988 30524 258040 30530
rect 257988 30466 258040 30472
rect 257896 13796 257948 13802
rect 257896 13738 257948 13744
rect 258000 12170 258028 30466
rect 258552 27334 258580 34054
rect 259104 30530 259132 34054
rect 259196 34054 259348 34082
rect 259900 34054 260236 34082
rect 260452 34054 260696 34082
rect 261096 34054 261432 34082
rect 261648 34054 261984 34082
rect 259092 30524 259144 30530
rect 259092 30466 259144 30472
rect 258540 27328 258592 27334
rect 258540 27270 258592 27276
rect 259196 13734 259224 34054
rect 260208 30530 260236 34054
rect 259276 30524 259328 30530
rect 259276 30466 259328 30472
rect 260196 30524 260248 30530
rect 260196 30466 260248 30472
rect 259184 13728 259236 13734
rect 259184 13670 259236 13676
rect 257988 12164 258040 12170
rect 257988 12106 258040 12112
rect 259288 12102 259316 30466
rect 259368 27328 259420 27334
rect 259368 27270 259420 27276
rect 259276 12096 259328 12102
rect 259276 12038 259328 12044
rect 259380 8634 259408 27270
rect 260668 12034 260696 34054
rect 261404 30530 261432 34054
rect 261956 31822 261984 34054
rect 262048 34054 262200 34082
rect 262752 34054 263088 34082
rect 263304 34054 263456 34082
rect 263856 34054 264192 34082
rect 264408 34054 264744 34082
rect 261944 31816 261996 31822
rect 261944 31758 261996 31764
rect 260748 30524 260800 30530
rect 260748 30466 260800 30472
rect 261392 30524 261444 30530
rect 261392 30466 261444 30472
rect 261944 30524 261996 30530
rect 261944 30466 261996 30472
rect 260656 12028 260708 12034
rect 260656 11970 260708 11976
rect 259460 8696 259512 8702
rect 259460 8638 259512 8644
rect 259368 8628 259420 8634
rect 259368 8570 259420 8576
rect 256608 8560 256660 8566
rect 256608 8502 256660 8508
rect 258262 6488 258318 6497
rect 258262 6423 258318 6432
rect 257068 5092 257120 5098
rect 257068 5034 257120 5040
rect 257080 480 257108 5034
rect 258276 480 258304 6423
rect 259472 480 259500 8638
rect 260760 6526 260788 30466
rect 261956 13666 261984 30466
rect 261944 13660 261996 13666
rect 261944 13602 261996 13608
rect 262048 11966 262076 34054
rect 262128 31816 262180 31822
rect 262128 31758 262180 31764
rect 262036 11960 262088 11966
rect 262036 11902 262088 11908
rect 262140 8702 262168 31758
rect 263060 30530 263088 34054
rect 263048 30524 263100 30530
rect 263048 30466 263100 30472
rect 263428 8770 263456 34054
rect 264164 30530 264192 34054
rect 264716 31822 264744 34054
rect 264808 34054 264960 34082
rect 265512 34054 265940 34082
rect 266064 34054 266308 34082
rect 266616 34054 266952 34082
rect 267168 34054 267504 34082
rect 264704 31816 264756 31822
rect 264704 31758 264756 31764
rect 263508 30524 263560 30530
rect 263508 30466 263560 30472
rect 264152 30524 264204 30530
rect 264152 30466 264204 30472
rect 264704 30524 264756 30530
rect 264704 30466 264756 30472
rect 262956 8764 263008 8770
rect 262956 8706 263008 8712
rect 263416 8764 263468 8770
rect 263416 8706 263468 8712
rect 262128 8696 262180 8702
rect 262128 8638 262180 8644
rect 260748 6520 260800 6526
rect 260748 6462 260800 6468
rect 261760 6316 261812 6322
rect 261760 6258 261812 6264
rect 260654 4992 260710 5001
rect 260654 4927 260710 4936
rect 260668 480 260696 4927
rect 261772 480 261800 6258
rect 262968 480 262996 8706
rect 263520 4690 263548 30466
rect 264716 11898 264744 30466
rect 264704 11892 264756 11898
rect 264704 11834 264756 11840
rect 264808 6458 264836 34054
rect 264888 31816 264940 31822
rect 264888 31758 264940 31764
rect 264796 6452 264848 6458
rect 264796 6394 264848 6400
rect 264152 5024 264204 5030
rect 264152 4966 264204 4972
rect 263508 4684 263560 4690
rect 263508 4626 263560 4632
rect 264164 480 264192 4966
rect 264900 4622 264928 31758
rect 265912 26234 265940 34054
rect 265912 26206 266216 26234
rect 266188 11830 266216 26206
rect 266176 11824 266228 11830
rect 266176 11766 266228 11772
rect 265346 6352 265402 6361
rect 265346 6287 265402 6296
rect 264888 4616 264940 4622
rect 264888 4558 264940 4564
rect 265360 480 265388 6287
rect 266280 4214 266308 34054
rect 266924 30530 266952 34054
rect 266912 30524 266964 30530
rect 266912 30466 266964 30472
rect 267476 11762 267504 34054
rect 267660 34054 267720 34082
rect 268272 34054 268608 34082
rect 268824 34054 268976 34082
rect 269376 34054 269712 34082
rect 269928 34054 270356 34082
rect 267556 30524 267608 30530
rect 267556 30466 267608 30472
rect 267464 11756 267516 11762
rect 267464 11698 267516 11704
rect 267568 8838 267596 30466
rect 266544 8832 266596 8838
rect 266544 8774 266596 8780
rect 267556 8832 267608 8838
rect 267556 8774 267608 8780
rect 266268 4208 266320 4214
rect 266268 4150 266320 4156
rect 266556 480 266584 8774
rect 267660 4350 267688 34054
rect 268580 30530 268608 34054
rect 268568 30524 268620 30530
rect 268568 30466 268620 30472
rect 268948 12073 268976 34054
rect 269684 30666 269712 34054
rect 269672 30660 269724 30666
rect 269672 30602 269724 30608
rect 269028 30524 269080 30530
rect 269028 30466 269080 30472
rect 270224 30524 270276 30530
rect 270224 30466 270276 30472
rect 268934 12064 268990 12073
rect 268934 11999 268990 12008
rect 269040 6390 269068 30466
rect 270236 11801 270264 30466
rect 270222 11792 270278 11801
rect 270222 11727 270278 11736
rect 270328 8906 270356 34054
rect 270420 34054 270480 34082
rect 271032 34054 271368 34082
rect 270420 30530 270448 34054
rect 270500 30660 270552 30666
rect 270500 30602 270552 30608
rect 270408 30524 270460 30530
rect 270408 30466 270460 30472
rect 270512 30410 270540 30602
rect 271340 30530 271368 34054
rect 271662 33810 271690 34068
rect 272228 34054 272564 34082
rect 272780 34054 273208 34082
rect 273332 34054 273668 34082
rect 273884 34054 274312 34082
rect 274436 34054 274588 34082
rect 274988 34054 275324 34082
rect 275540 34054 275876 34082
rect 276092 34054 276428 34082
rect 276644 34054 276980 34082
rect 271662 33782 271736 33810
rect 271328 30524 271380 30530
rect 271328 30466 271380 30472
rect 270420 30382 270540 30410
rect 270040 8900 270092 8906
rect 270040 8842 270092 8848
rect 270316 8900 270368 8906
rect 270316 8842 270368 8848
rect 269028 6384 269080 6390
rect 269028 6326 269080 6332
rect 268844 6248 268896 6254
rect 268844 6190 268896 6196
rect 267738 4856 267794 4865
rect 267738 4791 267794 4800
rect 267648 4344 267700 4350
rect 267648 4286 267700 4292
rect 267752 480 267780 4791
rect 268856 480 268884 6190
rect 270052 480 270080 8842
rect 270420 5030 270448 30382
rect 271708 6322 271736 33782
rect 272536 30530 272564 34054
rect 271788 30524 271840 30530
rect 271788 30466 271840 30472
rect 272524 30524 272576 30530
rect 272524 30466 272576 30472
rect 273076 30524 273128 30530
rect 273076 30466 273128 30472
rect 271696 6316 271748 6322
rect 271696 6258 271748 6264
rect 271800 5098 271828 30466
rect 273088 11937 273116 30466
rect 273074 11928 273130 11937
rect 273074 11863 273130 11872
rect 272430 6216 272486 6225
rect 272430 6151 272486 6160
rect 271788 5092 271840 5098
rect 271788 5034 271840 5040
rect 270408 5024 270460 5030
rect 270408 4966 270460 4972
rect 271236 4956 271288 4962
rect 271236 4898 271288 4904
rect 271248 480 271276 4898
rect 272444 480 272472 6151
rect 273180 5166 273208 34054
rect 273640 30530 273668 34054
rect 273628 30524 273680 30530
rect 273628 30466 273680 30472
rect 274284 26234 274312 34054
rect 274456 30524 274508 30530
rect 274456 30466 274508 30472
rect 274284 26206 274404 26234
rect 274376 11665 274404 26206
rect 274362 11656 274418 11665
rect 274362 11591 274418 11600
rect 274468 9654 274496 30466
rect 273628 9648 273680 9654
rect 273628 9590 273680 9596
rect 274456 9648 274508 9654
rect 274456 9590 274508 9596
rect 273168 5160 273220 5166
rect 273168 5102 273220 5108
rect 273640 480 273668 9590
rect 274560 5030 274588 34054
rect 275296 30530 275324 34054
rect 275284 30524 275336 30530
rect 275284 30466 275336 30472
rect 275848 13598 275876 34054
rect 276400 30666 276428 34054
rect 276296 30660 276348 30666
rect 276296 30602 276348 30608
rect 276388 30660 276440 30666
rect 276388 30602 276440 30608
rect 275928 30524 275980 30530
rect 275928 30466 275980 30472
rect 275836 13592 275888 13598
rect 275836 13534 275888 13540
rect 274824 13456 274876 13462
rect 274824 13398 274876 13404
rect 274548 5024 274600 5030
rect 274548 4966 274600 4972
rect 274836 480 274864 13398
rect 275940 6254 275968 30466
rect 276308 26234 276336 30602
rect 276952 30530 276980 34054
rect 277136 34054 277196 34082
rect 277748 34054 278084 34082
rect 278300 34054 278636 34082
rect 278852 34054 279188 34082
rect 279404 34054 279740 34082
rect 276940 30524 276992 30530
rect 276940 30466 276992 30472
rect 276308 26206 276704 26234
rect 276676 7002 276704 26206
rect 277136 13462 277164 34054
rect 277308 30660 277360 30666
rect 277308 30602 277360 30608
rect 277216 30524 277268 30530
rect 277216 30466 277268 30472
rect 277124 13456 277176 13462
rect 277124 13398 277176 13404
rect 277228 9586 277256 30466
rect 277124 9580 277176 9586
rect 277124 9522 277176 9528
rect 277216 9580 277268 9586
rect 277216 9522 277268 9528
rect 276020 6996 276072 7002
rect 276020 6938 276072 6944
rect 276664 6996 276716 7002
rect 276664 6938 276716 6944
rect 275928 6248 275980 6254
rect 275928 6190 275980 6196
rect 276032 480 276060 6938
rect 277136 480 277164 9522
rect 277320 4962 277348 30602
rect 278056 30530 278084 34054
rect 278044 30524 278096 30530
rect 278044 30466 278096 30472
rect 278320 13388 278372 13394
rect 278320 13330 278372 13336
rect 277308 4956 277360 4962
rect 277308 4898 277360 4904
rect 278332 480 278360 13330
rect 278608 6633 278636 34054
rect 279160 30530 279188 34054
rect 279712 30666 279740 34054
rect 279942 33810 279970 34068
rect 280508 34054 280844 34082
rect 281060 34054 281488 34082
rect 281612 34054 281948 34082
rect 282256 34054 282684 34082
rect 279942 33782 280016 33810
rect 279700 30660 279752 30666
rect 279700 30602 279752 30608
rect 278688 30524 278740 30530
rect 278688 30466 278740 30472
rect 279148 30524 279200 30530
rect 279148 30466 279200 30472
rect 279884 30524 279936 30530
rect 279884 30466 279936 30472
rect 278594 6624 278650 6633
rect 278594 6559 278650 6568
rect 278700 5506 278728 30466
rect 279896 13530 279924 30466
rect 279884 13524 279936 13530
rect 279884 13466 279936 13472
rect 279988 9518 280016 33782
rect 280068 30660 280120 30666
rect 280068 30602 280120 30608
rect 279516 9512 279568 9518
rect 279516 9454 279568 9460
rect 279976 9512 280028 9518
rect 279976 9454 280028 9460
rect 278688 5500 278740 5506
rect 278688 5442 278740 5448
rect 279528 480 279556 9454
rect 280080 5438 280108 30602
rect 280816 30530 280844 34054
rect 280804 30524 280856 30530
rect 280804 30466 280856 30472
rect 281356 30524 281408 30530
rect 281356 30466 281408 30472
rect 281368 13394 281396 30466
rect 281356 13388 281408 13394
rect 281356 13330 281408 13336
rect 280712 9444 280764 9450
rect 280712 9386 280764 9392
rect 280068 5432 280120 5438
rect 280068 5374 280120 5380
rect 280724 480 280752 9386
rect 281460 5370 281488 34054
rect 281920 30530 281948 34054
rect 281908 30524 281960 30530
rect 281908 30466 281960 30472
rect 282656 13433 282684 34054
rect 282794 33810 282822 34068
rect 283360 34054 283696 34082
rect 283912 34054 284156 34082
rect 284464 34054 284800 34082
rect 285016 34054 285352 34082
rect 282794 33782 282868 33810
rect 282736 30524 282788 30530
rect 282736 30466 282788 30472
rect 282642 13424 282698 13433
rect 282642 13359 282698 13368
rect 282748 9518 282776 30466
rect 282736 9512 282788 9518
rect 282736 9454 282788 9460
rect 281448 5364 281500 5370
rect 281448 5306 281500 5312
rect 282840 5302 282868 33782
rect 283668 30530 283696 34054
rect 283656 30524 283708 30530
rect 283656 30466 283708 30472
rect 284128 13297 284156 34054
rect 284772 30666 284800 34054
rect 284760 30660 284812 30666
rect 284760 30602 284812 30608
rect 285324 30530 285352 34054
rect 285416 34054 285568 34082
rect 286120 34054 286456 34082
rect 286672 34054 286916 34082
rect 287224 34054 287560 34082
rect 287776 34054 288112 34082
rect 284208 30524 284260 30530
rect 284208 30466 284260 30472
rect 285312 30524 285364 30530
rect 285312 30466 285364 30472
rect 284114 13288 284170 13297
rect 284114 13223 284170 13232
rect 284220 9450 284248 30466
rect 285416 13326 285444 34054
rect 285588 30660 285640 30666
rect 285588 30602 285640 30608
rect 285496 30524 285548 30530
rect 285496 30466 285548 30472
rect 284944 13320 284996 13326
rect 284944 13262 284996 13268
rect 285404 13320 285456 13326
rect 285404 13262 285456 13268
rect 284208 9444 284260 9450
rect 284208 9386 284260 9392
rect 283104 9308 283156 9314
rect 283104 9250 283156 9256
rect 282828 5296 282880 5302
rect 282828 5238 282880 5244
rect 282276 5024 282328 5030
rect 281828 4950 282040 4978
rect 282328 4972 282408 4978
rect 282276 4966 282408 4972
rect 281828 4758 281856 4950
rect 282012 4944 282040 4950
rect 282092 4956 282144 4962
rect 282012 4916 282092 4944
rect 282288 4950 282408 4966
rect 282092 4898 282144 4904
rect 281908 4888 281960 4894
rect 281908 4830 281960 4836
rect 281816 4752 281868 4758
rect 281816 4694 281868 4700
rect 281920 480 281948 4830
rect 282380 4758 282408 4950
rect 282368 4752 282420 4758
rect 282368 4694 282420 4700
rect 283116 480 283144 9250
rect 284300 5228 284352 5234
rect 284300 5170 284352 5176
rect 284312 480 284340 5170
rect 284956 490 284984 13262
rect 285508 6497 285536 30466
rect 285494 6488 285550 6497
rect 285494 6423 285550 6432
rect 285600 5234 285628 30602
rect 286428 30530 286456 34054
rect 286416 30524 286468 30530
rect 286416 30466 286468 30472
rect 286600 9376 286652 9382
rect 286600 9318 286652 9324
rect 285588 5228 285640 5234
rect 285588 5170 285640 5176
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 9318
rect 286888 9314 286916 34054
rect 287532 30530 287560 34054
rect 288084 30666 288112 34054
rect 288268 34054 288328 34082
rect 288880 34054 289216 34082
rect 289432 34054 289768 34082
rect 289984 34054 290320 34082
rect 290536 34054 290964 34082
rect 288072 30660 288124 30666
rect 288072 30602 288124 30608
rect 286968 30524 287020 30530
rect 286968 30466 287020 30472
rect 287520 30524 287572 30530
rect 287520 30466 287572 30472
rect 288164 30524 288216 30530
rect 288164 30466 288216 30472
rect 286876 9308 286928 9314
rect 286876 9250 286928 9256
rect 286980 5166 287008 30466
rect 288176 13161 288204 30466
rect 288162 13152 288218 13161
rect 288162 13087 288218 13096
rect 287336 11144 287388 11150
rect 287336 11086 287388 11092
rect 286968 5160 287020 5166
rect 286968 5102 287020 5108
rect 287348 490 287376 11086
rect 288268 8945 288296 34054
rect 288348 30660 288400 30666
rect 288348 30602 288400 30608
rect 288254 8936 288310 8945
rect 288254 8871 288310 8880
rect 288360 5098 288388 30602
rect 289188 30530 289216 34054
rect 289176 30524 289228 30530
rect 289176 30466 289228 30472
rect 289636 30524 289688 30530
rect 289636 30466 289688 30472
rect 289648 13258 289676 30466
rect 288992 13252 289044 13258
rect 288992 13194 289044 13200
rect 289636 13252 289688 13258
rect 289636 13194 289688 13200
rect 288348 5092 288400 5098
rect 288348 5034 288400 5040
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 13194
rect 289740 5137 289768 34054
rect 290292 30530 290320 34054
rect 290280 30524 290332 30530
rect 290280 30466 290332 30472
rect 290936 14550 290964 34054
rect 291074 33810 291102 34068
rect 291640 34054 291976 34082
rect 292192 34054 292528 34082
rect 292836 34054 293172 34082
rect 293388 34054 293816 34082
rect 291074 33782 291148 33810
rect 291016 30524 291068 30530
rect 291016 30466 291068 30472
rect 290924 14544 290976 14550
rect 290924 14486 290976 14492
rect 290188 9240 290240 9246
rect 290188 9182 290240 9188
rect 289726 5128 289782 5137
rect 289726 5063 289782 5072
rect 290200 480 290228 9182
rect 291028 6361 291056 30466
rect 291014 6352 291070 6361
rect 291014 6287 291070 6296
rect 291120 5001 291148 33782
rect 291948 30530 291976 34054
rect 291936 30524 291988 30530
rect 291936 30466 291988 30472
rect 292396 30524 292448 30530
rect 292396 30466 292448 30472
rect 292408 14482 292436 30466
rect 292500 14793 292528 34054
rect 293144 30666 293172 34054
rect 293132 30660 293184 30666
rect 293132 30602 293184 30608
rect 293684 30524 293736 30530
rect 293684 30466 293736 30472
rect 292486 14784 292542 14793
rect 292486 14719 292542 14728
rect 292396 14476 292448 14482
rect 292396 14418 292448 14424
rect 293696 13025 293724 30466
rect 293682 13016 293738 13025
rect 293682 12951 293738 12960
rect 293788 9246 293816 34054
rect 293880 34054 293940 34082
rect 294492 34054 294828 34082
rect 295044 34054 295196 34082
rect 295596 34054 295932 34082
rect 296148 34054 296576 34082
rect 293880 30530 293908 34054
rect 293960 30660 294012 30666
rect 293960 30602 294012 30608
rect 293868 30524 293920 30530
rect 293868 30466 293920 30472
rect 293972 30410 294000 30602
rect 294800 30530 294828 34054
rect 294788 30524 294840 30530
rect 294788 30466 294840 30472
rect 293880 30382 294000 30410
rect 293776 9240 293828 9246
rect 293776 9182 293828 9188
rect 293684 9172 293736 9178
rect 293684 9114 293736 9120
rect 291106 4992 291162 5001
rect 291106 4927 291162 4936
rect 291384 4888 291436 4894
rect 291384 4830 291436 4836
rect 291396 480 291424 4830
rect 292580 4820 292632 4826
rect 292580 4762 292632 4768
rect 292592 480 292620 4762
rect 293696 480 293724 9114
rect 293880 4826 293908 30382
rect 295168 9178 295196 34054
rect 295904 30530 295932 34054
rect 295248 30524 295300 30530
rect 295248 30466 295300 30472
rect 295892 30524 295944 30530
rect 295892 30466 295944 30472
rect 296444 30524 296496 30530
rect 296444 30466 296496 30472
rect 295156 9172 295208 9178
rect 295156 9114 295208 9120
rect 295260 4962 295288 30466
rect 296456 12510 296484 30466
rect 296548 30138 296576 34054
rect 296640 34054 296700 34082
rect 297252 34054 297680 34082
rect 297804 34054 298048 34082
rect 298356 34054 298692 34082
rect 298908 34054 299244 34082
rect 296640 30258 296668 34054
rect 296628 30252 296680 30258
rect 296628 30194 296680 30200
rect 296548 30110 296668 30138
rect 296536 30048 296588 30054
rect 296536 29990 296588 29996
rect 295616 12504 295668 12510
rect 295616 12446 295668 12452
rect 296444 12504 296496 12510
rect 296444 12446 296496 12452
rect 294880 4956 294932 4962
rect 294880 4898 294932 4904
rect 295248 4956 295300 4962
rect 295248 4898 295300 4904
rect 293868 4820 293920 4826
rect 293868 4762 293920 4768
rect 294892 480 294920 4898
rect 295628 490 295656 12446
rect 296548 6225 296576 29990
rect 296534 6216 296590 6225
rect 296534 6151 296590 6160
rect 296640 4894 296668 30110
rect 297652 26234 297680 34054
rect 297652 26206 297956 26234
rect 297928 14657 297956 26206
rect 297914 14648 297970 14657
rect 297914 14583 297970 14592
rect 297272 9036 297324 9042
rect 297272 8978 297324 8984
rect 296628 4888 296680 4894
rect 296628 4830 296680 4836
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 8978
rect 298020 4865 298048 34054
rect 298664 30530 298692 34054
rect 298652 30524 298704 30530
rect 298652 30466 298704 30472
rect 299216 14521 299244 34054
rect 299400 34054 299460 34082
rect 300012 34054 300440 34082
rect 300564 34054 300808 34082
rect 301116 34054 301452 34082
rect 301668 34054 302004 34082
rect 299296 30524 299348 30530
rect 299296 30466 299348 30472
rect 299202 14512 299258 14521
rect 299202 14447 299258 14456
rect 299308 9042 299336 30466
rect 299296 9036 299348 9042
rect 299296 8978 299348 8984
rect 299400 5030 299428 34054
rect 300412 26234 300440 34054
rect 300412 26206 300716 26234
rect 300688 13190 300716 26206
rect 299664 13184 299716 13190
rect 299664 13126 299716 13132
rect 300676 13184 300728 13190
rect 300676 13126 300728 13132
rect 298468 5024 298520 5030
rect 298468 4966 298520 4972
rect 299388 5024 299440 5030
rect 299388 4966 299440 4972
rect 298006 4856 298062 4865
rect 298006 4791 298062 4800
rect 298480 480 298508 4966
rect 299676 480 299704 13126
rect 300780 12730 300808 34054
rect 301424 30666 301452 34054
rect 301504 30728 301556 30734
rect 301504 30670 301556 30676
rect 301412 30660 301464 30666
rect 301412 30602 301464 30608
rect 300688 12702 300808 12730
rect 300688 9042 300716 12702
rect 300676 9036 300728 9042
rect 300676 8978 300728 8984
rect 300768 8968 300820 8974
rect 300768 8910 300820 8916
rect 300780 480 300808 8910
rect 301516 6866 301544 30670
rect 301976 30530 302004 34054
rect 302160 34054 302220 34082
rect 302160 31385 302188 34054
rect 302896 33114 302924 310490
rect 302974 309496 303030 309505
rect 302974 309431 303030 309440
rect 302988 46918 303016 309431
rect 303080 86970 303108 312015
rect 303160 310276 303212 310282
rect 303160 310218 303212 310224
rect 303172 167006 303200 310218
rect 303160 167000 303212 167006
rect 303160 166942 303212 166948
rect 303264 126954 303292 312151
rect 303344 310344 303396 310350
rect 303344 310286 303396 310292
rect 303356 206990 303384 310286
rect 303448 259418 303476 312938
rect 303528 312928 303580 312934
rect 303528 312870 303580 312876
rect 303540 273222 303568 312870
rect 304446 312352 304502 312361
rect 304446 312287 304502 312296
rect 304356 310208 304408 310214
rect 304356 310150 304408 310156
rect 304264 310072 304316 310078
rect 304264 310014 304316 310020
rect 303528 273216 303580 273222
rect 303528 273158 303580 273164
rect 303436 259412 303488 259418
rect 303436 259354 303488 259360
rect 303344 206984 303396 206990
rect 303344 206926 303396 206932
rect 303252 126948 303304 126954
rect 303252 126890 303304 126896
rect 303068 86964 303120 86970
rect 303068 86906 303120 86912
rect 304276 73166 304304 310014
rect 304368 153202 304396 310150
rect 304460 233238 304488 312287
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 304632 310480 304684 310486
rect 304632 310422 304684 310428
rect 304540 310412 304592 310418
rect 304540 310354 304592 310360
rect 304552 245614 304580 310354
rect 304644 299470 304672 310422
rect 580908 309596 580960 309602
rect 580908 309538 580960 309544
rect 580724 309528 580776 309534
rect 580724 309470 580776 309476
rect 580632 309392 580684 309398
rect 315302 309360 315358 309369
rect 580632 309334 580684 309340
rect 315302 309295 315358 309304
rect 580448 309324 580500 309330
rect 304632 299464 304684 299470
rect 304632 299406 304684 299412
rect 304540 245608 304592 245614
rect 304540 245550 304592 245556
rect 304448 233232 304500 233238
rect 304448 233174 304500 233180
rect 304356 153196 304408 153202
rect 304356 153138 304408 153144
rect 304264 73160 304316 73166
rect 304264 73102 304316 73108
rect 302976 46912 303028 46918
rect 302976 46854 303028 46860
rect 302884 33108 302936 33114
rect 302884 33050 302936 33056
rect 302146 31376 302202 31385
rect 302146 31311 302202 31320
rect 308404 30660 308456 30666
rect 308404 30602 308456 30608
rect 301964 30524 302016 30530
rect 301964 30466 302016 30472
rect 304264 30524 304316 30530
rect 304264 30466 304316 30472
rect 304276 13122 304304 30466
rect 307760 13864 307812 13870
rect 307760 13806 307812 13812
rect 303160 13116 303212 13122
rect 303160 13058 303212 13064
rect 304264 13116 304316 13122
rect 304264 13058 304316 13064
rect 301412 6860 301464 6866
rect 301412 6802 301464 6808
rect 301504 6860 301556 6866
rect 301504 6802 301556 6808
rect 301424 490 301452 6802
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301424 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 13058
rect 306380 12640 306432 12646
rect 306380 12582 306432 12588
rect 305552 9716 305604 9722
rect 305552 9658 305604 9664
rect 304356 8356 304408 8362
rect 304356 8298 304408 8304
rect 304368 480 304396 8298
rect 305564 480 305592 9658
rect 306392 490 306420 12582
rect 307772 3126 307800 13806
rect 308416 9110 308444 30602
rect 309784 30592 309836 30598
rect 309784 30534 309836 30540
rect 309692 12572 309744 12578
rect 309692 12514 309744 12520
rect 307944 9104 307996 9110
rect 307944 9046 307996 9052
rect 308404 9104 308456 9110
rect 308404 9046 308456 9052
rect 307760 3120 307812 3126
rect 307760 3062 307812 3068
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 9046
rect 309048 3120 309100 3126
rect 309048 3062 309100 3068
rect 309060 480 309088 3062
rect 309704 490 309732 12514
rect 309796 3126 309824 30534
rect 312544 30388 312596 30394
rect 312544 30330 312596 30336
rect 311440 8424 311492 8430
rect 311440 8366 311492 8372
rect 309784 3120 309836 3126
rect 309784 3062 309836 3068
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309704 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 8366
rect 312556 2854 312584 30330
rect 313832 12708 313884 12714
rect 313832 12650 313884 12656
rect 312636 6860 312688 6866
rect 312636 6802 312688 6808
rect 312544 2848 312596 2854
rect 312544 2790 312596 2796
rect 312648 480 312676 6802
rect 313844 480 313872 12650
rect 315026 9344 315082 9353
rect 315026 9279 315082 9288
rect 315040 480 315068 9279
rect 315316 6866 315344 309295
rect 580448 309266 580500 309272
rect 580262 309224 580318 309233
rect 580262 309159 580318 309168
rect 580356 309188 580408 309194
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 579988 273216 580040 273222
rect 579988 273158 580040 273164
rect 580000 272241 580028 273158
rect 579986 272232 580042 272241
rect 579986 272167 580042 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 579620 167000 579672 167006
rect 579620 166942 579672 166948
rect 579632 165889 579660 166942
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 579712 126948 579764 126954
rect 579712 126890 579764 126896
rect 579724 126041 579752 126890
rect 579710 126032 579766 126041
rect 579710 125967 579766 125976
rect 579620 86964 579672 86970
rect 579620 86906 579672 86912
rect 579632 86193 579660 86906
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 358084 31748 358136 31754
rect 358084 31690 358136 31696
rect 344284 31680 344336 31686
rect 344284 31622 344336 31628
rect 330484 31612 330536 31618
rect 330484 31554 330536 31560
rect 322202 31376 322258 31385
rect 322202 31311 322258 31320
rect 315396 30456 315448 30462
rect 315396 30398 315448 30404
rect 315304 6860 315356 6866
rect 315304 6802 315356 6808
rect 315408 2990 315436 30398
rect 316040 13932 316092 13938
rect 316040 13874 316092 13880
rect 316052 3482 316080 13874
rect 317328 12776 317380 12782
rect 317328 12718 317380 12724
rect 316052 3454 316264 3482
rect 315396 2984 315448 2990
rect 315396 2926 315448 2932
rect 316236 480 316264 3454
rect 317340 480 317368 12718
rect 318522 9208 318578 9217
rect 318522 9143 318578 9152
rect 318536 480 318564 9143
rect 322110 9072 322166 9081
rect 322110 9007 322166 9016
rect 319720 6996 319772 7002
rect 319720 6938 319772 6944
rect 319732 480 319760 6938
rect 320916 6180 320968 6186
rect 320916 6122 320968 6128
rect 320928 480 320956 6122
rect 322124 480 322152 9007
rect 322216 6186 322244 31311
rect 323582 31240 323638 31249
rect 323582 31175 323638 31184
rect 322204 6180 322256 6186
rect 322204 6122 322256 6128
rect 323596 3641 323624 31175
rect 323676 30796 323728 30802
rect 323676 30738 323728 30744
rect 323582 3632 323638 3641
rect 323582 3567 323638 3576
rect 323688 2922 323716 30738
rect 328736 14136 328788 14142
rect 328736 14078 328788 14084
rect 326344 14068 326396 14074
rect 326344 14010 326396 14016
rect 324320 14000 324372 14006
rect 324320 13942 324372 13948
rect 323308 2916 323360 2922
rect 323308 2858 323360 2864
rect 323676 2916 323728 2922
rect 323676 2858 323728 2864
rect 323320 480 323348 2858
rect 324332 2786 324360 13942
rect 324412 5568 324464 5574
rect 324412 5510 324464 5516
rect 324320 2780 324372 2786
rect 324320 2722 324372 2728
rect 324424 480 324452 5510
rect 325608 2780 325660 2786
rect 325608 2722 325660 2728
rect 325620 480 325648 2722
rect 326356 490 326384 14010
rect 328000 5636 328052 5642
rect 328000 5578 328052 5584
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 5578
rect 328748 490 328776 14078
rect 330496 3058 330524 31554
rect 341524 31204 341576 31210
rect 341524 31146 341576 31152
rect 337384 31000 337436 31006
rect 337384 30942 337436 30948
rect 333244 30864 333296 30870
rect 333244 30806 333296 30812
rect 332692 14204 332744 14210
rect 332692 14146 332744 14152
rect 331588 5704 331640 5710
rect 331588 5646 331640 5652
rect 330392 3052 330444 3058
rect 330392 2994 330444 3000
rect 330484 3052 330536 3058
rect 330484 2994 330536 3000
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 2994
rect 331600 480 331628 5646
rect 332704 480 332732 14146
rect 333256 3058 333284 30806
rect 337396 16574 337424 30942
rect 337396 16546 337608 16574
rect 336280 14272 336332 14278
rect 336280 14214 336332 14220
rect 335084 5772 335136 5778
rect 335084 5714 335136 5720
rect 333244 3052 333296 3058
rect 333244 2994 333296 3000
rect 333888 2916 333940 2922
rect 333888 2858 333940 2864
rect 333900 480 333928 2858
rect 335096 480 335124 5714
rect 336292 480 336320 14214
rect 337580 3194 337608 16546
rect 339500 9784 339552 9790
rect 339500 9726 339552 9732
rect 338672 5840 338724 5846
rect 338672 5782 338724 5788
rect 337476 3188 337528 3194
rect 337476 3130 337528 3136
rect 337568 3188 337620 3194
rect 337568 3130 337620 3136
rect 337488 480 337516 3130
rect 338684 480 338712 5782
rect 339512 490 339540 9726
rect 341536 2922 341564 31146
rect 342904 9852 342956 9858
rect 342904 9794 342956 9800
rect 342168 5908 342220 5914
rect 342168 5850 342220 5856
rect 340972 2916 341024 2922
rect 340972 2858 341024 2864
rect 341524 2916 341576 2922
rect 341524 2858 341576 2864
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 2858
rect 342180 480 342208 5850
rect 342916 490 342944 9794
rect 344296 3194 344324 31622
rect 355324 31340 355376 31346
rect 355324 31282 355376 31288
rect 348424 31272 348476 31278
rect 348424 31214 348476 31220
rect 346952 9920 347004 9926
rect 346952 9862 347004 9868
rect 345756 5976 345808 5982
rect 345756 5918 345808 5924
rect 344560 3256 344612 3262
rect 344560 3198 344612 3204
rect 344284 3188 344336 3194
rect 344284 3130 344336 3136
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3198
rect 345768 480 345796 5918
rect 346964 480 346992 9862
rect 348436 3233 348464 31214
rect 351184 30932 351236 30938
rect 351184 30874 351236 30880
rect 349160 9988 349212 9994
rect 349160 9930 349212 9936
rect 349172 3330 349200 9930
rect 349252 6044 349304 6050
rect 349252 5986 349304 5992
rect 349160 3324 349212 3330
rect 349160 3266 349212 3272
rect 348422 3224 348478 3233
rect 348422 3159 348478 3168
rect 348056 3052 348108 3058
rect 348056 2994 348108 3000
rect 348068 480 348096 2994
rect 349264 480 349292 5986
rect 351196 3330 351224 30874
rect 353576 10056 353628 10062
rect 353576 9998 353628 10004
rect 352840 6112 352892 6118
rect 352840 6054 352892 6060
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 351184 3324 351236 3330
rect 351184 3266 351236 3272
rect 351828 3324 351880 3330
rect 351828 3266 351880 3272
rect 350460 480 350488 3266
rect 351644 3256 351696 3262
rect 351840 3233 351868 3266
rect 351644 3198 351696 3204
rect 351826 3224 351882 3233
rect 351656 480 351684 3198
rect 351826 3159 351882 3168
rect 352852 480 352880 6054
rect 353588 490 353616 9998
rect 355336 2922 355364 31282
rect 357532 10124 357584 10130
rect 357532 10066 357584 10072
rect 356334 5264 356390 5273
rect 356334 5199 356390 5208
rect 355968 3392 356020 3398
rect 355888 3340 355968 3346
rect 355888 3334 356020 3340
rect 355888 3318 356008 3334
rect 355888 3262 355916 3318
rect 355876 3256 355928 3262
rect 355876 3198 355928 3204
rect 355232 2916 355284 2922
rect 355232 2858 355284 2864
rect 355324 2916 355376 2922
rect 355324 2858 355376 2864
rect 353864 598 354076 626
rect 353864 490 353892 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 462 353892 490
rect 354048 480 354076 598
rect 355244 480 355272 2858
rect 356348 480 356376 5199
rect 357544 480 357572 10066
rect 358096 3398 358124 31690
rect 362224 31544 362276 31550
rect 362224 31486 362276 31492
rect 362236 16574 362264 31486
rect 376024 31476 376076 31482
rect 376024 31418 376076 31424
rect 369124 31408 369176 31414
rect 369124 31350 369176 31356
rect 366364 31136 366416 31142
rect 366364 31078 366416 31084
rect 362236 16546 362448 16574
rect 361120 10192 361172 10198
rect 361120 10134 361172 10140
rect 359924 6792 359976 6798
rect 359924 6734 359976 6740
rect 358084 3392 358136 3398
rect 358084 3334 358136 3340
rect 358728 2916 358780 2922
rect 358728 2858 358780 2864
rect 358740 480 358768 2858
rect 359936 480 359964 6734
rect 361132 480 361160 10134
rect 362420 3058 362448 16546
rect 364616 10260 364668 10266
rect 364616 10202 364668 10208
rect 363512 6724 363564 6730
rect 363512 6666 363564 6672
rect 362316 3052 362368 3058
rect 362316 2994 362368 3000
rect 362408 3052 362460 3058
rect 362408 2994 362460 3000
rect 362328 480 362356 2994
rect 363524 480 363552 6666
rect 364628 480 364656 10202
rect 366376 4146 366404 31078
rect 369136 16574 369164 31350
rect 373264 31068 373316 31074
rect 373264 31010 373316 31016
rect 369136 16546 369532 16574
rect 367744 11008 367796 11014
rect 367744 10950 367796 10956
rect 367008 6656 367060 6662
rect 367008 6598 367060 6604
rect 365812 4140 365864 4146
rect 365812 4082 365864 4088
rect 366364 4140 366416 4146
rect 366364 4082 366416 4088
rect 365824 480 365852 4082
rect 367020 480 367048 6598
rect 367756 490 367784 10950
rect 369504 3398 369532 16546
rect 370136 12844 370188 12850
rect 370136 12786 370188 12792
rect 369492 3392 369544 3398
rect 369492 3334 369544 3340
rect 369400 3256 369452 3262
rect 369400 3198 369452 3204
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 3198
rect 370148 490 370176 12786
rect 371240 10940 371292 10946
rect 371240 10882 371292 10888
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371252 490 371280 10882
rect 372896 4072 372948 4078
rect 372896 4014 372948 4020
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 370566 -960 370678 480
rect 371252 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 4014
rect 373276 3398 373304 31010
rect 376036 16574 376064 31418
rect 382922 31104 382978 31113
rect 382922 31039 382978 31048
rect 380162 30968 380218 30977
rect 380162 30903 380218 30912
rect 376036 16546 376616 16574
rect 374092 12912 374144 12918
rect 374092 12854 374144 12860
rect 373264 3392 373316 3398
rect 373264 3334 373316 3340
rect 374104 480 374132 12854
rect 375288 10872 375340 10878
rect 375288 10814 375340 10820
rect 375300 480 375328 10814
rect 376588 4078 376616 16546
rect 377680 14340 377732 14346
rect 377680 14282 377732 14288
rect 376484 4072 376536 4078
rect 376484 4014 376536 4020
rect 376576 4072 376628 4078
rect 376576 4014 376628 4020
rect 376496 480 376524 4014
rect 377692 480 377720 14282
rect 378416 10804 378468 10810
rect 378416 10746 378468 10752
rect 378428 490 378456 10746
rect 380176 4078 380204 30903
rect 381176 14408 381228 14414
rect 381176 14350 381228 14356
rect 380164 4072 380216 4078
rect 380164 4014 380216 4020
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 3946
rect 381188 480 381216 14350
rect 382372 10736 382424 10742
rect 382372 10678 382424 10684
rect 382384 480 382412 10678
rect 382936 4010 382964 31039
rect 580276 19825 580304 309159
rect 580356 309130 580408 309136
rect 580368 59673 580396 309130
rect 580460 99521 580488 309266
rect 580540 309256 580592 309262
rect 580540 309198 580592 309204
rect 580552 112849 580580 309198
rect 580644 139369 580672 309334
rect 580736 179217 580764 309470
rect 580816 309460 580868 309466
rect 580816 309402 580868 309408
rect 580828 192545 580856 309402
rect 580920 219065 580948 309538
rect 580906 219056 580962 219065
rect 580906 218991 580962 219000
rect 580814 192536 580870 192545
rect 580814 192471 580870 192480
rect 580722 179208 580778 179217
rect 580722 179143 580778 179152
rect 580630 139360 580686 139369
rect 580630 139295 580686 139304
rect 580538 112840 580594 112849
rect 580538 112775 580594 112784
rect 580446 99512 580502 99521
rect 580446 99447 580502 99456
rect 580354 59664 580410 59673
rect 580354 59599 580410 59608
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 436744 16108 436796 16114
rect 436744 16050 436796 16056
rect 420920 15156 420972 15162
rect 420920 15098 420972 15104
rect 418804 12504 418856 12510
rect 418804 12446 418856 12452
rect 407210 10704 407266 10713
rect 385960 10668 386012 10674
rect 407210 10639 407266 10648
rect 385960 10610 386012 10616
rect 384764 7064 384816 7070
rect 384764 7006 384816 7012
rect 383476 4140 383528 4146
rect 383476 4082 383528 4088
rect 382924 4004 382976 4010
rect 382924 3946 382976 3952
rect 383488 3754 383516 4082
rect 383488 3726 383608 3754
rect 383580 3330 383608 3726
rect 383476 3324 383528 3330
rect 383476 3266 383528 3272
rect 383568 3324 383620 3330
rect 383568 3266 383620 3272
rect 383488 1714 383516 3266
rect 383488 1686 383608 1714
rect 383580 480 383608 1686
rect 384776 480 384804 7006
rect 385972 480 386000 10610
rect 389456 10600 389508 10606
rect 389456 10542 389508 10548
rect 388260 7132 388312 7138
rect 388260 7074 388312 7080
rect 387156 3936 387208 3942
rect 387156 3878 387208 3884
rect 387168 480 387196 3878
rect 388272 480 388300 7074
rect 389468 480 389496 10542
rect 392584 10532 392636 10538
rect 392584 10474 392636 10480
rect 391848 7200 391900 7206
rect 391848 7142 391900 7148
rect 390652 2916 390704 2922
rect 390652 2858 390704 2864
rect 390664 480 390692 2858
rect 391860 480 391888 7142
rect 392596 490 392624 10474
rect 396080 10464 396132 10470
rect 396080 10406 396132 10412
rect 395344 7268 395396 7274
rect 395344 7210 395396 7216
rect 394240 3868 394292 3874
rect 394240 3810 394292 3816
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 3810
rect 395356 480 395384 7210
rect 396092 490 396120 10406
rect 398840 10396 398892 10402
rect 398840 10338 398892 10344
rect 398852 3806 398880 10338
rect 403624 10328 403676 10334
rect 403624 10270 403676 10276
rect 402520 7404 402572 7410
rect 402520 7346 402572 7352
rect 398932 7336 398984 7342
rect 398932 7278 398984 7284
rect 398840 3800 398892 3806
rect 398840 3742 398892 3748
rect 397736 3052 397788 3058
rect 397736 2994 397788 3000
rect 396368 598 396580 626
rect 396368 490 396396 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 2994
rect 398944 480 398972 7278
rect 401324 3868 401376 3874
rect 401324 3810 401376 3816
rect 400128 3800 400180 3806
rect 400128 3742 400180 3748
rect 400140 480 400168 3742
rect 401336 480 401364 3810
rect 402532 480 402560 7346
rect 403636 480 403664 10270
rect 406016 7540 406068 7546
rect 406016 7482 406068 7488
rect 404820 3188 404872 3194
rect 404820 3130 404872 3136
rect 404832 480 404860 3130
rect 406028 480 406056 7482
rect 407224 480 407252 10639
rect 410798 10568 410854 10577
rect 410798 10503 410854 10512
rect 409604 7472 409656 7478
rect 409604 7414 409656 7420
rect 408408 3732 408460 3738
rect 408408 3674 408460 3680
rect 408420 480 408448 3674
rect 409616 480 409644 7414
rect 410812 480 410840 10503
rect 414294 10432 414350 10441
rect 414294 10367 414350 10376
rect 413100 8288 413152 8294
rect 413100 8230 413152 8236
rect 411904 3256 411956 3262
rect 411904 3198 411956 3204
rect 411916 480 411944 3198
rect 413112 480 413140 8230
rect 414308 480 414336 10367
rect 417422 10296 417478 10305
rect 417422 10231 417478 10240
rect 416688 8220 416740 8226
rect 416688 8162 416740 8168
rect 415492 3664 415544 3670
rect 415492 3606 415544 3612
rect 415504 480 415532 3606
rect 416700 480 416728 8162
rect 417436 490 417464 10231
rect 418816 3670 418844 12446
rect 420184 8152 420236 8158
rect 420184 8094 420236 8100
rect 418804 3664 418856 3670
rect 418804 3606 418856 3612
rect 418988 3324 419040 3330
rect 418988 3266 419040 3272
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 419000 480 419028 3266
rect 420196 480 420224 8094
rect 420932 490 420960 15098
rect 423680 15088 423732 15094
rect 423680 15030 423732 15036
rect 422576 3596 422628 3602
rect 422576 3538 422628 3544
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 3538
rect 423692 3534 423720 15030
rect 428464 15020 428516 15026
rect 428464 14962 428516 14968
rect 427268 8084 427320 8090
rect 427268 8026 427320 8032
rect 423772 8016 423824 8022
rect 423772 7958 423824 7964
rect 423680 3528 423732 3534
rect 423680 3470 423732 3476
rect 423784 480 423812 7958
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 424980 480 425008 3470
rect 426164 3392 426216 3398
rect 426164 3334 426216 3340
rect 426176 480 426204 3334
rect 427280 480 427308 8026
rect 428476 480 428504 14962
rect 432052 14952 432104 14958
rect 432052 14894 432104 14900
rect 430856 7948 430908 7954
rect 430856 7890 430908 7896
rect 429660 3596 429712 3602
rect 429660 3538 429712 3544
rect 429672 480 429700 3538
rect 430868 480 430896 7890
rect 432064 480 432092 14894
rect 435088 14884 435140 14890
rect 435088 14826 435140 14832
rect 434444 7880 434496 7886
rect 434444 7822 434496 7828
rect 433248 4140 433300 4146
rect 433248 4082 433300 4088
rect 433260 480 433288 4082
rect 434456 480 434484 7822
rect 435100 490 435128 14826
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 16050
rect 450912 16040 450964 16046
rect 450912 15982 450964 15988
rect 448520 11348 448572 11354
rect 448520 11290 448572 11296
rect 445760 11280 445812 11286
rect 445760 11222 445812 11228
rect 439136 11212 439188 11218
rect 439136 11154 439188 11160
rect 437940 7812 437992 7818
rect 437940 7754 437992 7760
rect 437952 480 437980 7754
rect 439148 480 439176 11154
rect 445022 7984 445078 7993
rect 445022 7919 445078 7928
rect 441528 7744 441580 7750
rect 441528 7686 441580 7692
rect 440332 2848 440384 2854
rect 440332 2790 440384 2796
rect 440344 480 440372 2790
rect 441540 480 441568 7686
rect 442632 6588 442684 6594
rect 442632 6530 442684 6536
rect 442644 480 442672 6530
rect 443828 3460 443880 3466
rect 443828 3402 443880 3408
rect 443840 480 443868 3402
rect 445036 480 445064 7919
rect 445772 490 445800 11222
rect 447416 4072 447468 4078
rect 447416 4014 447468 4020
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 4014
rect 448532 3534 448560 11290
rect 448610 7848 448666 7857
rect 448610 7783 448666 7792
rect 448520 3528 448572 3534
rect 448520 3470 448572 3476
rect 448624 480 448652 7783
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 449820 480 449848 3470
rect 450924 480 450952 15982
rect 456800 15972 456852 15978
rect 456800 15914 456852 15920
rect 453304 11416 453356 11422
rect 453304 11358 453356 11364
rect 452106 7712 452162 7721
rect 452106 7647 452162 7656
rect 452120 480 452148 7647
rect 453316 480 453344 11358
rect 455696 7676 455748 7682
rect 455696 7618 455748 7624
rect 454500 2984 454552 2990
rect 454500 2926 454552 2932
rect 454512 480 454540 2926
rect 455708 480 455736 7618
rect 456812 3534 456840 15914
rect 465172 15904 465224 15910
rect 465172 15846 465224 15852
rect 463976 11620 464028 11626
rect 463976 11562 464028 11568
rect 459928 11552 459980 11558
rect 459928 11494 459980 11500
rect 456892 11484 456944 11490
rect 456892 11426 456944 11432
rect 456800 3528 456852 3534
rect 456800 3470 456852 3476
rect 456904 480 456932 11426
rect 459192 7608 459244 7614
rect 459192 7550 459244 7556
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 458100 480 458128 3470
rect 459204 480 459232 7550
rect 459940 490 459968 11494
rect 462778 7576 462834 7585
rect 462778 7511 462834 7520
rect 461584 3120 461636 3126
rect 461584 3062 461636 3068
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3062
rect 462792 480 462820 7511
rect 463988 480 464016 11562
rect 465184 480 465212 15846
rect 465816 14816 465868 14822
rect 465816 14758 465868 14764
rect 560390 14784 560446 14793
rect 465828 490 465856 14758
rect 469864 14748 469916 14754
rect 560390 14719 560446 14728
rect 469864 14690 469916 14696
rect 467472 11688 467524 11694
rect 467472 11630 467524 11636
rect 466104 598 466316 626
rect 466104 490 466132 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 462 466132 490
rect 466288 480 466316 598
rect 467484 480 467512 11630
rect 468666 3632 468722 3641
rect 468666 3567 468722 3576
rect 468680 480 468708 3567
rect 469876 480 469904 14690
rect 476488 14680 476540 14686
rect 476488 14622 476540 14628
rect 473452 14612 473504 14618
rect 473452 14554 473504 14560
rect 470600 12436 470652 12442
rect 470600 12378 470652 12384
rect 470612 490 470640 12378
rect 472254 3496 472310 3505
rect 472254 3431 472310 3440
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 3431
rect 473464 480 473492 14554
rect 474096 12368 474148 12374
rect 474096 12310 474148 12316
rect 474108 490 474136 12310
rect 475752 4004 475804 4010
rect 475752 3946 475804 3952
rect 474384 598 474596 626
rect 474384 490 474412 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 462 474412 490
rect 474568 480 474596 598
rect 475764 480 475792 3946
rect 476500 490 476528 14622
rect 556896 14544 556948 14550
rect 556896 14486 556948 14492
rect 487160 13796 487212 13802
rect 487160 13738 487212 13744
rect 484032 13048 484084 13054
rect 484032 12990 484084 12996
rect 480536 12980 480588 12986
rect 480536 12922 480588 12928
rect 478144 12300 478196 12306
rect 478144 12242 478196 12248
rect 476776 598 476988 626
rect 476776 490 476804 598
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 462 476804 490
rect 476960 480 476988 598
rect 478156 480 478184 12242
rect 479338 3360 479394 3369
rect 479338 3295 479394 3304
rect 479352 480 479380 3295
rect 480548 480 480576 12922
rect 482376 12232 482428 12238
rect 482376 12174 482428 12180
rect 481732 8492 481784 8498
rect 481732 8434 481784 8440
rect 481744 480 481772 8434
rect 482388 490 482416 12174
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 12990
rect 486424 12164 486476 12170
rect 486424 12106 486476 12112
rect 485228 8560 485280 8566
rect 485228 8502 485280 8508
rect 485240 480 485268 8502
rect 486436 480 486464 12106
rect 487172 490 487200 13738
rect 489920 13728 489972 13734
rect 489920 13670 489972 13676
rect 488816 8628 488868 8634
rect 488816 8570 488868 8576
rect 487448 598 487660 626
rect 487448 490 487476 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 462 487476 490
rect 487632 480 487660 598
rect 488828 480 488856 8570
rect 489932 3602 489960 13670
rect 494704 13660 494756 13666
rect 494704 13602 494756 13608
rect 490012 12096 490064 12102
rect 490012 12038 490064 12044
rect 489920 3596 489972 3602
rect 489920 3538 489972 3544
rect 490024 3482 490052 12038
rect 493048 12028 493100 12034
rect 493048 11970 493100 11976
rect 492312 6520 492364 6526
rect 492312 6462 492364 6468
rect 491116 3596 491168 3602
rect 491116 3538 491168 3544
rect 489932 3454 490052 3482
rect 489932 480 489960 3454
rect 491128 480 491156 3538
rect 492324 480 492352 6462
rect 493060 490 493088 11970
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 13602
rect 525432 13592 525484 13598
rect 525432 13534 525484 13540
rect 511262 12064 511318 12073
rect 511262 11999 511318 12008
rect 497096 11960 497148 11966
rect 497096 11902 497148 11908
rect 495900 8696 495952 8702
rect 495900 8638 495952 8644
rect 495912 480 495940 8638
rect 497108 480 497136 11902
rect 500592 11892 500644 11898
rect 500592 11834 500644 11840
rect 499396 8764 499448 8770
rect 499396 8706 499448 8712
rect 498200 4208 498252 4214
rect 498200 4150 498252 4156
rect 498212 480 498240 4150
rect 499408 480 499436 8706
rect 500604 480 500632 11834
rect 503720 11824 503772 11830
rect 503720 11766 503772 11772
rect 502984 6452 503036 6458
rect 502984 6394 503036 6400
rect 501788 4276 501840 4282
rect 501788 4218 501840 4224
rect 501800 480 501828 4218
rect 502996 480 503024 6394
rect 503732 490 503760 11766
rect 507216 11756 507268 11762
rect 507216 11698 507268 11704
rect 506480 8832 506532 8838
rect 506480 8774 506532 8780
rect 505376 4344 505428 4350
rect 505376 4286 505428 4292
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 4286
rect 506492 480 506520 8774
rect 507228 490 507256 11698
rect 510068 6384 510120 6390
rect 510068 6326 510120 6332
rect 508872 4412 508924 4418
rect 508872 4354 508924 4360
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 4354
rect 510080 480 510108 6326
rect 511276 480 511304 11999
rect 517886 11928 517942 11937
rect 517886 11863 517942 11872
rect 514758 11792 514814 11801
rect 514758 11727 514814 11736
rect 513564 8900 513616 8906
rect 513564 8842 513616 8848
rect 512460 4480 512512 4486
rect 512460 4422 512512 4428
rect 512472 480 512500 4422
rect 513576 480 513604 8842
rect 514772 480 514800 11727
rect 517152 6316 517204 6322
rect 517152 6258 517204 6264
rect 515956 4548 516008 4554
rect 515956 4490 516008 4496
rect 515968 480 515996 4490
rect 517164 480 517192 6258
rect 517900 490 517928 11863
rect 521842 11656 521898 11665
rect 521842 11591 521898 11600
rect 520740 9648 520792 9654
rect 520740 9590 520792 9596
rect 519544 4616 519596 4622
rect 519544 4558 519596 4564
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 4558
rect 520752 480 520780 9590
rect 521856 480 521884 11591
rect 524236 6248 524288 6254
rect 524236 6190 524288 6196
rect 523040 4752 523092 4758
rect 523040 4694 523092 4700
rect 523052 480 523080 4694
rect 524248 480 524276 6190
rect 525444 480 525472 13534
rect 532056 13524 532108 13530
rect 532056 13466 532108 13472
rect 528560 13456 528612 13462
rect 528560 13398 528612 13404
rect 527824 9580 527876 9586
rect 527824 9522 527876 9528
rect 526628 4684 526680 4690
rect 526628 4626 526680 4632
rect 526640 480 526668 4626
rect 527836 480 527864 9522
rect 528572 490 528600 13398
rect 531318 6624 531374 6633
rect 531318 6559 531374 6568
rect 530124 5500 530176 5506
rect 530124 5442 530176 5448
rect 528848 598 529060 626
rect 528848 490 528876 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 5442
rect 531332 480 531360 6559
rect 532068 490 532096 13466
rect 539598 13424 539654 13433
rect 536104 13388 536156 13394
rect 539598 13359 539654 13368
rect 536104 13330 536156 13336
rect 534908 9512 534960 9518
rect 534908 9454 534960 9460
rect 533712 5432 533764 5438
rect 533712 5374 533764 5380
rect 532344 598 532556 626
rect 532344 490 532372 598
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 462 532372 490
rect 532528 480 532556 598
rect 533724 480 533752 5374
rect 534920 480 534948 9454
rect 536116 480 536144 13330
rect 538404 9444 538456 9450
rect 538404 9386 538456 9392
rect 537208 5364 537260 5370
rect 537208 5306 537260 5312
rect 537220 480 537248 5306
rect 538416 480 538444 9386
rect 539612 480 539640 13359
rect 546684 13320 546736 13326
rect 542726 13288 542782 13297
rect 546684 13262 546736 13268
rect 542726 13223 542782 13232
rect 541992 9376 542044 9382
rect 541992 9318 542044 9324
rect 540796 5296 540848 5302
rect 540796 5238 540848 5244
rect 540808 480 540836 5238
rect 542004 480 542032 9318
rect 542740 490 542768 13223
rect 545486 6488 545542 6497
rect 545486 6423 545542 6432
rect 544384 5228 544436 5234
rect 544384 5170 544436 5176
rect 543016 598 543228 626
rect 543016 490 543044 598
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 5170
rect 545500 480 545528 6423
rect 546696 480 546724 13262
rect 553768 13252 553820 13258
rect 553768 13194 553820 13200
rect 550270 13152 550326 13161
rect 550270 13087 550326 13096
rect 549076 9308 549128 9314
rect 549076 9250 549128 9256
rect 547880 5160 547932 5166
rect 547880 5102 547932 5108
rect 547892 480 547920 5102
rect 549088 480 549116 9250
rect 550284 480 550312 13087
rect 552662 8936 552718 8945
rect 552662 8871 552718 8880
rect 551468 5092 551520 5098
rect 551468 5034 551520 5040
rect 551480 480 551508 5034
rect 552676 480 552704 8871
rect 553780 480 553808 13194
rect 556158 6352 556214 6361
rect 556158 6287 556214 6296
rect 554962 5128 555018 5137
rect 554962 5063 555018 5072
rect 554976 480 555004 5063
rect 556172 480 556200 6287
rect 556908 490 556936 14486
rect 559288 14476 559340 14482
rect 559288 14418 559340 14424
rect 558550 4992 558606 5001
rect 558550 4927 558606 4936
rect 557184 598 557396 626
rect 557184 490 557212 598
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 462 557212 490
rect 557368 480 557396 598
rect 558564 480 558592 4927
rect 559300 490 559328 14418
rect 559576 598 559788 626
rect 559576 490 559604 598
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 462 559604 490
rect 559760 480 559788 598
rect 560404 490 560432 14719
rect 571522 14648 571578 14657
rect 571522 14583 571578 14592
rect 564438 13016 564494 13025
rect 564438 12951 564494 12960
rect 563244 9240 563296 9246
rect 563244 9182 563296 9188
rect 562048 5024 562100 5030
rect 562048 4966 562100 4972
rect 560680 598 560892 626
rect 560680 490 560708 598
rect 559718 -960 559830 480
rect 560404 462 560708 490
rect 560864 480 560892 598
rect 562060 480 562088 4966
rect 563256 480 563284 9182
rect 564452 480 564480 12951
rect 566832 9172 566884 9178
rect 566832 9114 566884 9120
rect 565636 4956 565688 4962
rect 565636 4898 565688 4904
rect 565648 480 565676 4898
rect 566844 480 566872 9114
rect 570326 6216 570382 6225
rect 570326 6151 570382 6160
rect 569132 4888 569184 4894
rect 569132 4830 569184 4836
rect 568028 3664 568080 3670
rect 568028 3606 568080 3612
rect 568040 480 568068 3606
rect 569144 480 569172 4830
rect 570340 480 570368 6151
rect 571536 480 571564 14583
rect 575110 14512 575166 14521
rect 575110 14447 575166 14456
rect 573916 9036 573968 9042
rect 573916 8978 573968 8984
rect 572718 4856 572774 4865
rect 572718 4791 572774 4800
rect 572732 480 572760 4791
rect 573928 480 573956 8978
rect 575124 480 575152 14447
rect 576952 13184 577004 13190
rect 576952 13126 577004 13132
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 576320 480 576348 4762
rect 576964 490 576992 13126
rect 581736 13116 581788 13122
rect 581736 13058 581788 13064
rect 581000 9104 581052 9110
rect 581000 9046 581052 9052
rect 578608 8968 578660 8974
rect 578608 8910 578660 8916
rect 577240 598 577452 626
rect 577240 490 577268 598
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 462 577268 490
rect 577424 480 577452 598
rect 578620 480 578648 8910
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 9046
rect 581748 490 581776 13058
rect 583392 3120 583444 3126
rect 583392 3062 583444 3068
rect 582024 598 582236 626
rect 582024 490 582052 598
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 462 582052 490
rect 582208 480 582236 598
rect 583404 480 583432 3062
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2870 658144 2926 658200
rect 3514 671200 3570 671256
rect 32034 645924 32090 645960
rect 32034 645904 32036 645924
rect 32036 645904 32088 645924
rect 32088 645904 32090 645924
rect 3698 639920 3754 639976
rect 3422 634888 3478 634944
rect 3238 632032 3294 632088
rect 3422 619112 3478 619168
rect 3422 607144 3478 607200
rect 3422 606056 3478 606112
rect 3422 593000 3478 593056
rect 3422 579944 3478 580000
rect 3330 553832 3386 553888
rect 3330 540776 3386 540832
rect 3330 527856 3386 527912
rect 3330 514800 3386 514856
rect 2870 501744 2926 501800
rect 3054 475632 3110 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 2870 410488 2926 410544
rect 3330 319232 3386 319288
rect 3698 566888 3754 566944
rect 3606 488688 3662 488744
rect 3514 436600 3570 436656
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 371320 3570 371376
rect 3606 358400 3662 358456
rect 3974 345344 4030 345400
rect 2962 306212 2964 306232
rect 2964 306212 3016 306232
rect 3016 306212 3018 306232
rect 2962 306176 3018 306212
rect 2778 293120 2834 293176
rect 2778 267180 2780 267200
rect 2780 267180 2832 267200
rect 2832 267180 2834 267200
rect 2778 267144 2834 267180
rect 3146 254088 3202 254144
rect 2778 241068 2780 241088
rect 2780 241068 2832 241088
rect 2832 241068 2834 241088
rect 2778 241032 2834 241068
rect 2778 214956 2780 214976
rect 2780 214956 2832 214976
rect 2832 214956 2834 214976
rect 2778 214920 2834 214956
rect 3514 311888 3570 311944
rect 3330 201864 3386 201920
rect 3146 149776 3202 149832
rect 2778 123664 2834 123720
rect 2778 110608 2834 110664
rect 2778 84632 2834 84688
rect 2778 71612 2780 71632
rect 2780 71612 2832 71632
rect 2832 71612 2834 71632
rect 2778 71576 2834 71612
rect 2778 45500 2780 45520
rect 2780 45500 2832 45520
rect 2832 45500 2834 45520
rect 2778 45464 2834 45500
rect 4066 188808 4122 188864
rect 3974 162832 4030 162888
rect 3882 136720 3938 136776
rect 90822 639940 90878 639976
rect 90822 639920 90824 639940
rect 90824 639920 90876 639940
rect 90876 639920 90878 639940
rect 96342 639940 96398 639976
rect 96342 639920 96344 639940
rect 96344 639920 96396 639940
rect 96396 639920 96398 639940
rect 90822 634924 90824 634944
rect 90824 634924 90876 634944
rect 90876 634924 90878 634944
rect 90822 634888 90878 634924
rect 96986 634924 96988 634944
rect 96988 634924 97040 634944
rect 97040 634924 97042 634944
rect 96986 634888 97042 634924
rect 97906 633256 97962 633312
rect 31758 622104 31814 622160
rect 31758 619676 31814 619712
rect 31758 619656 31760 619676
rect 31760 619656 31812 619676
rect 31812 619656 31814 619676
rect 120262 634908 120318 634944
rect 120262 634888 120264 634908
rect 120264 634888 120316 634908
rect 120316 634888 120318 634908
rect 99746 633256 99802 633312
rect 31758 602248 31814 602304
rect 98458 601976 98514 602032
rect 126794 634908 126850 634944
rect 126794 634888 126796 634908
rect 126796 634888 126848 634908
rect 126848 634888 126850 634908
rect 126886 632304 126942 632360
rect 98642 601568 98698 601624
rect 31850 578312 31906 578368
rect 118606 590688 118662 590744
rect 3790 97552 3846 97608
rect 3698 58520 3754 58576
rect 68006 312296 68062 312352
rect 50986 312160 51042 312216
rect 43994 312024 44050 312080
rect 121366 576816 121422 576872
rect 139490 576816 139546 576872
rect 153106 639784 153162 639840
rect 160006 640056 160062 640112
rect 159546 590688 159602 590744
rect 160098 607164 160154 607200
rect 160098 607144 160100 607164
rect 160100 607144 160152 607164
rect 160152 607144 160154 607164
rect 160926 607164 160982 607200
rect 160926 607144 160928 607164
rect 160928 607144 160980 607164
rect 160980 607144 160982 607164
rect 182914 639240 182970 639296
rect 184018 639104 184074 639160
rect 182546 638988 182602 639024
rect 182546 638968 182548 638988
rect 182548 638968 182600 638988
rect 182600 638968 182602 638988
rect 252466 669296 252522 669352
rect 194690 639240 194746 639296
rect 194598 639104 194654 639160
rect 176198 635160 176254 635216
rect 176566 634888 176622 634944
rect 184202 634888 184258 634944
rect 184754 634888 184810 634944
rect 184202 632440 184258 632496
rect 184754 632440 184810 632496
rect 197450 638968 197506 639024
rect 189262 634908 189318 634944
rect 189262 634888 189264 634908
rect 189264 634888 189316 634908
rect 189316 634888 189318 634908
rect 191562 634908 191618 634944
rect 191562 634888 191564 634908
rect 191564 634888 191616 634908
rect 191616 634888 191618 634908
rect 205362 638968 205418 639024
rect 233882 639240 233938 639296
rect 218886 638968 218942 639024
rect 201866 634888 201922 634944
rect 196162 633936 196218 633992
rect 196346 633936 196402 633992
rect 196346 633664 196402 633720
rect 196254 633528 196310 633584
rect 189814 632460 189870 632496
rect 189814 632440 189816 632460
rect 189816 632440 189868 632460
rect 189868 632440 189870 632460
rect 191562 632304 191618 632360
rect 191562 631388 191564 631408
rect 191564 631388 191616 631408
rect 191616 631388 191618 631408
rect 191562 631352 191618 631388
rect 192942 631352 192998 631408
rect 210238 632168 210294 632224
rect 215390 631216 215446 631272
rect 221094 631216 221150 631272
rect 204902 607144 204958 607200
rect 364338 639104 364394 639160
rect 404266 632032 404322 632088
rect 463330 692844 463386 692880
rect 463330 692824 463332 692844
rect 463332 692824 463384 692844
rect 463384 692824 463386 692844
rect 465538 692824 465594 692880
rect 580170 697176 580226 697232
rect 580354 683848 580410 683904
rect 580262 670656 580318 670712
rect 459558 644544 459614 644600
rect 468666 644544 468722 644600
rect 469034 644544 469090 644600
rect 471886 644544 471942 644600
rect 415306 640192 415362 640248
rect 423586 640192 423642 640248
rect 424230 640192 424286 640248
rect 429198 640192 429254 640248
rect 414662 631216 414718 631272
rect 422666 631216 422722 631272
rect 423402 631216 423458 631272
rect 436742 631216 436798 631272
rect 391846 559408 391902 559464
rect 391386 543496 391442 543552
rect 427818 551520 427874 551576
rect 496082 631080 496138 631136
rect 506662 631080 506718 631136
rect 579618 644000 579674 644056
rect 579802 630808 579858 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 579986 577632 580042 577688
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 579986 484608 580042 484664
rect 580170 471416 580226 471472
rect 579618 458088 579674 458144
rect 579894 431568 579950 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 580354 564304 580410 564360
rect 303250 312160 303306 312216
rect 303066 312024 303122 312080
rect 300950 311888 301006 311944
rect 29550 310120 29606 310176
rect 34334 309984 34390 310040
rect 36726 309984 36782 310040
rect 3606 32408 3662 32464
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 79782 3576 79838 3632
rect 84014 3440 84070 3496
rect 84106 3304 84162 3360
rect 110510 3576 110566 3632
rect 117594 3440 117650 3496
rect 118790 3304 118846 3360
rect 131026 3712 131082 3768
rect 133786 3576 133842 3632
rect 135166 3440 135222 3496
rect 139306 5072 139362 5128
rect 140686 3304 140742 3360
rect 148966 6568 149022 6624
rect 150254 6432 150310 6488
rect 153014 6296 153070 6352
rect 151726 4936 151782 4992
rect 154486 4800 154542 4856
rect 157246 6160 157302 6216
rect 176566 9288 176622 9344
rect 179234 9152 179290 9208
rect 180706 9016 180762 9072
rect 195886 5208 195942 5264
rect 216862 3712 216918 3768
rect 220634 10648 220690 10704
rect 222014 10512 222070 10568
rect 223394 10376 223450 10432
rect 224682 10240 224738 10296
rect 223946 3576 224002 3632
rect 227534 3440 227590 3496
rect 235814 5072 235870 5128
rect 238758 30912 238814 30968
rect 238666 7928 238722 7984
rect 240046 7792 240102 7848
rect 241426 7656 241482 7712
rect 238114 3304 238170 3360
rect 249062 31184 249118 31240
rect 246946 7520 247002 7576
rect 252466 31048 252522 31104
rect 251086 3440 251142 3496
rect 254674 6568 254730 6624
rect 253846 3304 253902 3360
rect 258262 6432 258318 6488
rect 260654 4936 260710 4992
rect 265346 6296 265402 6352
rect 268934 12008 268990 12064
rect 270222 11736 270278 11792
rect 267738 4800 267794 4856
rect 273074 11872 273130 11928
rect 272430 6160 272486 6216
rect 274362 11600 274418 11656
rect 278594 6568 278650 6624
rect 282642 13368 282698 13424
rect 284114 13232 284170 13288
rect 285494 6432 285550 6488
rect 288162 13096 288218 13152
rect 288254 8880 288310 8936
rect 289726 5072 289782 5128
rect 291014 6296 291070 6352
rect 292486 14728 292542 14784
rect 293682 12960 293738 13016
rect 291106 4936 291162 4992
rect 296534 6160 296590 6216
rect 297914 14592 297970 14648
rect 299202 14456 299258 14512
rect 298006 4800 298062 4856
rect 302974 309440 303030 309496
rect 304446 312296 304502 312352
rect 580170 312024 580226 312080
rect 315302 309304 315358 309360
rect 302146 31320 302202 31376
rect 315026 9288 315082 9344
rect 580262 309168 580318 309224
rect 580170 298696 580226 298752
rect 579986 272176 580042 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 205672 580226 205728
rect 579618 165824 579674 165880
rect 579802 152632 579858 152688
rect 579710 125976 579766 126032
rect 579618 86128 579674 86184
rect 580170 72936 580226 72992
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 322202 31320 322258 31376
rect 318522 9152 318578 9208
rect 322110 9016 322166 9072
rect 323582 31184 323638 31240
rect 323582 3576 323638 3632
rect 348422 3168 348478 3224
rect 351826 3168 351882 3224
rect 356334 5208 356390 5264
rect 382922 31048 382978 31104
rect 380162 30912 380218 30968
rect 580906 219000 580962 219056
rect 580814 192480 580870 192536
rect 580722 179152 580778 179208
rect 580630 139304 580686 139360
rect 580538 112784 580594 112840
rect 580446 99456 580502 99512
rect 580354 59608 580410 59664
rect 580262 19760 580318 19816
rect 407210 10648 407266 10704
rect 410798 10512 410854 10568
rect 414294 10376 414350 10432
rect 417422 10240 417478 10296
rect 445022 7928 445078 7984
rect 448610 7792 448666 7848
rect 452106 7656 452162 7712
rect 462778 7520 462834 7576
rect 560390 14728 560446 14784
rect 468666 3576 468722 3632
rect 472254 3440 472310 3496
rect 479338 3304 479394 3360
rect 511262 12008 511318 12064
rect 517886 11872 517942 11928
rect 514758 11736 514814 11792
rect 521842 11600 521898 11656
rect 531318 6568 531374 6624
rect 539598 13368 539654 13424
rect 542726 13232 542782 13288
rect 545486 6432 545542 6488
rect 550270 13096 550326 13152
rect 552662 8880 552718 8936
rect 556158 6296 556214 6352
rect 554962 5072 555018 5128
rect 558550 4936 558606 4992
rect 571522 14592 571578 14648
rect 564438 12960 564494 13016
rect 570326 6160 570382 6216
rect 575110 14456 575166 14512
rect 572718 4800 572774 4856
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect 463325 692882 463391 692885
rect 465533 692882 465599 692885
rect 463325 692880 465599 692882
rect 463325 692824 463330 692880
rect 463386 692824 465538 692880
rect 465594 692824 465599 692880
rect 463325 692822 465599 692824
rect 463325 692819 463391 692822
rect 465533 692819 465599 692822
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580349 683906 580415 683909
rect 583520 683906 584960 683996
rect 580349 683904 584960 683906
rect 580349 683848 580354 683904
rect 580410 683848 584960 683904
rect 580349 683846 584960 683848
rect 580349 683843 580415 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect 252461 669354 252527 669357
rect 252461 669352 528570 669354
rect 252461 669296 252466 669352
rect 252522 669296 528570 669352
rect 252461 669294 528570 669296
rect 252461 669291 252527 669294
rect 528510 668916 528570 669294
rect -960 658202 480 658292
rect 2865 658202 2931 658205
rect -960 658200 2931 658202
rect -960 658144 2870 658200
rect 2926 658144 2931 658200
rect -960 658142 2931 658144
rect -960 658052 480 658142
rect 2865 658139 2931 658142
rect 583520 657236 584960 657476
rect 32078 645965 32138 646340
rect 32029 645960 32138 645965
rect 32029 645904 32034 645960
rect 32090 645904 32138 645960
rect 32029 645902 32138 645904
rect 32029 645899 32095 645902
rect -960 644996 480 645236
rect 459553 644602 459619 644605
rect 468661 644602 468727 644605
rect 459553 644600 468727 644602
rect 459553 644544 459558 644600
rect 459614 644544 468666 644600
rect 468722 644544 468727 644600
rect 459553 644542 468727 644544
rect 459553 644539 459619 644542
rect 468661 644539 468727 644542
rect 469029 644602 469095 644605
rect 471881 644602 471947 644605
rect 469029 644600 471947 644602
rect 469029 644544 469034 644600
rect 469090 644544 471886 644600
rect 471942 644544 471947 644600
rect 469029 644542 471947 644544
rect 469029 644539 469095 644542
rect 471881 644539 471947 644542
rect 579613 644058 579679 644061
rect 583520 644058 584960 644148
rect 579613 644056 584960 644058
rect 579613 644000 579618 644056
rect 579674 644000 584960 644056
rect 579613 643998 584960 644000
rect 579613 643995 579679 643998
rect 583520 643908 584960 643998
rect 415301 640250 415367 640253
rect 423581 640250 423647 640253
rect 415301 640248 423647 640250
rect 415301 640192 415306 640248
rect 415362 640192 423586 640248
rect 423642 640192 423647 640248
rect 415301 640190 423647 640192
rect 415301 640187 415367 640190
rect 423581 640187 423647 640190
rect 424225 640250 424291 640253
rect 429193 640250 429259 640253
rect 424225 640248 429259 640250
rect 424225 640192 424230 640248
rect 424286 640192 429198 640248
rect 429254 640192 429259 640248
rect 424225 640190 429259 640192
rect 424225 640187 424291 640190
rect 429193 640187 429259 640190
rect 160001 640114 160067 640117
rect 160001 640112 183202 640114
rect 160001 640056 160006 640112
rect 160062 640056 183202 640112
rect 160001 640054 183202 640056
rect 160001 640051 160067 640054
rect 3693 639978 3759 639981
rect 90817 639978 90883 639981
rect 3693 639976 90883 639978
rect 3693 639920 3698 639976
rect 3754 639920 90822 639976
rect 90878 639920 90883 639976
rect 3693 639918 90883 639920
rect 3693 639915 3759 639918
rect 90817 639915 90883 639918
rect 96337 639978 96403 639981
rect 96337 639976 182834 639978
rect 96337 639920 96342 639976
rect 96398 639920 182834 639976
rect 96337 639918 182834 639920
rect 96337 639915 96403 639918
rect 153101 639842 153167 639845
rect 153101 639840 181546 639842
rect 153101 639784 153106 639840
rect 153162 639784 181546 639840
rect 153101 639782 181546 639784
rect 153101 639779 153167 639782
rect 181486 639298 181546 639782
rect 182774 639298 182834 639918
rect 182909 639298 182975 639301
rect 181486 639268 182068 639298
rect 182774 639296 182975 639298
rect 181516 639238 182098 639268
rect 182774 639240 182914 639296
rect 182970 639240 182975 639296
rect 182774 639238 182975 639240
rect 182038 639026 182098 639238
rect 182909 639235 182975 639238
rect 183142 639162 183202 640054
rect 194685 639298 194751 639301
rect 233877 639298 233943 639301
rect 194685 639296 233943 639298
rect 194685 639240 194690 639296
rect 194746 639240 233882 639296
rect 233938 639240 233943 639296
rect 194685 639238 233943 639240
rect 194685 639235 194751 639238
rect 233877 639235 233943 639238
rect 184013 639162 184079 639165
rect 183142 639160 184079 639162
rect 183142 639132 184018 639160
rect 183172 639104 184018 639132
rect 184074 639104 184079 639160
rect 183172 639102 184079 639104
rect 184013 639099 184079 639102
rect 194593 639162 194659 639165
rect 364333 639162 364399 639165
rect 194593 639160 364399 639162
rect 194593 639104 194598 639160
rect 194654 639104 364338 639160
rect 364394 639104 364399 639160
rect 194593 639102 364399 639104
rect 194593 639099 194659 639102
rect 364333 639099 364399 639102
rect 182541 639026 182607 639029
rect 182038 639024 182607 639026
rect 182038 638996 182546 639024
rect 182068 638968 182546 638996
rect 182602 638968 182607 639024
rect 182068 638966 182607 638968
rect 182541 638963 182607 638966
rect 197445 639026 197511 639029
rect 205357 639026 205423 639029
rect 218881 639026 218947 639029
rect 197445 639024 218947 639026
rect 197445 638968 197450 639024
rect 197506 638968 205362 639024
rect 205418 638968 218886 639024
rect 218942 638968 218947 639024
rect 197445 638966 218947 638968
rect 197445 638963 197511 638966
rect 205357 638963 205423 638966
rect 218881 638963 218947 638966
rect 176193 635218 176259 635221
rect 161430 635216 176259 635218
rect 161430 635160 176198 635216
rect 176254 635160 176259 635216
rect 161430 635158 176259 635160
rect 3417 634946 3483 634949
rect 90817 634946 90883 634949
rect 3417 634944 90883 634946
rect 3417 634888 3422 634944
rect 3478 634888 90822 634944
rect 90878 634888 90883 634944
rect 3417 634886 90883 634888
rect 3417 634883 3483 634886
rect 90817 634883 90883 634886
rect 96981 634946 97047 634949
rect 120257 634946 120323 634949
rect 96981 634944 120323 634946
rect 96981 634888 96986 634944
rect 97042 634888 120262 634944
rect 120318 634888 120323 634944
rect 96981 634886 120323 634888
rect 96981 634883 97047 634886
rect 120257 634883 120323 634886
rect 126789 634946 126855 634949
rect 161430 634946 161490 635158
rect 176193 635155 176259 635158
rect 126789 634944 161490 634946
rect 126789 634888 126794 634944
rect 126850 634888 161490 634944
rect 126789 634886 161490 634888
rect 176561 634946 176627 634949
rect 184197 634946 184263 634949
rect 176561 634944 184263 634946
rect 176561 634888 176566 634944
rect 176622 634888 184202 634944
rect 184258 634888 184263 634944
rect 176561 634886 184263 634888
rect 126789 634883 126855 634886
rect 176561 634883 176627 634886
rect 184197 634883 184263 634886
rect 184749 634946 184815 634949
rect 189257 634946 189323 634949
rect 184749 634944 189323 634946
rect 184749 634888 184754 634944
rect 184810 634888 189262 634944
rect 189318 634888 189323 634944
rect 184749 634886 189323 634888
rect 184749 634883 184815 634886
rect 189257 634883 189323 634886
rect 191557 634946 191623 634949
rect 201861 634946 201927 634949
rect 191557 634944 201927 634946
rect 191557 634888 191562 634944
rect 191618 634888 201866 634944
rect 201922 634888 201927 634944
rect 191557 634886 201927 634888
rect 191557 634883 191623 634886
rect 201861 634883 201927 634886
rect 196157 633994 196223 633997
rect 196341 633994 196407 633997
rect 196157 633992 196266 633994
rect 196157 633936 196162 633992
rect 196218 633936 196266 633992
rect 196157 633931 196266 633936
rect 196341 633992 196450 633994
rect 196341 633936 196346 633992
rect 196402 633936 196450 633992
rect 196341 633931 196450 633936
rect 196206 633589 196266 633931
rect 196390 633725 196450 633931
rect 196341 633720 196450 633725
rect 196341 633664 196346 633720
rect 196402 633664 196450 633720
rect 196341 633662 196450 633664
rect 196341 633659 196407 633662
rect 196206 633584 196315 633589
rect 196206 633528 196254 633584
rect 196310 633528 196315 633584
rect 196206 633526 196315 633528
rect 196249 633523 196315 633526
rect 97901 633314 97967 633317
rect 99741 633314 99807 633317
rect 97901 633312 99807 633314
rect 97901 633256 97906 633312
rect 97962 633256 99746 633312
rect 99802 633256 99807 633312
rect 97901 633254 99807 633256
rect 97901 633251 97967 633254
rect 99741 633251 99807 633254
rect 184197 632498 184263 632501
rect 180750 632496 184263 632498
rect 180750 632440 184202 632496
rect 184258 632440 184263 632496
rect 180750 632438 184263 632440
rect 126881 632362 126947 632365
rect 180750 632362 180810 632438
rect 184197 632435 184263 632438
rect 184749 632498 184815 632501
rect 189809 632498 189875 632501
rect 184749 632496 189875 632498
rect 184749 632440 184754 632496
rect 184810 632440 189814 632496
rect 189870 632440 189875 632496
rect 184749 632438 189875 632440
rect 184749 632435 184815 632438
rect 189809 632435 189875 632438
rect 126881 632360 180810 632362
rect 126881 632304 126886 632360
rect 126942 632304 180810 632360
rect 126881 632302 180810 632304
rect 191557 632362 191623 632365
rect 191557 632360 195990 632362
rect 191557 632304 191562 632360
rect 191618 632304 195990 632360
rect 191557 632302 195990 632304
rect 126881 632299 126947 632302
rect 191557 632299 191623 632302
rect 195930 632226 195990 632302
rect 210233 632226 210299 632229
rect 195930 632224 210299 632226
rect -960 632090 480 632180
rect 195930 632168 210238 632224
rect 210294 632168 210299 632224
rect 195930 632166 210299 632168
rect 210233 632163 210299 632166
rect 3233 632090 3299 632093
rect -960 632088 3299 632090
rect -960 632032 3238 632088
rect 3294 632032 3299 632088
rect -960 632030 3299 632032
rect -960 631940 480 632030
rect 3233 632027 3299 632030
rect 404261 632090 404327 632093
rect 404261 632088 406364 632090
rect 404261 632032 404266 632088
rect 404322 632032 406364 632088
rect 404261 632030 406364 632032
rect 404261 632027 404327 632030
rect 191557 631410 191623 631413
rect 192937 631410 193003 631413
rect 191557 631408 193003 631410
rect 191557 631352 191562 631408
rect 191618 631352 192942 631408
rect 192998 631352 193003 631408
rect 191557 631350 193003 631352
rect 191557 631347 191623 631350
rect 192937 631347 193003 631350
rect 215385 631274 215451 631277
rect 221089 631274 221155 631277
rect 215385 631272 221155 631274
rect 215385 631216 215390 631272
rect 215446 631216 221094 631272
rect 221150 631216 221155 631272
rect 215385 631214 221155 631216
rect 215385 631211 215451 631214
rect 221089 631211 221155 631214
rect 414657 631274 414723 631277
rect 422661 631274 422727 631277
rect 414657 631272 422727 631274
rect 414657 631216 414662 631272
rect 414718 631216 422666 631272
rect 422722 631216 422727 631272
rect 414657 631214 422727 631216
rect 414657 631211 414723 631214
rect 422661 631211 422727 631214
rect 423397 631274 423463 631277
rect 436737 631274 436803 631277
rect 423397 631272 436803 631274
rect 423397 631216 423402 631272
rect 423458 631216 436742 631272
rect 436798 631216 436803 631272
rect 423397 631214 436803 631216
rect 423397 631211 423463 631214
rect 436737 631211 436803 631214
rect 496077 631138 496143 631141
rect 506657 631138 506723 631141
rect 496077 631136 506723 631138
rect 496077 631080 496082 631136
rect 496138 631080 506662 631136
rect 506718 631080 506723 631136
rect 496077 631078 506723 631080
rect 496077 631075 496143 631078
rect 506657 631075 506723 631078
rect 579797 630866 579863 630869
rect 583520 630866 584960 630956
rect 579797 630864 584960 630866
rect 579797 630808 579802 630864
rect 579858 630808 584960 630864
rect 579797 630806 584960 630808
rect 579797 630803 579863 630806
rect 583520 630716 584960 630806
rect 31753 622162 31819 622165
rect 31753 622160 32108 622162
rect 31753 622104 31758 622160
rect 31814 622104 32108 622160
rect 31753 622102 32108 622104
rect 31753 622099 31819 622102
rect 31753 619714 31819 619717
rect 31753 619712 32108 619714
rect 31753 619656 31758 619712
rect 31814 619656 32108 619712
rect 31753 619654 32108 619656
rect 31753 619651 31819 619654
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 3417 607202 3483 607205
rect 160093 607202 160159 607205
rect 3417 607200 160159 607202
rect 3417 607144 3422 607200
rect 3478 607144 160098 607200
rect 160154 607144 160159 607200
rect 3417 607142 160159 607144
rect 3417 607139 3483 607142
rect 160093 607139 160159 607142
rect 160921 607202 160987 607205
rect 204897 607202 204963 607205
rect 160921 607200 204963 607202
rect 160921 607144 160926 607200
rect 160982 607144 204902 607200
rect 204958 607144 204963 607200
rect 160921 607142 204963 607144
rect 160921 607139 160987 607142
rect 204897 607139 204963 607142
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect 31753 602306 31819 602309
rect 31753 602304 32108 602306
rect 31753 602248 31758 602304
rect 31814 602248 32108 602304
rect 31753 602246 32108 602248
rect 31753 602243 31819 602246
rect 98453 602034 98519 602037
rect 98453 602032 98562 602034
rect 98453 601976 98458 602032
rect 98514 601976 98562 602032
rect 98453 601971 98562 601976
rect 98502 601626 98562 601971
rect 98637 601626 98703 601629
rect 98502 601624 98703 601626
rect 98502 601568 98642 601624
rect 98698 601568 98703 601624
rect 98502 601566 98703 601568
rect 98637 601563 98703 601566
rect -960 593058 480 593148
rect 3417 593058 3483 593061
rect -960 593056 3483 593058
rect -960 593000 3422 593056
rect 3478 593000 3483 593056
rect -960 592998 3483 593000
rect -960 592908 480 592998
rect 3417 592995 3483 592998
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect 118601 590746 118667 590749
rect 159541 590746 159607 590749
rect 118601 590744 159607 590746
rect 118601 590688 118606 590744
rect 118662 590688 159546 590744
rect 159602 590688 159607 590744
rect 118601 590686 159607 590688
rect 118601 590683 118667 590686
rect 159541 590683 159607 590686
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 31845 578370 31911 578373
rect 31845 578368 32108 578370
rect 31845 578312 31850 578368
rect 31906 578312 32108 578368
rect 31845 578310 32108 578312
rect 31845 578307 31911 578310
rect 579981 577690 580047 577693
rect 583520 577690 584960 577780
rect 579981 577688 584960 577690
rect 579981 577632 579986 577688
rect 580042 577632 584960 577688
rect 579981 577630 584960 577632
rect 579981 577627 580047 577630
rect 583520 577540 584960 577630
rect 121361 576874 121427 576877
rect 139485 576874 139551 576877
rect 121361 576872 139551 576874
rect 121361 576816 121366 576872
rect 121422 576816 139490 576872
rect 139546 576816 139551 576872
rect 121361 576814 139551 576816
rect 121361 576811 121427 576814
rect 139485 576811 139551 576814
rect -960 566946 480 567036
rect 3693 566946 3759 566949
rect -960 566944 3759 566946
rect -960 566888 3698 566944
rect 3754 566888 3759 566944
rect -960 566886 3759 566888
rect -960 566796 480 566886
rect 3693 566883 3759 566886
rect 580349 564362 580415 564365
rect 583520 564362 584960 564452
rect 580349 564360 584960 564362
rect 580349 564304 580354 564360
rect 580410 564304 584960 564360
rect 580349 564302 584960 564304
rect 580349 564299 580415 564302
rect 583520 564212 584960 564302
rect 391841 559466 391907 559469
rect 391841 559464 394036 559466
rect 391841 559408 391846 559464
rect 391902 559408 394036 559464
rect 391841 559406 394036 559408
rect 391841 559403 391907 559406
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 427813 551578 427879 551581
rect 425868 551576 427879 551578
rect 425868 551520 427818 551576
rect 427874 551520 427879 551576
rect 425868 551518 427879 551520
rect 427813 551515 427879 551518
rect 583520 551020 584960 551260
rect 391381 543554 391447 543557
rect 391381 543552 394036 543554
rect 391381 543496 391386 543552
rect 391442 543496 394036 543552
rect 391381 543494 394036 543496
rect 391381 543491 391447 543494
rect -960 540834 480 540924
rect 3325 540834 3391 540837
rect -960 540832 3391 540834
rect -960 540776 3330 540832
rect 3386 540776 3391 540832
rect -960 540774 3391 540776
rect -960 540684 480 540774
rect 3325 540771 3391 540774
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2865 501802 2931 501805
rect -960 501800 2931 501802
rect -960 501744 2870 501800
rect 2926 501744 2931 501800
rect -960 501742 2931 501744
rect -960 501652 480 501742
rect 2865 501739 2931 501742
rect 583520 497844 584960 498084
rect -960 488746 480 488836
rect 3601 488746 3667 488749
rect -960 488744 3667 488746
rect -960 488688 3606 488744
rect 3662 488688 3667 488744
rect -960 488686 3667 488688
rect -960 488596 480 488686
rect 3601 488683 3667 488686
rect 579981 484666 580047 484669
rect 583520 484666 584960 484756
rect 579981 484664 584960 484666
rect 579981 484608 579986 484664
rect 580042 484608 584960 484664
rect 579981 484606 584960 484608
rect 579981 484603 580047 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 579613 458146 579679 458149
rect 583520 458146 584960 458236
rect 579613 458144 584960 458146
rect 579613 458088 579618 458144
rect 579674 458088 584960 458144
rect 579613 458086 584960 458088
rect 579613 458083 579679 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436658 480 436748
rect 3509 436658 3575 436661
rect -960 436656 3575 436658
rect -960 436600 3514 436656
rect 3570 436600 3575 436656
rect -960 436598 3575 436600
rect -960 436508 480 436598
rect 3509 436595 3575 436598
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3969 345402 4035 345405
rect -960 345400 4035 345402
rect -960 345344 3974 345400
rect 4030 345344 4035 345400
rect -960 345342 4035 345344
rect -960 345252 480 345342
rect 3969 345339 4035 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 68001 312354 68067 312357
rect 304441 312354 304507 312357
rect 68001 312352 304507 312354
rect 68001 312296 68006 312352
rect 68062 312296 304446 312352
rect 304502 312296 304507 312352
rect 68001 312294 304507 312296
rect 68001 312291 68067 312294
rect 304441 312291 304507 312294
rect 50981 312218 51047 312221
rect 303245 312218 303311 312221
rect 50981 312216 303311 312218
rect 50981 312160 50986 312216
rect 51042 312160 303250 312216
rect 303306 312160 303311 312216
rect 50981 312158 303311 312160
rect 50981 312155 51047 312158
rect 303245 312155 303311 312158
rect 43989 312082 44055 312085
rect 303061 312082 303127 312085
rect 43989 312080 303127 312082
rect 43989 312024 43994 312080
rect 44050 312024 303066 312080
rect 303122 312024 303127 312080
rect 43989 312022 303127 312024
rect 43989 312019 44055 312022
rect 303061 312019 303127 312022
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 3509 311946 3575 311949
rect 300945 311946 301011 311949
rect 3509 311944 301011 311946
rect 3509 311888 3514 311944
rect 3570 311888 300950 311944
rect 301006 311888 301011 311944
rect 583520 311932 584960 312022
rect 3509 311886 301011 311888
rect 3509 311883 3575 311886
rect 300945 311883 301011 311886
rect 29545 310178 29611 310181
rect 29545 310176 36554 310178
rect 29545 310120 29550 310176
rect 29606 310120 36554 310176
rect 29545 310118 36554 310120
rect 29545 310115 29611 310118
rect 34329 310042 34395 310045
rect 34329 310040 35910 310042
rect 34329 309984 34334 310040
rect 34390 309984 35910 310040
rect 34329 309982 35910 309984
rect 34329 309979 34395 309982
rect 35850 309226 35910 309982
rect 36494 309362 36554 310118
rect 36721 310042 36787 310045
rect 36721 310040 45570 310042
rect 36721 309984 36726 310040
rect 36782 309984 45570 310040
rect 36721 309982 45570 309984
rect 36721 309979 36787 309982
rect 45510 309498 45570 309982
rect 302969 309498 303035 309501
rect 45510 309496 303035 309498
rect 45510 309440 302974 309496
rect 303030 309440 303035 309496
rect 45510 309438 303035 309440
rect 302969 309435 303035 309438
rect 315297 309362 315363 309365
rect 36494 309360 315363 309362
rect 36494 309304 315302 309360
rect 315358 309304 315363 309360
rect 36494 309302 315363 309304
rect 315297 309299 315363 309302
rect 580257 309226 580323 309229
rect 35850 309224 580323 309226
rect 35850 309168 580262 309224
rect 580318 309168 580323 309224
rect 35850 309166 580323 309168
rect 580257 309163 580323 309166
rect -960 306234 480 306324
rect 2957 306234 3023 306237
rect -960 306232 3023 306234
rect -960 306176 2962 306232
rect 3018 306176 3023 306232
rect -960 306174 3023 306176
rect -960 306084 480 306174
rect 2957 306171 3023 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579981 272234 580047 272237
rect 583520 272234 584960 272324
rect 579981 272232 584960 272234
rect 579981 272176 579986 272232
rect 580042 272176 584960 272232
rect 579981 272174 584960 272176
rect 579981 272171 580047 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2773 267202 2839 267205
rect -960 267200 2839 267202
rect -960 267144 2778 267200
rect 2834 267144 2839 267200
rect -960 267142 2839 267144
rect -960 267052 480 267142
rect 2773 267139 2839 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580901 219058 580967 219061
rect 583520 219058 584960 219148
rect 580901 219056 584960 219058
rect 580901 219000 580906 219056
rect 580962 219000 584960 219056
rect 580901 218998 584960 219000
rect 580901 218995 580967 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580809 192538 580875 192541
rect 583520 192538 584960 192628
rect 580809 192536 584960 192538
rect 580809 192480 580814 192536
rect 580870 192480 584960 192536
rect 580809 192478 584960 192480
rect 580809 192475 580875 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 4061 188866 4127 188869
rect -960 188864 4127 188866
rect -960 188808 4066 188864
rect 4122 188808 4127 188864
rect -960 188806 4127 188808
rect -960 188716 480 188806
rect 4061 188803 4127 188806
rect 580717 179210 580783 179213
rect 583520 179210 584960 179300
rect 580717 179208 584960 179210
rect 580717 179152 580722 179208
rect 580778 179152 584960 179208
rect 580717 179150 584960 179152
rect 580717 179147 580783 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3969 162890 4035 162893
rect -960 162888 4035 162890
rect -960 162832 3974 162888
rect 4030 162832 4035 162888
rect -960 162830 4035 162832
rect -960 162740 480 162830
rect 3969 162827 4035 162830
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 580625 139362 580691 139365
rect 583520 139362 584960 139452
rect 580625 139360 584960 139362
rect 580625 139304 580630 139360
rect 580686 139304 584960 139360
rect 580625 139302 584960 139304
rect 580625 139299 580691 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3877 136778 3943 136781
rect -960 136776 3943 136778
rect -960 136720 3882 136776
rect 3938 136720 3943 136776
rect -960 136718 3943 136720
rect -960 136628 480 136718
rect 3877 136715 3943 136718
rect 579705 126034 579771 126037
rect 583520 126034 584960 126124
rect 579705 126032 584960 126034
rect 579705 125976 579710 126032
rect 579766 125976 584960 126032
rect 579705 125974 584960 125976
rect 579705 125971 579771 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 2773 123722 2839 123725
rect -960 123720 2839 123722
rect -960 123664 2778 123720
rect 2834 123664 2839 123720
rect -960 123662 2839 123664
rect -960 123572 480 123662
rect 2773 123659 2839 123662
rect 580533 112842 580599 112845
rect 583520 112842 584960 112932
rect 580533 112840 584960 112842
rect 580533 112784 580538 112840
rect 580594 112784 584960 112840
rect 580533 112782 584960 112784
rect 580533 112779 580599 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 2773 110666 2839 110669
rect -960 110664 2839 110666
rect -960 110608 2778 110664
rect 2834 110608 2839 110664
rect -960 110606 2839 110608
rect -960 110516 480 110606
rect 2773 110603 2839 110606
rect 580441 99514 580507 99517
rect 583520 99514 584960 99604
rect 580441 99512 584960 99514
rect 580441 99456 580446 99512
rect 580502 99456 584960 99512
rect 580441 99454 584960 99456
rect 580441 99451 580507 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3785 97610 3851 97613
rect -960 97608 3851 97610
rect -960 97552 3790 97608
rect 3846 97552 3851 97608
rect -960 97550 3851 97552
rect -960 97460 480 97550
rect 3785 97547 3851 97550
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2773 71634 2839 71637
rect -960 71632 2839 71634
rect -960 71576 2778 71632
rect 2834 71576 2839 71632
rect -960 71574 2839 71576
rect -960 71484 480 71574
rect 2773 71571 2839 71574
rect 580349 59666 580415 59669
rect 583520 59666 584960 59756
rect 580349 59664 584960 59666
rect 580349 59608 580354 59664
rect 580410 59608 584960 59664
rect 580349 59606 584960 59608
rect 580349 59603 580415 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3693 58578 3759 58581
rect -960 58576 3759 58578
rect -960 58520 3698 58576
rect 3754 58520 3759 58576
rect -960 58518 3759 58520
rect -960 58428 480 58518
rect 3693 58515 3759 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3601 32466 3667 32469
rect -960 32464 3667 32466
rect -960 32408 3606 32464
rect 3662 32408 3667 32464
rect -960 32406 3667 32408
rect -960 32316 480 32406
rect 3601 32403 3667 32406
rect 302141 31378 302207 31381
rect 322197 31378 322263 31381
rect 302141 31376 322263 31378
rect 302141 31320 302146 31376
rect 302202 31320 322202 31376
rect 322258 31320 322263 31376
rect 302141 31318 322263 31320
rect 302141 31315 302207 31318
rect 322197 31315 322263 31318
rect 249057 31242 249123 31245
rect 323577 31242 323643 31245
rect 249057 31240 323643 31242
rect 249057 31184 249062 31240
rect 249118 31184 323582 31240
rect 323638 31184 323643 31240
rect 249057 31182 323643 31184
rect 249057 31179 249123 31182
rect 323577 31179 323643 31182
rect 252461 31106 252527 31109
rect 382917 31106 382983 31109
rect 252461 31104 382983 31106
rect 252461 31048 252466 31104
rect 252522 31048 382922 31104
rect 382978 31048 382983 31104
rect 252461 31046 382983 31048
rect 252461 31043 252527 31046
rect 382917 31043 382983 31046
rect 238753 30970 238819 30973
rect 380157 30970 380223 30973
rect 238753 30968 380223 30970
rect 238753 30912 238758 30968
rect 238814 30912 380162 30968
rect 380218 30912 380223 30968
rect 238753 30910 380223 30912
rect 238753 30907 238819 30910
rect 380157 30907 380223 30910
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 292481 14786 292547 14789
rect 560385 14786 560451 14789
rect 292481 14784 560451 14786
rect 292481 14728 292486 14784
rect 292542 14728 560390 14784
rect 560446 14728 560451 14784
rect 292481 14726 560451 14728
rect 292481 14723 292547 14726
rect 560385 14723 560451 14726
rect 297909 14650 297975 14653
rect 571517 14650 571583 14653
rect 297909 14648 571583 14650
rect 297909 14592 297914 14648
rect 297970 14592 571522 14648
rect 571578 14592 571583 14648
rect 297909 14590 571583 14592
rect 297909 14587 297975 14590
rect 571517 14587 571583 14590
rect 299197 14514 299263 14517
rect 575105 14514 575171 14517
rect 299197 14512 575171 14514
rect 299197 14456 299202 14512
rect 299258 14456 575110 14512
rect 575166 14456 575171 14512
rect 299197 14454 575171 14456
rect 299197 14451 299263 14454
rect 575105 14451 575171 14454
rect 282637 13426 282703 13429
rect 539593 13426 539659 13429
rect 282637 13424 539659 13426
rect 282637 13368 282642 13424
rect 282698 13368 539598 13424
rect 539654 13368 539659 13424
rect 282637 13366 539659 13368
rect 282637 13363 282703 13366
rect 539593 13363 539659 13366
rect 284109 13290 284175 13293
rect 542721 13290 542787 13293
rect 284109 13288 542787 13290
rect 284109 13232 284114 13288
rect 284170 13232 542726 13288
rect 542782 13232 542787 13288
rect 284109 13230 542787 13232
rect 284109 13227 284175 13230
rect 542721 13227 542787 13230
rect 288157 13154 288223 13157
rect 550265 13154 550331 13157
rect 288157 13152 550331 13154
rect 288157 13096 288162 13152
rect 288218 13096 550270 13152
rect 550326 13096 550331 13152
rect 288157 13094 550331 13096
rect 288157 13091 288223 13094
rect 550265 13091 550331 13094
rect 293677 13018 293743 13021
rect 564433 13018 564499 13021
rect 293677 13016 564499 13018
rect 293677 12960 293682 13016
rect 293738 12960 564438 13016
rect 564494 12960 564499 13016
rect 293677 12958 564499 12960
rect 293677 12955 293743 12958
rect 564433 12955 564499 12958
rect 268929 12066 268995 12069
rect 511257 12066 511323 12069
rect 268929 12064 511323 12066
rect 268929 12008 268934 12064
rect 268990 12008 511262 12064
rect 511318 12008 511323 12064
rect 268929 12006 511323 12008
rect 268929 12003 268995 12006
rect 511257 12003 511323 12006
rect 273069 11930 273135 11933
rect 517881 11930 517947 11933
rect 273069 11928 517947 11930
rect 273069 11872 273074 11928
rect 273130 11872 517886 11928
rect 517942 11872 517947 11928
rect 273069 11870 517947 11872
rect 273069 11867 273135 11870
rect 517881 11867 517947 11870
rect 270217 11794 270283 11797
rect 514753 11794 514819 11797
rect 270217 11792 514819 11794
rect 270217 11736 270222 11792
rect 270278 11736 514758 11792
rect 514814 11736 514819 11792
rect 270217 11734 514819 11736
rect 270217 11731 270283 11734
rect 514753 11731 514819 11734
rect 274357 11658 274423 11661
rect 521837 11658 521903 11661
rect 274357 11656 521903 11658
rect 274357 11600 274362 11656
rect 274418 11600 521842 11656
rect 521898 11600 521903 11656
rect 274357 11598 521903 11600
rect 274357 11595 274423 11598
rect 521837 11595 521903 11598
rect 220629 10706 220695 10709
rect 407205 10706 407271 10709
rect 220629 10704 407271 10706
rect 220629 10648 220634 10704
rect 220690 10648 407210 10704
rect 407266 10648 407271 10704
rect 220629 10646 407271 10648
rect 220629 10643 220695 10646
rect 407205 10643 407271 10646
rect 222009 10570 222075 10573
rect 410793 10570 410859 10573
rect 222009 10568 410859 10570
rect 222009 10512 222014 10568
rect 222070 10512 410798 10568
rect 410854 10512 410859 10568
rect 222009 10510 410859 10512
rect 222009 10507 222075 10510
rect 410793 10507 410859 10510
rect 223389 10434 223455 10437
rect 414289 10434 414355 10437
rect 223389 10432 414355 10434
rect 223389 10376 223394 10432
rect 223450 10376 414294 10432
rect 414350 10376 414355 10432
rect 223389 10374 414355 10376
rect 223389 10371 223455 10374
rect 414289 10371 414355 10374
rect 224677 10298 224743 10301
rect 417417 10298 417483 10301
rect 224677 10296 417483 10298
rect 224677 10240 224682 10296
rect 224738 10240 417422 10296
rect 417478 10240 417483 10296
rect 224677 10238 417483 10240
rect 224677 10235 224743 10238
rect 417417 10235 417483 10238
rect 176561 9346 176627 9349
rect 315021 9346 315087 9349
rect 176561 9344 315087 9346
rect 176561 9288 176566 9344
rect 176622 9288 315026 9344
rect 315082 9288 315087 9344
rect 176561 9286 315087 9288
rect 176561 9283 176627 9286
rect 315021 9283 315087 9286
rect 179229 9210 179295 9213
rect 318517 9210 318583 9213
rect 179229 9208 318583 9210
rect 179229 9152 179234 9208
rect 179290 9152 318522 9208
rect 318578 9152 318583 9208
rect 179229 9150 318583 9152
rect 179229 9147 179295 9150
rect 318517 9147 318583 9150
rect 180701 9074 180767 9077
rect 322105 9074 322171 9077
rect 180701 9072 322171 9074
rect 180701 9016 180706 9072
rect 180762 9016 322110 9072
rect 322166 9016 322171 9072
rect 180701 9014 322171 9016
rect 180701 9011 180767 9014
rect 322105 9011 322171 9014
rect 288249 8938 288315 8941
rect 552657 8938 552723 8941
rect 288249 8936 552723 8938
rect 288249 8880 288254 8936
rect 288310 8880 552662 8936
rect 552718 8880 552723 8936
rect 288249 8878 552723 8880
rect 288249 8875 288315 8878
rect 552657 8875 552723 8878
rect 238661 7986 238727 7989
rect 445017 7986 445083 7989
rect 238661 7984 445083 7986
rect 238661 7928 238666 7984
rect 238722 7928 445022 7984
rect 445078 7928 445083 7984
rect 238661 7926 445083 7928
rect 238661 7923 238727 7926
rect 445017 7923 445083 7926
rect 240041 7850 240107 7853
rect 448605 7850 448671 7853
rect 240041 7848 448671 7850
rect 240041 7792 240046 7848
rect 240102 7792 448610 7848
rect 448666 7792 448671 7848
rect 240041 7790 448671 7792
rect 240041 7787 240107 7790
rect 448605 7787 448671 7790
rect 241421 7714 241487 7717
rect 452101 7714 452167 7717
rect 241421 7712 452167 7714
rect 241421 7656 241426 7712
rect 241482 7656 452106 7712
rect 452162 7656 452167 7712
rect 241421 7654 452167 7656
rect 241421 7651 241487 7654
rect 452101 7651 452167 7654
rect 246941 7578 247007 7581
rect 462773 7578 462839 7581
rect 246941 7576 462839 7578
rect 246941 7520 246946 7576
rect 247002 7520 462778 7576
rect 462834 7520 462839 7576
rect 246941 7518 462839 7520
rect 246941 7515 247007 7518
rect 462773 7515 462839 7518
rect 148961 6626 149027 6629
rect 254669 6626 254735 6629
rect 148961 6624 254735 6626
rect -960 6490 480 6580
rect 148961 6568 148966 6624
rect 149022 6568 254674 6624
rect 254730 6568 254735 6624
rect 148961 6566 254735 6568
rect 148961 6563 149027 6566
rect 254669 6563 254735 6566
rect 278589 6626 278655 6629
rect 531313 6626 531379 6629
rect 278589 6624 531379 6626
rect 278589 6568 278594 6624
rect 278650 6568 531318 6624
rect 531374 6568 531379 6624
rect 278589 6566 531379 6568
rect 278589 6563 278655 6566
rect 531313 6563 531379 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 150249 6490 150315 6493
rect 258257 6490 258323 6493
rect 150249 6488 258323 6490
rect 150249 6432 150254 6488
rect 150310 6432 258262 6488
rect 258318 6432 258323 6488
rect 150249 6430 258323 6432
rect 150249 6427 150315 6430
rect 258257 6427 258323 6430
rect 285489 6490 285555 6493
rect 545481 6490 545547 6493
rect 285489 6488 545547 6490
rect 285489 6432 285494 6488
rect 285550 6432 545486 6488
rect 545542 6432 545547 6488
rect 583520 6476 584960 6566
rect 285489 6430 545547 6432
rect 285489 6427 285555 6430
rect 545481 6427 545547 6430
rect 153009 6354 153075 6357
rect 265341 6354 265407 6357
rect 153009 6352 265407 6354
rect 153009 6296 153014 6352
rect 153070 6296 265346 6352
rect 265402 6296 265407 6352
rect 153009 6294 265407 6296
rect 153009 6291 153075 6294
rect 265341 6291 265407 6294
rect 291009 6354 291075 6357
rect 556153 6354 556219 6357
rect 291009 6352 556219 6354
rect 291009 6296 291014 6352
rect 291070 6296 556158 6352
rect 556214 6296 556219 6352
rect 291009 6294 556219 6296
rect 291009 6291 291075 6294
rect 556153 6291 556219 6294
rect 157241 6218 157307 6221
rect 272425 6218 272491 6221
rect 157241 6216 272491 6218
rect 157241 6160 157246 6216
rect 157302 6160 272430 6216
rect 272486 6160 272491 6216
rect 157241 6158 272491 6160
rect 157241 6155 157307 6158
rect 272425 6155 272491 6158
rect 296529 6218 296595 6221
rect 570321 6218 570387 6221
rect 296529 6216 570387 6218
rect 296529 6160 296534 6216
rect 296590 6160 570326 6216
rect 570382 6160 570387 6216
rect 296529 6158 570387 6160
rect 296529 6155 296595 6158
rect 570321 6155 570387 6158
rect 195881 5266 195947 5269
rect 356329 5266 356395 5269
rect 195881 5264 356395 5266
rect 195881 5208 195886 5264
rect 195942 5208 356334 5264
rect 356390 5208 356395 5264
rect 195881 5206 356395 5208
rect 195881 5203 195947 5206
rect 356329 5203 356395 5206
rect 139301 5130 139367 5133
rect 235809 5130 235875 5133
rect 139301 5128 235875 5130
rect 139301 5072 139306 5128
rect 139362 5072 235814 5128
rect 235870 5072 235875 5128
rect 139301 5070 235875 5072
rect 139301 5067 139367 5070
rect 235809 5067 235875 5070
rect 289721 5130 289787 5133
rect 554957 5130 555023 5133
rect 289721 5128 555023 5130
rect 289721 5072 289726 5128
rect 289782 5072 554962 5128
rect 555018 5072 555023 5128
rect 289721 5070 555023 5072
rect 289721 5067 289787 5070
rect 554957 5067 555023 5070
rect 151721 4994 151787 4997
rect 260649 4994 260715 4997
rect 151721 4992 260715 4994
rect 151721 4936 151726 4992
rect 151782 4936 260654 4992
rect 260710 4936 260715 4992
rect 151721 4934 260715 4936
rect 151721 4931 151787 4934
rect 260649 4931 260715 4934
rect 291101 4994 291167 4997
rect 558545 4994 558611 4997
rect 291101 4992 558611 4994
rect 291101 4936 291106 4992
rect 291162 4936 558550 4992
rect 558606 4936 558611 4992
rect 291101 4934 558611 4936
rect 291101 4931 291167 4934
rect 558545 4931 558611 4934
rect 154481 4858 154547 4861
rect 267733 4858 267799 4861
rect 154481 4856 267799 4858
rect 154481 4800 154486 4856
rect 154542 4800 267738 4856
rect 267794 4800 267799 4856
rect 154481 4798 267799 4800
rect 154481 4795 154547 4798
rect 267733 4795 267799 4798
rect 298001 4858 298067 4861
rect 572713 4858 572779 4861
rect 298001 4856 572779 4858
rect 298001 4800 298006 4856
rect 298062 4800 572718 4856
rect 572774 4800 572779 4856
rect 298001 4798 572779 4800
rect 298001 4795 298067 4798
rect 572713 4795 572779 4798
rect 131021 3770 131087 3773
rect 216857 3770 216923 3773
rect 131021 3768 216923 3770
rect 131021 3712 131026 3768
rect 131082 3712 216862 3768
rect 216918 3712 216923 3768
rect 131021 3710 216923 3712
rect 131021 3707 131087 3710
rect 216857 3707 216923 3710
rect 79777 3634 79843 3637
rect 110505 3634 110571 3637
rect 79777 3632 110571 3634
rect 79777 3576 79782 3632
rect 79838 3576 110510 3632
rect 110566 3576 110571 3632
rect 79777 3574 110571 3576
rect 79777 3571 79843 3574
rect 110505 3571 110571 3574
rect 133781 3634 133847 3637
rect 223941 3634 224007 3637
rect 133781 3632 224007 3634
rect 133781 3576 133786 3632
rect 133842 3576 223946 3632
rect 224002 3576 224007 3632
rect 133781 3574 224007 3576
rect 133781 3571 133847 3574
rect 223941 3571 224007 3574
rect 323577 3634 323643 3637
rect 468661 3634 468727 3637
rect 323577 3632 468727 3634
rect 323577 3576 323582 3632
rect 323638 3576 468666 3632
rect 468722 3576 468727 3632
rect 323577 3574 468727 3576
rect 323577 3571 323643 3574
rect 468661 3571 468727 3574
rect 84009 3498 84075 3501
rect 117589 3498 117655 3501
rect 84009 3496 117655 3498
rect 84009 3440 84014 3496
rect 84070 3440 117594 3496
rect 117650 3440 117655 3496
rect 84009 3438 117655 3440
rect 84009 3435 84075 3438
rect 117589 3435 117655 3438
rect 135161 3498 135227 3501
rect 227529 3498 227595 3501
rect 135161 3496 227595 3498
rect 135161 3440 135166 3496
rect 135222 3440 227534 3496
rect 227590 3440 227595 3496
rect 135161 3438 227595 3440
rect 135161 3435 135227 3438
rect 227529 3435 227595 3438
rect 251081 3498 251147 3501
rect 472249 3498 472315 3501
rect 251081 3496 472315 3498
rect 251081 3440 251086 3496
rect 251142 3440 472254 3496
rect 472310 3440 472315 3496
rect 251081 3438 472315 3440
rect 251081 3435 251147 3438
rect 472249 3435 472315 3438
rect 84101 3362 84167 3365
rect 118785 3362 118851 3365
rect 84101 3360 118851 3362
rect 84101 3304 84106 3360
rect 84162 3304 118790 3360
rect 118846 3304 118851 3360
rect 84101 3302 118851 3304
rect 84101 3299 84167 3302
rect 118785 3299 118851 3302
rect 140681 3362 140747 3365
rect 238109 3362 238175 3365
rect 140681 3360 238175 3362
rect 140681 3304 140686 3360
rect 140742 3304 238114 3360
rect 238170 3304 238175 3360
rect 140681 3302 238175 3304
rect 140681 3299 140747 3302
rect 238109 3299 238175 3302
rect 253841 3362 253907 3365
rect 479333 3362 479399 3365
rect 253841 3360 479399 3362
rect 253841 3304 253846 3360
rect 253902 3304 479338 3360
rect 479394 3304 479399 3360
rect 253841 3302 479399 3304
rect 253841 3299 253907 3302
rect 479333 3299 479399 3302
rect 348417 3226 348483 3229
rect 351821 3226 351887 3229
rect 348417 3224 351887 3226
rect 348417 3168 348422 3224
rect 348478 3168 351826 3224
rect 351882 3168 351887 3224
rect 348417 3166 351887 3168
rect 348417 3163 348483 3166
rect 351821 3163 351887 3166
<< metal4 >>
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 675364 38414 686898
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 675364 56414 705242
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 675364 74414 686898
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 675364 92414 705242
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 675364 110414 686898
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 675364 128414 705242
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 675364 146414 686898
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 675364 164414 705242
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 675364 182414 686898
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 675364 200414 705242
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 675364 218414 686898
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 675364 236414 705242
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 675364 254414 686898
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 53494 669454 55628 669486
rect 53494 669218 53643 669454
rect 53879 669218 53963 669454
rect 54199 669218 54283 669454
rect 54519 669218 54603 669454
rect 54839 669218 54923 669454
rect 55159 669218 55243 669454
rect 55479 669218 55628 669454
rect 53494 669134 55628 669218
rect 53494 668898 53643 669134
rect 53879 668898 53963 669134
rect 54199 668898 54283 669134
rect 54519 668898 54603 669134
rect 54839 668898 54923 669134
rect 55159 668898 55243 669134
rect 55479 668898 55628 669134
rect 53494 668866 55628 668898
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 36912 633454 44282 633486
rect 36912 633218 36959 633454
rect 37195 633218 37279 633454
rect 37515 633218 37599 633454
rect 37835 633218 37919 633454
rect 38155 633218 38239 633454
rect 38475 633218 38559 633454
rect 38795 633218 38879 633454
rect 39115 633218 39199 633454
rect 39435 633218 39519 633454
rect 39755 633218 39839 633454
rect 40075 633218 40159 633454
rect 40395 633218 40479 633454
rect 40715 633218 40799 633454
rect 41035 633218 41119 633454
rect 41355 633218 41439 633454
rect 41675 633218 41759 633454
rect 41995 633218 42079 633454
rect 42315 633218 42399 633454
rect 42635 633218 42719 633454
rect 42955 633218 43039 633454
rect 43275 633218 43359 633454
rect 43595 633218 43679 633454
rect 43915 633218 43999 633454
rect 44235 633218 44282 633454
rect 36912 633134 44282 633218
rect 36912 632898 36959 633134
rect 37195 632898 37279 633134
rect 37515 632898 37599 633134
rect 37835 632898 37919 633134
rect 38155 632898 38239 633134
rect 38475 632898 38559 633134
rect 38795 632898 38879 633134
rect 39115 632898 39199 633134
rect 39435 632898 39519 633134
rect 39755 632898 39839 633134
rect 40075 632898 40159 633134
rect 40395 632898 40479 633134
rect 40715 632898 40799 633134
rect 41035 632898 41119 633134
rect 41355 632898 41439 633134
rect 41675 632898 41759 633134
rect 41995 632898 42079 633134
rect 42315 632898 42399 633134
rect 42635 632898 42719 633134
rect 42955 632898 43039 633134
rect 43275 632898 43359 633134
rect 43595 632898 43679 633134
rect 43915 632898 43999 633134
rect 44235 632898 44282 633134
rect 36912 632866 44282 632898
rect 261496 633454 266930 633486
rect 261496 633218 261535 633454
rect 261771 633218 261855 633454
rect 262091 633218 262175 633454
rect 262411 633218 262495 633454
rect 262731 633218 262815 633454
rect 263051 633218 263135 633454
rect 263371 633218 263455 633454
rect 263691 633218 263775 633454
rect 264011 633218 264095 633454
rect 264331 633218 264415 633454
rect 264651 633218 264735 633454
rect 264971 633218 265055 633454
rect 265291 633218 265375 633454
rect 265611 633218 265695 633454
rect 265931 633218 266015 633454
rect 266251 633218 266335 633454
rect 266571 633218 266655 633454
rect 266891 633218 266930 633454
rect 261496 633134 266930 633218
rect 261496 632898 261535 633134
rect 261771 632898 261855 633134
rect 262091 632898 262175 633134
rect 262411 632898 262495 633134
rect 262731 632898 262815 633134
rect 263051 632898 263135 633134
rect 263371 632898 263455 633134
rect 263691 632898 263775 633134
rect 264011 632898 264095 633134
rect 264331 632898 264415 633134
rect 264651 632898 264735 633134
rect 264971 632898 265055 633134
rect 265291 632898 265375 633134
rect 265611 632898 265695 633134
rect 265931 632898 266015 633134
rect 266251 632898 266335 633134
rect 266571 632898 266655 633134
rect 266891 632898 266930 633134
rect 261496 632866 266930 632898
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 47300 615454 53316 615486
rect 47300 615218 47470 615454
rect 47706 615218 47790 615454
rect 48026 615218 48110 615454
rect 48346 615218 48430 615454
rect 48666 615218 48750 615454
rect 48986 615218 49070 615454
rect 49306 615218 49390 615454
rect 49626 615218 49710 615454
rect 49946 615218 50030 615454
rect 50266 615218 50350 615454
rect 50586 615218 50670 615454
rect 50906 615218 50990 615454
rect 51226 615218 51310 615454
rect 51546 615218 51630 615454
rect 51866 615218 51950 615454
rect 52186 615218 52270 615454
rect 52506 615218 52590 615454
rect 52826 615218 52910 615454
rect 53146 615218 53316 615454
rect 47300 615134 53316 615218
rect 47300 614898 47470 615134
rect 47706 614898 47790 615134
rect 48026 614898 48110 615134
rect 48346 614898 48430 615134
rect 48666 614898 48750 615134
rect 48986 614898 49070 615134
rect 49306 614898 49390 615134
rect 49626 614898 49710 615134
rect 49946 614898 50030 615134
rect 50266 614898 50350 615134
rect 50586 614898 50670 615134
rect 50906 614898 50990 615134
rect 51226 614898 51310 615134
rect 51546 614898 51630 615134
rect 51866 614898 51950 615134
rect 52186 614898 52270 615134
rect 52506 614898 52590 615134
rect 52826 614898 52910 615134
rect 53146 614898 53316 615134
rect 47300 614866 53316 614898
rect 253294 615454 258068 615486
rect 253294 615218 253323 615454
rect 253559 615218 253643 615454
rect 253879 615218 253963 615454
rect 254199 615218 254283 615454
rect 254519 615218 254603 615454
rect 254839 615218 254923 615454
rect 255159 615218 255243 615454
rect 255479 615218 255563 615454
rect 255799 615218 255883 615454
rect 256119 615218 256203 615454
rect 256439 615218 256523 615454
rect 256759 615218 256843 615454
rect 257079 615218 257163 615454
rect 257399 615218 257483 615454
rect 257719 615218 257803 615454
rect 258039 615218 258068 615454
rect 253294 615134 258068 615218
rect 253294 614898 253323 615134
rect 253559 614898 253643 615134
rect 253879 614898 253963 615134
rect 254199 614898 254283 615134
rect 254519 614898 254603 615134
rect 254839 614898 254923 615134
rect 255159 614898 255243 615134
rect 255479 614898 255563 615134
rect 255799 614898 255883 615134
rect 256119 614898 256203 615134
rect 256439 614898 256523 615134
rect 256759 614898 256843 615134
rect 257079 614898 257163 615134
rect 257399 614898 257483 615134
rect 257719 614898 257803 615134
rect 258039 614898 258068 615134
rect 253294 614866 258068 614898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 36912 597454 44282 597486
rect 36912 597218 36959 597454
rect 37195 597218 37279 597454
rect 37515 597218 37599 597454
rect 37835 597218 37919 597454
rect 38155 597218 38239 597454
rect 38475 597218 38559 597454
rect 38795 597218 38879 597454
rect 39115 597218 39199 597454
rect 39435 597218 39519 597454
rect 39755 597218 39839 597454
rect 40075 597218 40159 597454
rect 40395 597218 40479 597454
rect 40715 597218 40799 597454
rect 41035 597218 41119 597454
rect 41355 597218 41439 597454
rect 41675 597218 41759 597454
rect 41995 597218 42079 597454
rect 42315 597218 42399 597454
rect 42635 597218 42719 597454
rect 42955 597218 43039 597454
rect 43275 597218 43359 597454
rect 43595 597218 43679 597454
rect 43915 597218 43999 597454
rect 44235 597218 44282 597454
rect 36912 597134 44282 597218
rect 36912 596898 36959 597134
rect 37195 596898 37279 597134
rect 37515 596898 37599 597134
rect 37835 596898 37919 597134
rect 38155 596898 38239 597134
rect 38475 596898 38559 597134
rect 38795 596898 38879 597134
rect 39115 596898 39199 597134
rect 39435 596898 39519 597134
rect 39755 596898 39839 597134
rect 40075 596898 40159 597134
rect 40395 596898 40479 597134
rect 40715 596898 40799 597134
rect 41035 596898 41119 597134
rect 41355 596898 41439 597134
rect 41675 596898 41759 597134
rect 41995 596898 42079 597134
rect 42315 596898 42399 597134
rect 42635 596898 42719 597134
rect 42955 596898 43039 597134
rect 43275 596898 43359 597134
rect 43595 596898 43679 597134
rect 43915 596898 43999 597134
rect 44235 596898 44282 597134
rect 36912 596866 44282 596898
rect 167626 597454 167862 597486
rect 167626 597134 167862 597218
rect 167626 596866 167862 596898
rect 171918 597454 172154 597486
rect 171918 597134 172154 597218
rect 171918 596866 172154 596898
rect 176210 597454 176446 597486
rect 176210 597134 176446 597218
rect 176210 596866 176446 596898
rect 180502 597454 180738 597486
rect 180502 597134 180738 597218
rect 180502 596866 180738 596898
rect 184794 597454 185030 597486
rect 184794 597134 185030 597218
rect 184794 596866 185030 596898
rect 189366 597454 189602 597486
rect 189366 597134 189602 597218
rect 189366 596866 189602 596898
rect 193658 597454 193894 597486
rect 193658 597134 193894 597218
rect 193658 596866 193894 596898
rect 197950 597454 198186 597486
rect 197950 597134 198186 597218
rect 197950 596866 198186 596898
rect 202242 597454 202478 597486
rect 202242 597134 202478 597218
rect 202242 596866 202478 596898
rect 206534 597454 206770 597486
rect 206534 597134 206770 597218
rect 206534 596866 206770 596898
rect 211138 597454 211374 597486
rect 211138 597134 211374 597218
rect 211138 596866 211374 596898
rect 215430 597454 215666 597486
rect 215430 597134 215666 597218
rect 215430 596866 215666 596898
rect 219722 597454 219958 597486
rect 219722 597134 219958 597218
rect 219722 596866 219958 596898
rect 224014 597454 224250 597486
rect 224014 597134 224250 597218
rect 224014 596866 224250 596898
rect 228306 597454 228542 597486
rect 228306 597134 228542 597218
rect 228306 596866 228542 596898
rect 232826 597454 233062 597486
rect 232826 597134 233062 597218
rect 232826 596866 233062 596898
rect 237118 597454 237354 597486
rect 237118 597134 237354 597218
rect 237118 596866 237354 596898
rect 241410 597454 241646 597486
rect 241410 597134 241646 597218
rect 241410 596866 241646 596898
rect 245702 597454 245938 597486
rect 245702 597134 245938 597218
rect 245702 596866 245938 596898
rect 249994 597454 250230 597486
rect 249994 597134 250230 597218
rect 249994 596866 250230 596898
rect 261496 597454 266930 597486
rect 261496 597218 261535 597454
rect 261771 597218 261855 597454
rect 262091 597218 262175 597454
rect 262411 597218 262495 597454
rect 262731 597218 262815 597454
rect 263051 597218 263135 597454
rect 263371 597218 263455 597454
rect 263691 597218 263775 597454
rect 264011 597218 264095 597454
rect 264331 597218 264415 597454
rect 264651 597218 264735 597454
rect 264971 597218 265055 597454
rect 265291 597218 265375 597454
rect 265611 597218 265695 597454
rect 265931 597218 266015 597454
rect 266251 597218 266335 597454
rect 266571 597218 266655 597454
rect 266891 597218 266930 597454
rect 261496 597134 266930 597218
rect 261496 596898 261535 597134
rect 261771 596898 261855 597134
rect 262091 596898 262175 597134
rect 262411 596898 262495 597134
rect 262731 596898 262815 597134
rect 263051 596898 263135 597134
rect 263371 596898 263455 597134
rect 263691 596898 263775 597134
rect 264011 596898 264095 597134
rect 264331 596898 264415 597134
rect 264651 596898 264735 597134
rect 264971 596898 265055 597134
rect 265291 596898 265375 597134
rect 265611 596898 265695 597134
rect 265931 596898 266015 597134
rect 266251 596898 266335 597134
rect 266571 596898 266655 597134
rect 266891 596898 266930 597134
rect 261496 596866 266930 596898
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 47300 579454 53316 579486
rect 47300 579218 47470 579454
rect 47706 579218 47790 579454
rect 48026 579218 48110 579454
rect 48346 579218 48430 579454
rect 48666 579218 48750 579454
rect 48986 579218 49070 579454
rect 49306 579218 49390 579454
rect 49626 579218 49710 579454
rect 49946 579218 50030 579454
rect 50266 579218 50350 579454
rect 50586 579218 50670 579454
rect 50906 579218 50990 579454
rect 51226 579218 51310 579454
rect 51546 579218 51630 579454
rect 51866 579218 51950 579454
rect 52186 579218 52270 579454
rect 52506 579218 52590 579454
rect 52826 579218 52910 579454
rect 53146 579218 53316 579454
rect 47300 579134 53316 579218
rect 47300 578898 47470 579134
rect 47706 578898 47790 579134
rect 48026 578898 48110 579134
rect 48346 578898 48430 579134
rect 48666 578898 48750 579134
rect 48986 578898 49070 579134
rect 49306 578898 49390 579134
rect 49626 578898 49710 579134
rect 49946 578898 50030 579134
rect 50266 578898 50350 579134
rect 50586 578898 50670 579134
rect 50906 578898 50990 579134
rect 51226 578898 51310 579134
rect 51546 578898 51630 579134
rect 51866 578898 51950 579134
rect 52186 578898 52270 579134
rect 52506 578898 52590 579134
rect 52826 578898 52910 579134
rect 53146 578898 53316 579134
rect 47300 578866 53316 578898
rect 253294 579454 258068 579486
rect 253294 579218 253323 579454
rect 253559 579218 253643 579454
rect 253879 579218 253963 579454
rect 254199 579218 254283 579454
rect 254519 579218 254603 579454
rect 254839 579218 254923 579454
rect 255159 579218 255243 579454
rect 255479 579218 255563 579454
rect 255799 579218 255883 579454
rect 256119 579218 256203 579454
rect 256439 579218 256523 579454
rect 256759 579218 256843 579454
rect 257079 579218 257163 579454
rect 257399 579218 257483 579454
rect 257719 579218 257803 579454
rect 258039 579218 258068 579454
rect 253294 579134 258068 579218
rect 253294 578898 253323 579134
rect 253559 578898 253643 579134
rect 253879 578898 253963 579134
rect 254199 578898 254283 579134
rect 254519 578898 254603 579134
rect 254839 578898 254923 579134
rect 255159 578898 255243 579134
rect 255479 578898 255563 579134
rect 255799 578898 255883 579134
rect 256119 578898 256203 579134
rect 256439 578898 256523 579134
rect 256759 578898 256843 579134
rect 257079 578898 257163 579134
rect 257399 578898 257483 579134
rect 257719 578898 257803 579134
rect 258039 578898 258068 579134
rect 253294 578866 258068 578898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 37794 543454 38414 552000
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 312712 38414 326898
rect 55794 525454 56414 552000
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 312712 56414 344898
rect 73794 543454 74414 552000
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 312712 74414 326898
rect 91794 525454 92414 552000
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 312712 92414 344898
rect 109794 543454 110414 552000
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 312712 110414 326898
rect 127794 525454 128414 552000
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 312712 128414 344898
rect 145794 543454 146414 552000
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 312712 146414 326898
rect 163794 525454 164414 552000
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 312712 164414 344898
rect 181794 543454 182414 552000
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 312712 182414 326898
rect 199794 525454 200414 552000
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 312712 200414 344898
rect 217794 543454 218414 552000
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 312712 218414 326898
rect 235794 525454 236414 552000
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 312712 236414 344898
rect 253794 543454 254414 552000
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 312712 254414 326898
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 312712 272414 344898
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 312712 290414 326898
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 32208 291454 32528 291486
rect 32208 291218 32250 291454
rect 32486 291218 32528 291454
rect 32208 291134 32528 291218
rect 32208 290898 32250 291134
rect 32486 290898 32528 291134
rect 32208 290866 32528 290898
rect 62928 291454 63248 291486
rect 62928 291218 62970 291454
rect 63206 291218 63248 291454
rect 62928 291134 63248 291218
rect 62928 290898 62970 291134
rect 63206 290898 63248 291134
rect 62928 290866 63248 290898
rect 93648 291454 93968 291486
rect 93648 291218 93690 291454
rect 93926 291218 93968 291454
rect 93648 291134 93968 291218
rect 93648 290898 93690 291134
rect 93926 290898 93968 291134
rect 93648 290866 93968 290898
rect 124368 291454 124688 291486
rect 124368 291218 124410 291454
rect 124646 291218 124688 291454
rect 124368 291134 124688 291218
rect 124368 290898 124410 291134
rect 124646 290898 124688 291134
rect 124368 290866 124688 290898
rect 155088 291454 155408 291486
rect 155088 291218 155130 291454
rect 155366 291218 155408 291454
rect 155088 291134 155408 291218
rect 155088 290898 155130 291134
rect 155366 290898 155408 291134
rect 155088 290866 155408 290898
rect 185808 291454 186128 291486
rect 185808 291218 185850 291454
rect 186086 291218 186128 291454
rect 185808 291134 186128 291218
rect 185808 290898 185850 291134
rect 186086 290898 186128 291134
rect 185808 290866 186128 290898
rect 216528 291454 216848 291486
rect 216528 291218 216570 291454
rect 216806 291218 216848 291454
rect 216528 291134 216848 291218
rect 216528 290898 216570 291134
rect 216806 290898 216848 291134
rect 216528 290866 216848 290898
rect 247248 291454 247568 291486
rect 247248 291218 247290 291454
rect 247526 291218 247568 291454
rect 247248 291134 247568 291218
rect 247248 290898 247290 291134
rect 247526 290898 247568 291134
rect 247248 290866 247568 290898
rect 277968 291454 278288 291486
rect 277968 291218 278010 291454
rect 278246 291218 278288 291454
rect 277968 291134 278288 291218
rect 277968 290898 278010 291134
rect 278246 290898 278288 291134
rect 277968 290866 278288 290898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 47568 273454 47888 273486
rect 47568 273218 47610 273454
rect 47846 273218 47888 273454
rect 47568 273134 47888 273218
rect 47568 272898 47610 273134
rect 47846 272898 47888 273134
rect 47568 272866 47888 272898
rect 78288 273454 78608 273486
rect 78288 273218 78330 273454
rect 78566 273218 78608 273454
rect 78288 273134 78608 273218
rect 78288 272898 78330 273134
rect 78566 272898 78608 273134
rect 78288 272866 78608 272898
rect 109008 273454 109328 273486
rect 109008 273218 109050 273454
rect 109286 273218 109328 273454
rect 109008 273134 109328 273218
rect 109008 272898 109050 273134
rect 109286 272898 109328 273134
rect 109008 272866 109328 272898
rect 139728 273454 140048 273486
rect 139728 273218 139770 273454
rect 140006 273218 140048 273454
rect 139728 273134 140048 273218
rect 139728 272898 139770 273134
rect 140006 272898 140048 273134
rect 139728 272866 140048 272898
rect 170448 273454 170768 273486
rect 170448 273218 170490 273454
rect 170726 273218 170768 273454
rect 170448 273134 170768 273218
rect 170448 272898 170490 273134
rect 170726 272898 170768 273134
rect 170448 272866 170768 272898
rect 201168 273454 201488 273486
rect 201168 273218 201210 273454
rect 201446 273218 201488 273454
rect 201168 273134 201488 273218
rect 201168 272898 201210 273134
rect 201446 272898 201488 273134
rect 201168 272866 201488 272898
rect 231888 273454 232208 273486
rect 231888 273218 231930 273454
rect 232166 273218 232208 273454
rect 231888 273134 232208 273218
rect 231888 272898 231930 273134
rect 232166 272898 232208 273134
rect 231888 272866 232208 272898
rect 262608 273454 262928 273486
rect 262608 273218 262650 273454
rect 262886 273218 262928 273454
rect 262608 273134 262928 273218
rect 262608 272898 262650 273134
rect 262886 272898 262928 273134
rect 262608 272866 262928 272898
rect 293328 273454 293648 273486
rect 293328 273218 293370 273454
rect 293606 273218 293648 273454
rect 293328 273134 293648 273218
rect 293328 272898 293370 273134
rect 293606 272898 293648 273134
rect 293328 272866 293648 272898
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 32208 255454 32528 255486
rect 32208 255218 32250 255454
rect 32486 255218 32528 255454
rect 32208 255134 32528 255218
rect 32208 254898 32250 255134
rect 32486 254898 32528 255134
rect 32208 254866 32528 254898
rect 62928 255454 63248 255486
rect 62928 255218 62970 255454
rect 63206 255218 63248 255454
rect 62928 255134 63248 255218
rect 62928 254898 62970 255134
rect 63206 254898 63248 255134
rect 62928 254866 63248 254898
rect 93648 255454 93968 255486
rect 93648 255218 93690 255454
rect 93926 255218 93968 255454
rect 93648 255134 93968 255218
rect 93648 254898 93690 255134
rect 93926 254898 93968 255134
rect 93648 254866 93968 254898
rect 124368 255454 124688 255486
rect 124368 255218 124410 255454
rect 124646 255218 124688 255454
rect 124368 255134 124688 255218
rect 124368 254898 124410 255134
rect 124646 254898 124688 255134
rect 124368 254866 124688 254898
rect 155088 255454 155408 255486
rect 155088 255218 155130 255454
rect 155366 255218 155408 255454
rect 155088 255134 155408 255218
rect 155088 254898 155130 255134
rect 155366 254898 155408 255134
rect 155088 254866 155408 254898
rect 185808 255454 186128 255486
rect 185808 255218 185850 255454
rect 186086 255218 186128 255454
rect 185808 255134 186128 255218
rect 185808 254898 185850 255134
rect 186086 254898 186128 255134
rect 185808 254866 186128 254898
rect 216528 255454 216848 255486
rect 216528 255218 216570 255454
rect 216806 255218 216848 255454
rect 216528 255134 216848 255218
rect 216528 254898 216570 255134
rect 216806 254898 216848 255134
rect 216528 254866 216848 254898
rect 247248 255454 247568 255486
rect 247248 255218 247290 255454
rect 247526 255218 247568 255454
rect 247248 255134 247568 255218
rect 247248 254898 247290 255134
rect 247526 254898 247568 255134
rect 247248 254866 247568 254898
rect 277968 255454 278288 255486
rect 277968 255218 278010 255454
rect 278246 255218 278288 255454
rect 277968 255134 278288 255218
rect 277968 254898 278010 255134
rect 278246 254898 278288 255134
rect 277968 254866 278288 254898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 47568 237454 47888 237486
rect 47568 237218 47610 237454
rect 47846 237218 47888 237454
rect 47568 237134 47888 237218
rect 47568 236898 47610 237134
rect 47846 236898 47888 237134
rect 47568 236866 47888 236898
rect 78288 237454 78608 237486
rect 78288 237218 78330 237454
rect 78566 237218 78608 237454
rect 78288 237134 78608 237218
rect 78288 236898 78330 237134
rect 78566 236898 78608 237134
rect 78288 236866 78608 236898
rect 109008 237454 109328 237486
rect 109008 237218 109050 237454
rect 109286 237218 109328 237454
rect 109008 237134 109328 237218
rect 109008 236898 109050 237134
rect 109286 236898 109328 237134
rect 109008 236866 109328 236898
rect 139728 237454 140048 237486
rect 139728 237218 139770 237454
rect 140006 237218 140048 237454
rect 139728 237134 140048 237218
rect 139728 236898 139770 237134
rect 140006 236898 140048 237134
rect 139728 236866 140048 236898
rect 170448 237454 170768 237486
rect 170448 237218 170490 237454
rect 170726 237218 170768 237454
rect 170448 237134 170768 237218
rect 170448 236898 170490 237134
rect 170726 236898 170768 237134
rect 170448 236866 170768 236898
rect 201168 237454 201488 237486
rect 201168 237218 201210 237454
rect 201446 237218 201488 237454
rect 201168 237134 201488 237218
rect 201168 236898 201210 237134
rect 201446 236898 201488 237134
rect 201168 236866 201488 236898
rect 231888 237454 232208 237486
rect 231888 237218 231930 237454
rect 232166 237218 232208 237454
rect 231888 237134 232208 237218
rect 231888 236898 231930 237134
rect 232166 236898 232208 237134
rect 231888 236866 232208 236898
rect 262608 237454 262928 237486
rect 262608 237218 262650 237454
rect 262886 237218 262928 237454
rect 262608 237134 262928 237218
rect 262608 236898 262650 237134
rect 262886 236898 262928 237134
rect 262608 236866 262928 236898
rect 293328 237454 293648 237486
rect 293328 237218 293370 237454
rect 293606 237218 293648 237454
rect 293328 237134 293648 237218
rect 293328 236898 293370 237134
rect 293606 236898 293648 237134
rect 293328 236866 293648 236898
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 32208 219454 32528 219486
rect 32208 219218 32250 219454
rect 32486 219218 32528 219454
rect 32208 219134 32528 219218
rect 32208 218898 32250 219134
rect 32486 218898 32528 219134
rect 32208 218866 32528 218898
rect 62928 219454 63248 219486
rect 62928 219218 62970 219454
rect 63206 219218 63248 219454
rect 62928 219134 63248 219218
rect 62928 218898 62970 219134
rect 63206 218898 63248 219134
rect 62928 218866 63248 218898
rect 93648 219454 93968 219486
rect 93648 219218 93690 219454
rect 93926 219218 93968 219454
rect 93648 219134 93968 219218
rect 93648 218898 93690 219134
rect 93926 218898 93968 219134
rect 93648 218866 93968 218898
rect 124368 219454 124688 219486
rect 124368 219218 124410 219454
rect 124646 219218 124688 219454
rect 124368 219134 124688 219218
rect 124368 218898 124410 219134
rect 124646 218898 124688 219134
rect 124368 218866 124688 218898
rect 155088 219454 155408 219486
rect 155088 219218 155130 219454
rect 155366 219218 155408 219454
rect 155088 219134 155408 219218
rect 155088 218898 155130 219134
rect 155366 218898 155408 219134
rect 155088 218866 155408 218898
rect 185808 219454 186128 219486
rect 185808 219218 185850 219454
rect 186086 219218 186128 219454
rect 185808 219134 186128 219218
rect 185808 218898 185850 219134
rect 186086 218898 186128 219134
rect 185808 218866 186128 218898
rect 216528 219454 216848 219486
rect 216528 219218 216570 219454
rect 216806 219218 216848 219454
rect 216528 219134 216848 219218
rect 216528 218898 216570 219134
rect 216806 218898 216848 219134
rect 216528 218866 216848 218898
rect 247248 219454 247568 219486
rect 247248 219218 247290 219454
rect 247526 219218 247568 219454
rect 247248 219134 247568 219218
rect 247248 218898 247290 219134
rect 247526 218898 247568 219134
rect 247248 218866 247568 218898
rect 277968 219454 278288 219486
rect 277968 219218 278010 219454
rect 278246 219218 278288 219454
rect 277968 219134 278288 219218
rect 277968 218898 278010 219134
rect 278246 218898 278288 219134
rect 277968 218866 278288 218898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 47568 201454 47888 201486
rect 47568 201218 47610 201454
rect 47846 201218 47888 201454
rect 47568 201134 47888 201218
rect 47568 200898 47610 201134
rect 47846 200898 47888 201134
rect 47568 200866 47888 200898
rect 78288 201454 78608 201486
rect 78288 201218 78330 201454
rect 78566 201218 78608 201454
rect 78288 201134 78608 201218
rect 78288 200898 78330 201134
rect 78566 200898 78608 201134
rect 78288 200866 78608 200898
rect 109008 201454 109328 201486
rect 109008 201218 109050 201454
rect 109286 201218 109328 201454
rect 109008 201134 109328 201218
rect 109008 200898 109050 201134
rect 109286 200898 109328 201134
rect 109008 200866 109328 200898
rect 139728 201454 140048 201486
rect 139728 201218 139770 201454
rect 140006 201218 140048 201454
rect 139728 201134 140048 201218
rect 139728 200898 139770 201134
rect 140006 200898 140048 201134
rect 139728 200866 140048 200898
rect 170448 201454 170768 201486
rect 170448 201218 170490 201454
rect 170726 201218 170768 201454
rect 170448 201134 170768 201218
rect 170448 200898 170490 201134
rect 170726 200898 170768 201134
rect 170448 200866 170768 200898
rect 201168 201454 201488 201486
rect 201168 201218 201210 201454
rect 201446 201218 201488 201454
rect 201168 201134 201488 201218
rect 201168 200898 201210 201134
rect 201446 200898 201488 201134
rect 201168 200866 201488 200898
rect 231888 201454 232208 201486
rect 231888 201218 231930 201454
rect 232166 201218 232208 201454
rect 231888 201134 232208 201218
rect 231888 200898 231930 201134
rect 232166 200898 232208 201134
rect 231888 200866 232208 200898
rect 262608 201454 262928 201486
rect 262608 201218 262650 201454
rect 262886 201218 262928 201454
rect 262608 201134 262928 201218
rect 262608 200898 262650 201134
rect 262886 200898 262928 201134
rect 262608 200866 262928 200898
rect 293328 201454 293648 201486
rect 293328 201218 293370 201454
rect 293606 201218 293648 201454
rect 293328 201134 293648 201218
rect 293328 200898 293370 201134
rect 293606 200898 293648 201134
rect 293328 200866 293648 200898
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 32208 183454 32528 183486
rect 32208 183218 32250 183454
rect 32486 183218 32528 183454
rect 32208 183134 32528 183218
rect 32208 182898 32250 183134
rect 32486 182898 32528 183134
rect 32208 182866 32528 182898
rect 62928 183454 63248 183486
rect 62928 183218 62970 183454
rect 63206 183218 63248 183454
rect 62928 183134 63248 183218
rect 62928 182898 62970 183134
rect 63206 182898 63248 183134
rect 62928 182866 63248 182898
rect 93648 183454 93968 183486
rect 93648 183218 93690 183454
rect 93926 183218 93968 183454
rect 93648 183134 93968 183218
rect 93648 182898 93690 183134
rect 93926 182898 93968 183134
rect 93648 182866 93968 182898
rect 124368 183454 124688 183486
rect 124368 183218 124410 183454
rect 124646 183218 124688 183454
rect 124368 183134 124688 183218
rect 124368 182898 124410 183134
rect 124646 182898 124688 183134
rect 124368 182866 124688 182898
rect 155088 183454 155408 183486
rect 155088 183218 155130 183454
rect 155366 183218 155408 183454
rect 155088 183134 155408 183218
rect 155088 182898 155130 183134
rect 155366 182898 155408 183134
rect 155088 182866 155408 182898
rect 185808 183454 186128 183486
rect 185808 183218 185850 183454
rect 186086 183218 186128 183454
rect 185808 183134 186128 183218
rect 185808 182898 185850 183134
rect 186086 182898 186128 183134
rect 185808 182866 186128 182898
rect 216528 183454 216848 183486
rect 216528 183218 216570 183454
rect 216806 183218 216848 183454
rect 216528 183134 216848 183218
rect 216528 182898 216570 183134
rect 216806 182898 216848 183134
rect 216528 182866 216848 182898
rect 247248 183454 247568 183486
rect 247248 183218 247290 183454
rect 247526 183218 247568 183454
rect 247248 183134 247568 183218
rect 247248 182898 247290 183134
rect 247526 182898 247568 183134
rect 247248 182866 247568 182898
rect 277968 183454 278288 183486
rect 277968 183218 278010 183454
rect 278246 183218 278288 183454
rect 277968 183134 278288 183218
rect 277968 182898 278010 183134
rect 278246 182898 278288 183134
rect 277968 182866 278288 182898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 47568 165454 47888 165486
rect 47568 165218 47610 165454
rect 47846 165218 47888 165454
rect 47568 165134 47888 165218
rect 47568 164898 47610 165134
rect 47846 164898 47888 165134
rect 47568 164866 47888 164898
rect 78288 165454 78608 165486
rect 78288 165218 78330 165454
rect 78566 165218 78608 165454
rect 78288 165134 78608 165218
rect 78288 164898 78330 165134
rect 78566 164898 78608 165134
rect 78288 164866 78608 164898
rect 109008 165454 109328 165486
rect 109008 165218 109050 165454
rect 109286 165218 109328 165454
rect 109008 165134 109328 165218
rect 109008 164898 109050 165134
rect 109286 164898 109328 165134
rect 109008 164866 109328 164898
rect 139728 165454 140048 165486
rect 139728 165218 139770 165454
rect 140006 165218 140048 165454
rect 139728 165134 140048 165218
rect 139728 164898 139770 165134
rect 140006 164898 140048 165134
rect 139728 164866 140048 164898
rect 170448 165454 170768 165486
rect 170448 165218 170490 165454
rect 170726 165218 170768 165454
rect 170448 165134 170768 165218
rect 170448 164898 170490 165134
rect 170726 164898 170768 165134
rect 170448 164866 170768 164898
rect 201168 165454 201488 165486
rect 201168 165218 201210 165454
rect 201446 165218 201488 165454
rect 201168 165134 201488 165218
rect 201168 164898 201210 165134
rect 201446 164898 201488 165134
rect 201168 164866 201488 164898
rect 231888 165454 232208 165486
rect 231888 165218 231930 165454
rect 232166 165218 232208 165454
rect 231888 165134 232208 165218
rect 231888 164898 231930 165134
rect 232166 164898 232208 165134
rect 231888 164866 232208 164898
rect 262608 165454 262928 165486
rect 262608 165218 262650 165454
rect 262886 165218 262928 165454
rect 262608 165134 262928 165218
rect 262608 164898 262650 165134
rect 262886 164898 262928 165134
rect 262608 164866 262928 164898
rect 293328 165454 293648 165486
rect 293328 165218 293370 165454
rect 293606 165218 293648 165454
rect 293328 165134 293648 165218
rect 293328 164898 293370 165134
rect 293606 164898 293648 165134
rect 293328 164866 293648 164898
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 32208 147454 32528 147486
rect 32208 147218 32250 147454
rect 32486 147218 32528 147454
rect 32208 147134 32528 147218
rect 32208 146898 32250 147134
rect 32486 146898 32528 147134
rect 32208 146866 32528 146898
rect 62928 147454 63248 147486
rect 62928 147218 62970 147454
rect 63206 147218 63248 147454
rect 62928 147134 63248 147218
rect 62928 146898 62970 147134
rect 63206 146898 63248 147134
rect 62928 146866 63248 146898
rect 93648 147454 93968 147486
rect 93648 147218 93690 147454
rect 93926 147218 93968 147454
rect 93648 147134 93968 147218
rect 93648 146898 93690 147134
rect 93926 146898 93968 147134
rect 93648 146866 93968 146898
rect 124368 147454 124688 147486
rect 124368 147218 124410 147454
rect 124646 147218 124688 147454
rect 124368 147134 124688 147218
rect 124368 146898 124410 147134
rect 124646 146898 124688 147134
rect 124368 146866 124688 146898
rect 155088 147454 155408 147486
rect 155088 147218 155130 147454
rect 155366 147218 155408 147454
rect 155088 147134 155408 147218
rect 155088 146898 155130 147134
rect 155366 146898 155408 147134
rect 155088 146866 155408 146898
rect 185808 147454 186128 147486
rect 185808 147218 185850 147454
rect 186086 147218 186128 147454
rect 185808 147134 186128 147218
rect 185808 146898 185850 147134
rect 186086 146898 186128 147134
rect 185808 146866 186128 146898
rect 216528 147454 216848 147486
rect 216528 147218 216570 147454
rect 216806 147218 216848 147454
rect 216528 147134 216848 147218
rect 216528 146898 216570 147134
rect 216806 146898 216848 147134
rect 216528 146866 216848 146898
rect 247248 147454 247568 147486
rect 247248 147218 247290 147454
rect 247526 147218 247568 147454
rect 247248 147134 247568 147218
rect 247248 146898 247290 147134
rect 247526 146898 247568 147134
rect 247248 146866 247568 146898
rect 277968 147454 278288 147486
rect 277968 147218 278010 147454
rect 278246 147218 278288 147454
rect 277968 147134 278288 147218
rect 277968 146898 278010 147134
rect 278246 146898 278288 147134
rect 277968 146866 278288 146898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 47568 129454 47888 129486
rect 47568 129218 47610 129454
rect 47846 129218 47888 129454
rect 47568 129134 47888 129218
rect 47568 128898 47610 129134
rect 47846 128898 47888 129134
rect 47568 128866 47888 128898
rect 78288 129454 78608 129486
rect 78288 129218 78330 129454
rect 78566 129218 78608 129454
rect 78288 129134 78608 129218
rect 78288 128898 78330 129134
rect 78566 128898 78608 129134
rect 78288 128866 78608 128898
rect 109008 129454 109328 129486
rect 109008 129218 109050 129454
rect 109286 129218 109328 129454
rect 109008 129134 109328 129218
rect 109008 128898 109050 129134
rect 109286 128898 109328 129134
rect 109008 128866 109328 128898
rect 139728 129454 140048 129486
rect 139728 129218 139770 129454
rect 140006 129218 140048 129454
rect 139728 129134 140048 129218
rect 139728 128898 139770 129134
rect 140006 128898 140048 129134
rect 139728 128866 140048 128898
rect 170448 129454 170768 129486
rect 170448 129218 170490 129454
rect 170726 129218 170768 129454
rect 170448 129134 170768 129218
rect 170448 128898 170490 129134
rect 170726 128898 170768 129134
rect 170448 128866 170768 128898
rect 201168 129454 201488 129486
rect 201168 129218 201210 129454
rect 201446 129218 201488 129454
rect 201168 129134 201488 129218
rect 201168 128898 201210 129134
rect 201446 128898 201488 129134
rect 201168 128866 201488 128898
rect 231888 129454 232208 129486
rect 231888 129218 231930 129454
rect 232166 129218 232208 129454
rect 231888 129134 232208 129218
rect 231888 128898 231930 129134
rect 232166 128898 232208 129134
rect 231888 128866 232208 128898
rect 262608 129454 262928 129486
rect 262608 129218 262650 129454
rect 262886 129218 262928 129454
rect 262608 129134 262928 129218
rect 262608 128898 262650 129134
rect 262886 128898 262928 129134
rect 262608 128866 262928 128898
rect 293328 129454 293648 129486
rect 293328 129218 293370 129454
rect 293606 129218 293648 129454
rect 293328 129134 293648 129218
rect 293328 128898 293370 129134
rect 293606 128898 293648 129134
rect 293328 128866 293648 128898
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 32208 111454 32528 111486
rect 32208 111218 32250 111454
rect 32486 111218 32528 111454
rect 32208 111134 32528 111218
rect 32208 110898 32250 111134
rect 32486 110898 32528 111134
rect 32208 110866 32528 110898
rect 62928 111454 63248 111486
rect 62928 111218 62970 111454
rect 63206 111218 63248 111454
rect 62928 111134 63248 111218
rect 62928 110898 62970 111134
rect 63206 110898 63248 111134
rect 62928 110866 63248 110898
rect 93648 111454 93968 111486
rect 93648 111218 93690 111454
rect 93926 111218 93968 111454
rect 93648 111134 93968 111218
rect 93648 110898 93690 111134
rect 93926 110898 93968 111134
rect 93648 110866 93968 110898
rect 124368 111454 124688 111486
rect 124368 111218 124410 111454
rect 124646 111218 124688 111454
rect 124368 111134 124688 111218
rect 124368 110898 124410 111134
rect 124646 110898 124688 111134
rect 124368 110866 124688 110898
rect 155088 111454 155408 111486
rect 155088 111218 155130 111454
rect 155366 111218 155408 111454
rect 155088 111134 155408 111218
rect 155088 110898 155130 111134
rect 155366 110898 155408 111134
rect 155088 110866 155408 110898
rect 185808 111454 186128 111486
rect 185808 111218 185850 111454
rect 186086 111218 186128 111454
rect 185808 111134 186128 111218
rect 185808 110898 185850 111134
rect 186086 110898 186128 111134
rect 185808 110866 186128 110898
rect 216528 111454 216848 111486
rect 216528 111218 216570 111454
rect 216806 111218 216848 111454
rect 216528 111134 216848 111218
rect 216528 110898 216570 111134
rect 216806 110898 216848 111134
rect 216528 110866 216848 110898
rect 247248 111454 247568 111486
rect 247248 111218 247290 111454
rect 247526 111218 247568 111454
rect 247248 111134 247568 111218
rect 247248 110898 247290 111134
rect 247526 110898 247568 111134
rect 247248 110866 247568 110898
rect 277968 111454 278288 111486
rect 277968 111218 278010 111454
rect 278246 111218 278288 111454
rect 277968 111134 278288 111218
rect 277968 110898 278010 111134
rect 278246 110898 278288 111134
rect 277968 110866 278288 110898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 47568 93454 47888 93486
rect 47568 93218 47610 93454
rect 47846 93218 47888 93454
rect 47568 93134 47888 93218
rect 47568 92898 47610 93134
rect 47846 92898 47888 93134
rect 47568 92866 47888 92898
rect 78288 93454 78608 93486
rect 78288 93218 78330 93454
rect 78566 93218 78608 93454
rect 78288 93134 78608 93218
rect 78288 92898 78330 93134
rect 78566 92898 78608 93134
rect 78288 92866 78608 92898
rect 109008 93454 109328 93486
rect 109008 93218 109050 93454
rect 109286 93218 109328 93454
rect 109008 93134 109328 93218
rect 109008 92898 109050 93134
rect 109286 92898 109328 93134
rect 109008 92866 109328 92898
rect 139728 93454 140048 93486
rect 139728 93218 139770 93454
rect 140006 93218 140048 93454
rect 139728 93134 140048 93218
rect 139728 92898 139770 93134
rect 140006 92898 140048 93134
rect 139728 92866 140048 92898
rect 170448 93454 170768 93486
rect 170448 93218 170490 93454
rect 170726 93218 170768 93454
rect 170448 93134 170768 93218
rect 170448 92898 170490 93134
rect 170726 92898 170768 93134
rect 170448 92866 170768 92898
rect 201168 93454 201488 93486
rect 201168 93218 201210 93454
rect 201446 93218 201488 93454
rect 201168 93134 201488 93218
rect 201168 92898 201210 93134
rect 201446 92898 201488 93134
rect 201168 92866 201488 92898
rect 231888 93454 232208 93486
rect 231888 93218 231930 93454
rect 232166 93218 232208 93454
rect 231888 93134 232208 93218
rect 231888 92898 231930 93134
rect 232166 92898 232208 93134
rect 231888 92866 232208 92898
rect 262608 93454 262928 93486
rect 262608 93218 262650 93454
rect 262886 93218 262928 93454
rect 262608 93134 262928 93218
rect 262608 92898 262650 93134
rect 262886 92898 262928 93134
rect 262608 92866 262928 92898
rect 293328 93454 293648 93486
rect 293328 93218 293370 93454
rect 293606 93218 293648 93454
rect 293328 93134 293648 93218
rect 293328 92898 293370 93134
rect 293606 92898 293648 93134
rect 293328 92866 293648 92898
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 32208 75454 32528 75486
rect 32208 75218 32250 75454
rect 32486 75218 32528 75454
rect 32208 75134 32528 75218
rect 32208 74898 32250 75134
rect 32486 74898 32528 75134
rect 32208 74866 32528 74898
rect 62928 75454 63248 75486
rect 62928 75218 62970 75454
rect 63206 75218 63248 75454
rect 62928 75134 63248 75218
rect 62928 74898 62970 75134
rect 63206 74898 63248 75134
rect 62928 74866 63248 74898
rect 93648 75454 93968 75486
rect 93648 75218 93690 75454
rect 93926 75218 93968 75454
rect 93648 75134 93968 75218
rect 93648 74898 93690 75134
rect 93926 74898 93968 75134
rect 93648 74866 93968 74898
rect 124368 75454 124688 75486
rect 124368 75218 124410 75454
rect 124646 75218 124688 75454
rect 124368 75134 124688 75218
rect 124368 74898 124410 75134
rect 124646 74898 124688 75134
rect 124368 74866 124688 74898
rect 155088 75454 155408 75486
rect 155088 75218 155130 75454
rect 155366 75218 155408 75454
rect 155088 75134 155408 75218
rect 155088 74898 155130 75134
rect 155366 74898 155408 75134
rect 155088 74866 155408 74898
rect 185808 75454 186128 75486
rect 185808 75218 185850 75454
rect 186086 75218 186128 75454
rect 185808 75134 186128 75218
rect 185808 74898 185850 75134
rect 186086 74898 186128 75134
rect 185808 74866 186128 74898
rect 216528 75454 216848 75486
rect 216528 75218 216570 75454
rect 216806 75218 216848 75454
rect 216528 75134 216848 75218
rect 216528 74898 216570 75134
rect 216806 74898 216848 75134
rect 216528 74866 216848 74898
rect 247248 75454 247568 75486
rect 247248 75218 247290 75454
rect 247526 75218 247568 75454
rect 247248 75134 247568 75218
rect 247248 74898 247290 75134
rect 247526 74898 247568 75134
rect 247248 74866 247568 74898
rect 277968 75454 278288 75486
rect 277968 75218 278010 75454
rect 278246 75218 278288 75454
rect 277968 75134 278288 75218
rect 277968 74898 278010 75134
rect 278246 74898 278288 75134
rect 277968 74866 278288 74898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 47568 57454 47888 57486
rect 47568 57218 47610 57454
rect 47846 57218 47888 57454
rect 47568 57134 47888 57218
rect 47568 56898 47610 57134
rect 47846 56898 47888 57134
rect 47568 56866 47888 56898
rect 78288 57454 78608 57486
rect 78288 57218 78330 57454
rect 78566 57218 78608 57454
rect 78288 57134 78608 57218
rect 78288 56898 78330 57134
rect 78566 56898 78608 57134
rect 78288 56866 78608 56898
rect 109008 57454 109328 57486
rect 109008 57218 109050 57454
rect 109286 57218 109328 57454
rect 109008 57134 109328 57218
rect 109008 56898 109050 57134
rect 109286 56898 109328 57134
rect 109008 56866 109328 56898
rect 139728 57454 140048 57486
rect 139728 57218 139770 57454
rect 140006 57218 140048 57454
rect 139728 57134 140048 57218
rect 139728 56898 139770 57134
rect 140006 56898 140048 57134
rect 139728 56866 140048 56898
rect 170448 57454 170768 57486
rect 170448 57218 170490 57454
rect 170726 57218 170768 57454
rect 170448 57134 170768 57218
rect 170448 56898 170490 57134
rect 170726 56898 170768 57134
rect 170448 56866 170768 56898
rect 201168 57454 201488 57486
rect 201168 57218 201210 57454
rect 201446 57218 201488 57454
rect 201168 57134 201488 57218
rect 201168 56898 201210 57134
rect 201446 56898 201488 57134
rect 201168 56866 201488 56898
rect 231888 57454 232208 57486
rect 231888 57218 231930 57454
rect 232166 57218 232208 57454
rect 231888 57134 232208 57218
rect 231888 56898 231930 57134
rect 232166 56898 232208 57134
rect 231888 56866 232208 56898
rect 262608 57454 262928 57486
rect 262608 57218 262650 57454
rect 262886 57218 262928 57454
rect 262608 57134 262928 57218
rect 262608 56898 262650 57134
rect 262886 56898 262928 57134
rect 262608 56866 262928 56898
rect 293328 57454 293648 57486
rect 293328 57218 293370 57454
rect 293606 57218 293648 57454
rect 293328 57134 293648 57218
rect 293328 56898 293370 57134
rect 293606 56898 293648 57134
rect 293328 56866 293648 56898
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 32208 39454 32528 39486
rect 32208 39218 32250 39454
rect 32486 39218 32528 39454
rect 32208 39134 32528 39218
rect 32208 38898 32250 39134
rect 32486 38898 32528 39134
rect 32208 38866 32528 38898
rect 62928 39454 63248 39486
rect 62928 39218 62970 39454
rect 63206 39218 63248 39454
rect 62928 39134 63248 39218
rect 62928 38898 62970 39134
rect 63206 38898 63248 39134
rect 62928 38866 63248 38898
rect 93648 39454 93968 39486
rect 93648 39218 93690 39454
rect 93926 39218 93968 39454
rect 93648 39134 93968 39218
rect 93648 38898 93690 39134
rect 93926 38898 93968 39134
rect 93648 38866 93968 38898
rect 124368 39454 124688 39486
rect 124368 39218 124410 39454
rect 124646 39218 124688 39454
rect 124368 39134 124688 39218
rect 124368 38898 124410 39134
rect 124646 38898 124688 39134
rect 124368 38866 124688 38898
rect 155088 39454 155408 39486
rect 155088 39218 155130 39454
rect 155366 39218 155408 39454
rect 155088 39134 155408 39218
rect 155088 38898 155130 39134
rect 155366 38898 155408 39134
rect 155088 38866 155408 38898
rect 185808 39454 186128 39486
rect 185808 39218 185850 39454
rect 186086 39218 186128 39454
rect 185808 39134 186128 39218
rect 185808 38898 185850 39134
rect 186086 38898 186128 39134
rect 185808 38866 186128 38898
rect 216528 39454 216848 39486
rect 216528 39218 216570 39454
rect 216806 39218 216848 39454
rect 216528 39134 216848 39218
rect 216528 38898 216570 39134
rect 216806 38898 216848 39134
rect 216528 38866 216848 38898
rect 247248 39454 247568 39486
rect 247248 39218 247290 39454
rect 247526 39218 247568 39454
rect 247248 39134 247568 39218
rect 247248 38898 247290 39134
rect 247526 38898 247568 39134
rect 247248 38866 247568 38898
rect 277968 39454 278288 39486
rect 277968 39218 278010 39454
rect 278246 39218 278288 39454
rect 277968 39134 278288 39218
rect 277968 38898 278010 39134
rect 278246 38898 278288 39134
rect 277968 38866 278288 38898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 37794 3454 38414 32000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 55794 21454 56414 32000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 73794 3454 74414 32000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 91794 21454 92414 32000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 109794 3454 110414 32000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 127794 21454 128414 32000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 145794 3454 146414 32000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 163794 21454 164414 32000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 181794 3454 182414 32000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 199794 21454 200414 32000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 217794 3454 218414 32000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 235794 21454 236414 32000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 253794 3454 254414 32000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 271794 21454 272414 32000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 289794 3454 290414 32000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 701262 398414 704282
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 701262 416414 705242
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 701262 434414 704282
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 701262 452414 705242
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 701262 470414 704282
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 701262 488414 705242
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 701262 506414 704282
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 701262 524414 705242
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 701262 542414 704282
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 701262 560414 705242
rect 577794 704838 578414 705830
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 394766 687454 398024 687486
rect 394766 687218 394837 687454
rect 395073 687218 395157 687454
rect 395393 687218 395477 687454
rect 395713 687218 395797 687454
rect 396033 687218 396117 687454
rect 396353 687218 396437 687454
rect 396673 687218 396757 687454
rect 396993 687218 397077 687454
rect 397313 687218 397397 687454
rect 397633 687218 397717 687454
rect 397953 687218 398024 687454
rect 394766 687134 398024 687218
rect 394766 686898 394837 687134
rect 395073 686898 395157 687134
rect 395393 686898 395477 687134
rect 395713 686898 395797 687134
rect 396033 686898 396117 687134
rect 396353 686898 396437 687134
rect 396673 686898 396757 687134
rect 396993 686898 397077 687134
rect 397313 686898 397397 687134
rect 397633 686898 397717 687134
rect 397953 686898 398024 687134
rect 394766 686866 398024 686898
rect 461456 687454 462396 687486
rect 461456 687218 461488 687454
rect 461724 687218 461808 687454
rect 462044 687218 462128 687454
rect 462364 687218 462396 687454
rect 461456 687134 462396 687218
rect 461456 686898 461488 687134
rect 461724 686898 461808 687134
rect 462044 686898 462128 687134
rect 462364 686898 462396 687134
rect 461456 686866 462396 686898
rect 538132 687454 546798 687486
rect 538132 687218 538187 687454
rect 538423 687218 538507 687454
rect 538743 687218 538827 687454
rect 539063 687218 539147 687454
rect 539383 687218 539467 687454
rect 539703 687218 539787 687454
rect 540023 687218 540107 687454
rect 540343 687218 540427 687454
rect 540663 687218 540747 687454
rect 540983 687218 541067 687454
rect 541303 687218 541387 687454
rect 541623 687218 541707 687454
rect 541943 687218 542027 687454
rect 542263 687218 542347 687454
rect 542583 687218 542667 687454
rect 542903 687218 542987 687454
rect 543223 687218 543307 687454
rect 543543 687218 543627 687454
rect 543863 687218 543947 687454
rect 544183 687218 544267 687454
rect 544503 687218 544587 687454
rect 544823 687218 544907 687454
rect 545143 687218 545227 687454
rect 545463 687218 545547 687454
rect 545783 687218 545867 687454
rect 546103 687218 546187 687454
rect 546423 687218 546507 687454
rect 546743 687218 546798 687454
rect 538132 687134 546798 687218
rect 538132 686898 538187 687134
rect 538423 686898 538507 687134
rect 538743 686898 538827 687134
rect 539063 686898 539147 687134
rect 539383 686898 539467 687134
rect 539703 686898 539787 687134
rect 540023 686898 540107 687134
rect 540343 686898 540427 687134
rect 540663 686898 540747 687134
rect 540983 686898 541067 687134
rect 541303 686898 541387 687134
rect 541623 686898 541707 687134
rect 541943 686898 542027 687134
rect 542263 686898 542347 687134
rect 542583 686898 542667 687134
rect 542903 686898 542987 687134
rect 543223 686898 543307 687134
rect 543543 686898 543627 687134
rect 543863 686898 543947 687134
rect 544183 686898 544267 687134
rect 544503 686898 544587 687134
rect 544823 686898 544907 687134
rect 545143 686898 545227 687134
rect 545463 686898 545547 687134
rect 545783 686898 545867 687134
rect 546103 686898 546187 687134
rect 546423 686898 546507 687134
rect 546743 686898 546798 687134
rect 538132 686866 546798 686898
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 399978 669454 403236 669486
rect 399978 669218 400049 669454
rect 400285 669218 400369 669454
rect 400605 669218 400689 669454
rect 400925 669218 401009 669454
rect 401245 669218 401329 669454
rect 401565 669218 401649 669454
rect 401885 669218 401969 669454
rect 402205 669218 402289 669454
rect 402525 669218 402609 669454
rect 402845 669218 402929 669454
rect 403165 669218 403236 669454
rect 399978 669134 403236 669218
rect 399978 668898 400049 669134
rect 400285 668898 400369 669134
rect 400605 668898 400689 669134
rect 400925 668898 401009 669134
rect 401245 668898 401329 669134
rect 401565 668898 401649 669134
rect 401885 668898 401969 669134
rect 402205 668898 402289 669134
rect 402525 668898 402609 669134
rect 402845 668898 402929 669134
rect 403165 668898 403236 669134
rect 399978 668866 403236 668898
rect 549206 669454 555800 669486
rect 549206 669218 549345 669454
rect 549581 669218 549665 669454
rect 549901 669218 549985 669454
rect 550221 669218 550305 669454
rect 550541 669218 550625 669454
rect 550861 669218 550945 669454
rect 551181 669218 551265 669454
rect 551501 669218 551585 669454
rect 551821 669218 551905 669454
rect 552141 669218 552225 669454
rect 552461 669218 552545 669454
rect 552781 669218 552865 669454
rect 553101 669218 553185 669454
rect 553421 669218 553505 669454
rect 553741 669218 553825 669454
rect 554061 669218 554145 669454
rect 554381 669218 554465 669454
rect 554701 669218 554785 669454
rect 555021 669218 555105 669454
rect 555341 669218 555425 669454
rect 555661 669218 555800 669454
rect 549206 669134 555800 669218
rect 549206 668898 549345 669134
rect 549581 668898 549665 669134
rect 549901 668898 549985 669134
rect 550221 668898 550305 669134
rect 550541 668898 550625 669134
rect 550861 668898 550945 669134
rect 551181 668898 551265 669134
rect 551501 668898 551585 669134
rect 551821 668898 551905 669134
rect 552141 668898 552225 669134
rect 552461 668898 552545 669134
rect 552781 668898 552865 669134
rect 553101 668898 553185 669134
rect 553421 668898 553505 669134
rect 553741 668898 553825 669134
rect 554061 668898 554145 669134
rect 554381 668898 554465 669134
rect 554701 668898 554785 669134
rect 555021 668898 555105 669134
rect 555341 668898 555425 669134
rect 555661 668898 555800 669134
rect 549206 668866 555800 668898
rect 394766 651454 398024 651486
rect 394766 651218 394837 651454
rect 395073 651218 395157 651454
rect 395393 651218 395477 651454
rect 395713 651218 395797 651454
rect 396033 651218 396117 651454
rect 396353 651218 396437 651454
rect 396673 651218 396757 651454
rect 396993 651218 397077 651454
rect 397313 651218 397397 651454
rect 397633 651218 397717 651454
rect 397953 651218 398024 651454
rect 394766 651134 398024 651218
rect 394766 650898 394837 651134
rect 395073 650898 395157 651134
rect 395393 650898 395477 651134
rect 395713 650898 395797 651134
rect 396033 650898 396117 651134
rect 396353 650898 396437 651134
rect 396673 650898 396757 651134
rect 396993 650898 397077 651134
rect 397313 650898 397397 651134
rect 397633 650898 397717 651134
rect 397953 650898 398024 651134
rect 394766 650866 398024 650898
rect 459760 651454 460720 651486
rect 459760 651218 459802 651454
rect 460038 651218 460122 651454
rect 460358 651218 460442 651454
rect 460678 651218 460720 651454
rect 459760 651134 460720 651218
rect 459760 650898 459802 651134
rect 460038 650898 460122 651134
rect 460358 650898 460442 651134
rect 460678 650898 460720 651134
rect 459760 650866 460720 650898
rect 538132 651454 546798 651486
rect 538132 651218 538187 651454
rect 538423 651218 538507 651454
rect 538743 651218 538827 651454
rect 539063 651218 539147 651454
rect 539383 651218 539467 651454
rect 539703 651218 539787 651454
rect 540023 651218 540107 651454
rect 540343 651218 540427 651454
rect 540663 651218 540747 651454
rect 540983 651218 541067 651454
rect 541303 651218 541387 651454
rect 541623 651218 541707 651454
rect 541943 651218 542027 651454
rect 542263 651218 542347 651454
rect 542583 651218 542667 651454
rect 542903 651218 542987 651454
rect 543223 651218 543307 651454
rect 543543 651218 543627 651454
rect 543863 651218 543947 651454
rect 544183 651218 544267 651454
rect 544503 651218 544587 651454
rect 544823 651218 544907 651454
rect 545143 651218 545227 651454
rect 545463 651218 545547 651454
rect 545783 651218 545867 651454
rect 546103 651218 546187 651454
rect 546423 651218 546507 651454
rect 546743 651218 546798 651454
rect 538132 651134 546798 651218
rect 538132 650898 538187 651134
rect 538423 650898 538507 651134
rect 538743 650898 538827 651134
rect 539063 650898 539147 651134
rect 539383 650898 539467 651134
rect 539703 650898 539787 651134
rect 540023 650898 540107 651134
rect 540343 650898 540427 651134
rect 540663 650898 540747 651134
rect 540983 650898 541067 651134
rect 541303 650898 541387 651134
rect 541623 650898 541707 651134
rect 541943 650898 542027 651134
rect 542263 650898 542347 651134
rect 542583 650898 542667 651134
rect 542903 650898 542987 651134
rect 543223 650898 543307 651134
rect 543543 650898 543627 651134
rect 543863 650898 543947 651134
rect 544183 650898 544267 651134
rect 544503 650898 544587 651134
rect 544823 650898 544907 651134
rect 545143 650898 545227 651134
rect 545463 650898 545547 651134
rect 545783 650898 545867 651134
rect 546103 650898 546187 651134
rect 546423 650898 546507 651134
rect 546743 650898 546798 651134
rect 538132 650866 546798 650898
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 399978 633454 403236 633486
rect 399978 633218 400049 633454
rect 400285 633218 400369 633454
rect 400605 633218 400689 633454
rect 400925 633218 401009 633454
rect 401245 633218 401329 633454
rect 401565 633218 401649 633454
rect 401885 633218 401969 633454
rect 402205 633218 402289 633454
rect 402525 633218 402609 633454
rect 402845 633218 402929 633454
rect 403165 633218 403236 633454
rect 399978 633134 403236 633218
rect 399978 632898 400049 633134
rect 400285 632898 400369 633134
rect 400605 632898 400689 633134
rect 400925 632898 401009 633134
rect 401245 632898 401329 633134
rect 401565 632898 401649 633134
rect 401885 632898 401969 633134
rect 402205 632898 402289 633134
rect 402525 632898 402609 633134
rect 402845 632898 402929 633134
rect 403165 632898 403236 633134
rect 399978 632866 403236 632898
rect 424725 633454 424961 633486
rect 424725 633134 424961 633218
rect 424725 632866 424961 632898
rect 427394 633454 427630 633486
rect 427394 633134 427630 633218
rect 427394 632866 427630 632898
rect 430063 633454 430299 633486
rect 430063 633134 430299 633218
rect 430063 632866 430299 632898
rect 436728 633454 437336 633486
rect 436728 633218 436754 633454
rect 436990 633218 437074 633454
rect 437310 633218 437336 633454
rect 436728 633134 437336 633218
rect 436728 632898 436754 633134
rect 436990 632898 437074 633134
rect 437310 632898 437336 633134
rect 436728 632866 437336 632898
rect 549206 633454 555800 633486
rect 549206 633218 549345 633454
rect 549581 633218 549665 633454
rect 549901 633218 549985 633454
rect 550221 633218 550305 633454
rect 550541 633218 550625 633454
rect 550861 633218 550945 633454
rect 551181 633218 551265 633454
rect 551501 633218 551585 633454
rect 551821 633218 551905 633454
rect 552141 633218 552225 633454
rect 552461 633218 552545 633454
rect 552781 633218 552865 633454
rect 553101 633218 553185 633454
rect 553421 633218 553505 633454
rect 553741 633218 553825 633454
rect 554061 633218 554145 633454
rect 554381 633218 554465 633454
rect 554701 633218 554785 633454
rect 555021 633218 555105 633454
rect 555341 633218 555425 633454
rect 555661 633218 555800 633454
rect 549206 633134 555800 633218
rect 549206 632898 549345 633134
rect 549581 632898 549665 633134
rect 549901 632898 549985 633134
rect 550221 632898 550305 633134
rect 550541 632898 550625 633134
rect 550861 632898 550945 633134
rect 551181 632898 551265 633134
rect 551501 632898 551585 633134
rect 551821 632898 551905 633134
rect 552141 632898 552225 633134
rect 552461 632898 552545 633134
rect 552781 632898 552865 633134
rect 553101 632898 553185 633134
rect 553421 632898 553505 633134
rect 553741 632898 553825 633134
rect 554061 632898 554145 633134
rect 554381 632898 554465 633134
rect 554701 632898 554785 633134
rect 555021 632898 555105 633134
rect 555341 632898 555425 633134
rect 555661 632898 555800 633134
rect 549206 632866 555800 632898
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 397794 579454 398414 609200
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 569600 398414 578898
rect 415794 597454 416414 609200
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 569600 416414 596898
rect 433794 579454 434414 609200
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 404874 561454 405194 561486
rect 404874 561218 404916 561454
rect 405152 561218 405194 561454
rect 404874 561134 405194 561218
rect 404874 560898 404916 561134
rect 405152 560898 405194 561134
rect 404874 560866 405194 560898
rect 414805 561454 415125 561486
rect 414805 561218 414847 561454
rect 415083 561218 415125 561454
rect 414805 561134 415125 561218
rect 414805 560898 414847 561134
rect 415083 560898 415125 561134
rect 414805 560866 415125 560898
rect 399909 543454 400229 543486
rect 399909 543218 399951 543454
rect 400187 543218 400229 543454
rect 399909 543134 400229 543218
rect 399909 542898 399951 543134
rect 400187 542898 400229 543134
rect 399909 542866 400229 542898
rect 409839 543454 410159 543486
rect 409839 543218 409881 543454
rect 410117 543218 410159 543454
rect 409839 543134 410159 543218
rect 409839 542898 409881 543134
rect 410117 542898 410159 543134
rect 409839 542866 410159 542898
rect 419770 543454 420090 543486
rect 419770 543218 419812 543454
rect 420048 543218 420090 543454
rect 419770 543134 420090 543218
rect 419770 542898 419812 543134
rect 420048 542898 420090 543134
rect 419770 542866 420090 542898
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 397794 507454 398414 533600
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 415794 525454 416414 533600
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 451794 597454 452414 609200
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 469794 579454 470414 609200
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 487794 597454 488414 609200
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 505794 579454 506414 609200
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 523794 597454 524414 609200
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 541794 579454 542414 609200
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 559794 597454 560414 609200
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
<< via4 >>
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 53643 669218 53879 669454
rect 53963 669218 54199 669454
rect 54283 669218 54519 669454
rect 54603 669218 54839 669454
rect 54923 669218 55159 669454
rect 55243 669218 55479 669454
rect 53643 668898 53879 669134
rect 53963 668898 54199 669134
rect 54283 668898 54519 669134
rect 54603 668898 54839 669134
rect 54923 668898 55159 669134
rect 55243 668898 55479 669134
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 36959 633218 37195 633454
rect 37279 633218 37515 633454
rect 37599 633218 37835 633454
rect 37919 633218 38155 633454
rect 38239 633218 38475 633454
rect 38559 633218 38795 633454
rect 38879 633218 39115 633454
rect 39199 633218 39435 633454
rect 39519 633218 39755 633454
rect 39839 633218 40075 633454
rect 40159 633218 40395 633454
rect 40479 633218 40715 633454
rect 40799 633218 41035 633454
rect 41119 633218 41355 633454
rect 41439 633218 41675 633454
rect 41759 633218 41995 633454
rect 42079 633218 42315 633454
rect 42399 633218 42635 633454
rect 42719 633218 42955 633454
rect 43039 633218 43275 633454
rect 43359 633218 43595 633454
rect 43679 633218 43915 633454
rect 43999 633218 44235 633454
rect 36959 632898 37195 633134
rect 37279 632898 37515 633134
rect 37599 632898 37835 633134
rect 37919 632898 38155 633134
rect 38239 632898 38475 633134
rect 38559 632898 38795 633134
rect 38879 632898 39115 633134
rect 39199 632898 39435 633134
rect 39519 632898 39755 633134
rect 39839 632898 40075 633134
rect 40159 632898 40395 633134
rect 40479 632898 40715 633134
rect 40799 632898 41035 633134
rect 41119 632898 41355 633134
rect 41439 632898 41675 633134
rect 41759 632898 41995 633134
rect 42079 632898 42315 633134
rect 42399 632898 42635 633134
rect 42719 632898 42955 633134
rect 43039 632898 43275 633134
rect 43359 632898 43595 633134
rect 43679 632898 43915 633134
rect 43999 632898 44235 633134
rect 261535 633218 261771 633454
rect 261855 633218 262091 633454
rect 262175 633218 262411 633454
rect 262495 633218 262731 633454
rect 262815 633218 263051 633454
rect 263135 633218 263371 633454
rect 263455 633218 263691 633454
rect 263775 633218 264011 633454
rect 264095 633218 264331 633454
rect 264415 633218 264651 633454
rect 264735 633218 264971 633454
rect 265055 633218 265291 633454
rect 265375 633218 265611 633454
rect 265695 633218 265931 633454
rect 266015 633218 266251 633454
rect 266335 633218 266571 633454
rect 266655 633218 266891 633454
rect 261535 632898 261771 633134
rect 261855 632898 262091 633134
rect 262175 632898 262411 633134
rect 262495 632898 262731 633134
rect 262815 632898 263051 633134
rect 263135 632898 263371 633134
rect 263455 632898 263691 633134
rect 263775 632898 264011 633134
rect 264095 632898 264331 633134
rect 264415 632898 264651 633134
rect 264735 632898 264971 633134
rect 265055 632898 265291 633134
rect 265375 632898 265611 633134
rect 265695 632898 265931 633134
rect 266015 632898 266251 633134
rect 266335 632898 266571 633134
rect 266655 632898 266891 633134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 47470 615218 47706 615454
rect 47790 615218 48026 615454
rect 48110 615218 48346 615454
rect 48430 615218 48666 615454
rect 48750 615218 48986 615454
rect 49070 615218 49306 615454
rect 49390 615218 49626 615454
rect 49710 615218 49946 615454
rect 50030 615218 50266 615454
rect 50350 615218 50586 615454
rect 50670 615218 50906 615454
rect 50990 615218 51226 615454
rect 51310 615218 51546 615454
rect 51630 615218 51866 615454
rect 51950 615218 52186 615454
rect 52270 615218 52506 615454
rect 52590 615218 52826 615454
rect 52910 615218 53146 615454
rect 47470 614898 47706 615134
rect 47790 614898 48026 615134
rect 48110 614898 48346 615134
rect 48430 614898 48666 615134
rect 48750 614898 48986 615134
rect 49070 614898 49306 615134
rect 49390 614898 49626 615134
rect 49710 614898 49946 615134
rect 50030 614898 50266 615134
rect 50350 614898 50586 615134
rect 50670 614898 50906 615134
rect 50990 614898 51226 615134
rect 51310 614898 51546 615134
rect 51630 614898 51866 615134
rect 51950 614898 52186 615134
rect 52270 614898 52506 615134
rect 52590 614898 52826 615134
rect 52910 614898 53146 615134
rect 253323 615218 253559 615454
rect 253643 615218 253879 615454
rect 253963 615218 254199 615454
rect 254283 615218 254519 615454
rect 254603 615218 254839 615454
rect 254923 615218 255159 615454
rect 255243 615218 255479 615454
rect 255563 615218 255799 615454
rect 255883 615218 256119 615454
rect 256203 615218 256439 615454
rect 256523 615218 256759 615454
rect 256843 615218 257079 615454
rect 257163 615218 257399 615454
rect 257483 615218 257719 615454
rect 257803 615218 258039 615454
rect 253323 614898 253559 615134
rect 253643 614898 253879 615134
rect 253963 614898 254199 615134
rect 254283 614898 254519 615134
rect 254603 614898 254839 615134
rect 254923 614898 255159 615134
rect 255243 614898 255479 615134
rect 255563 614898 255799 615134
rect 255883 614898 256119 615134
rect 256203 614898 256439 615134
rect 256523 614898 256759 615134
rect 256843 614898 257079 615134
rect 257163 614898 257399 615134
rect 257483 614898 257719 615134
rect 257803 614898 258039 615134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 36959 597218 37195 597454
rect 37279 597218 37515 597454
rect 37599 597218 37835 597454
rect 37919 597218 38155 597454
rect 38239 597218 38475 597454
rect 38559 597218 38795 597454
rect 38879 597218 39115 597454
rect 39199 597218 39435 597454
rect 39519 597218 39755 597454
rect 39839 597218 40075 597454
rect 40159 597218 40395 597454
rect 40479 597218 40715 597454
rect 40799 597218 41035 597454
rect 41119 597218 41355 597454
rect 41439 597218 41675 597454
rect 41759 597218 41995 597454
rect 42079 597218 42315 597454
rect 42399 597218 42635 597454
rect 42719 597218 42955 597454
rect 43039 597218 43275 597454
rect 43359 597218 43595 597454
rect 43679 597218 43915 597454
rect 43999 597218 44235 597454
rect 36959 596898 37195 597134
rect 37279 596898 37515 597134
rect 37599 596898 37835 597134
rect 37919 596898 38155 597134
rect 38239 596898 38475 597134
rect 38559 596898 38795 597134
rect 38879 596898 39115 597134
rect 39199 596898 39435 597134
rect 39519 596898 39755 597134
rect 39839 596898 40075 597134
rect 40159 596898 40395 597134
rect 40479 596898 40715 597134
rect 40799 596898 41035 597134
rect 41119 596898 41355 597134
rect 41439 596898 41675 597134
rect 41759 596898 41995 597134
rect 42079 596898 42315 597134
rect 42399 596898 42635 597134
rect 42719 596898 42955 597134
rect 43039 596898 43275 597134
rect 43359 596898 43595 597134
rect 43679 596898 43915 597134
rect 43999 596898 44235 597134
rect 167626 597218 167862 597454
rect 167626 596898 167862 597134
rect 171918 597218 172154 597454
rect 171918 596898 172154 597134
rect 176210 597218 176446 597454
rect 176210 596898 176446 597134
rect 180502 597218 180738 597454
rect 180502 596898 180738 597134
rect 184794 597218 185030 597454
rect 184794 596898 185030 597134
rect 189366 597218 189602 597454
rect 189366 596898 189602 597134
rect 193658 597218 193894 597454
rect 193658 596898 193894 597134
rect 197950 597218 198186 597454
rect 197950 596898 198186 597134
rect 202242 597218 202478 597454
rect 202242 596898 202478 597134
rect 206534 597218 206770 597454
rect 206534 596898 206770 597134
rect 211138 597218 211374 597454
rect 211138 596898 211374 597134
rect 215430 597218 215666 597454
rect 215430 596898 215666 597134
rect 219722 597218 219958 597454
rect 219722 596898 219958 597134
rect 224014 597218 224250 597454
rect 224014 596898 224250 597134
rect 228306 597218 228542 597454
rect 228306 596898 228542 597134
rect 232826 597218 233062 597454
rect 232826 596898 233062 597134
rect 237118 597218 237354 597454
rect 237118 596898 237354 597134
rect 241410 597218 241646 597454
rect 241410 596898 241646 597134
rect 245702 597218 245938 597454
rect 245702 596898 245938 597134
rect 249994 597218 250230 597454
rect 249994 596898 250230 597134
rect 261535 597218 261771 597454
rect 261855 597218 262091 597454
rect 262175 597218 262411 597454
rect 262495 597218 262731 597454
rect 262815 597218 263051 597454
rect 263135 597218 263371 597454
rect 263455 597218 263691 597454
rect 263775 597218 264011 597454
rect 264095 597218 264331 597454
rect 264415 597218 264651 597454
rect 264735 597218 264971 597454
rect 265055 597218 265291 597454
rect 265375 597218 265611 597454
rect 265695 597218 265931 597454
rect 266015 597218 266251 597454
rect 266335 597218 266571 597454
rect 266655 597218 266891 597454
rect 261535 596898 261771 597134
rect 261855 596898 262091 597134
rect 262175 596898 262411 597134
rect 262495 596898 262731 597134
rect 262815 596898 263051 597134
rect 263135 596898 263371 597134
rect 263455 596898 263691 597134
rect 263775 596898 264011 597134
rect 264095 596898 264331 597134
rect 264415 596898 264651 597134
rect 264735 596898 264971 597134
rect 265055 596898 265291 597134
rect 265375 596898 265611 597134
rect 265695 596898 265931 597134
rect 266015 596898 266251 597134
rect 266335 596898 266571 597134
rect 266655 596898 266891 597134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 47470 579218 47706 579454
rect 47790 579218 48026 579454
rect 48110 579218 48346 579454
rect 48430 579218 48666 579454
rect 48750 579218 48986 579454
rect 49070 579218 49306 579454
rect 49390 579218 49626 579454
rect 49710 579218 49946 579454
rect 50030 579218 50266 579454
rect 50350 579218 50586 579454
rect 50670 579218 50906 579454
rect 50990 579218 51226 579454
rect 51310 579218 51546 579454
rect 51630 579218 51866 579454
rect 51950 579218 52186 579454
rect 52270 579218 52506 579454
rect 52590 579218 52826 579454
rect 52910 579218 53146 579454
rect 47470 578898 47706 579134
rect 47790 578898 48026 579134
rect 48110 578898 48346 579134
rect 48430 578898 48666 579134
rect 48750 578898 48986 579134
rect 49070 578898 49306 579134
rect 49390 578898 49626 579134
rect 49710 578898 49946 579134
rect 50030 578898 50266 579134
rect 50350 578898 50586 579134
rect 50670 578898 50906 579134
rect 50990 578898 51226 579134
rect 51310 578898 51546 579134
rect 51630 578898 51866 579134
rect 51950 578898 52186 579134
rect 52270 578898 52506 579134
rect 52590 578898 52826 579134
rect 52910 578898 53146 579134
rect 253323 579218 253559 579454
rect 253643 579218 253879 579454
rect 253963 579218 254199 579454
rect 254283 579218 254519 579454
rect 254603 579218 254839 579454
rect 254923 579218 255159 579454
rect 255243 579218 255479 579454
rect 255563 579218 255799 579454
rect 255883 579218 256119 579454
rect 256203 579218 256439 579454
rect 256523 579218 256759 579454
rect 256843 579218 257079 579454
rect 257163 579218 257399 579454
rect 257483 579218 257719 579454
rect 257803 579218 258039 579454
rect 253323 578898 253559 579134
rect 253643 578898 253879 579134
rect 253963 578898 254199 579134
rect 254283 578898 254519 579134
rect 254603 578898 254839 579134
rect 254923 578898 255159 579134
rect 255243 578898 255479 579134
rect 255563 578898 255799 579134
rect 255883 578898 256119 579134
rect 256203 578898 256439 579134
rect 256523 578898 256759 579134
rect 256843 578898 257079 579134
rect 257163 578898 257399 579134
rect 257483 578898 257719 579134
rect 257803 578898 258039 579134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 32250 291218 32486 291454
rect 32250 290898 32486 291134
rect 62970 291218 63206 291454
rect 62970 290898 63206 291134
rect 93690 291218 93926 291454
rect 93690 290898 93926 291134
rect 124410 291218 124646 291454
rect 124410 290898 124646 291134
rect 155130 291218 155366 291454
rect 155130 290898 155366 291134
rect 185850 291218 186086 291454
rect 185850 290898 186086 291134
rect 216570 291218 216806 291454
rect 216570 290898 216806 291134
rect 247290 291218 247526 291454
rect 247290 290898 247526 291134
rect 278010 291218 278246 291454
rect 278010 290898 278246 291134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 47610 273218 47846 273454
rect 47610 272898 47846 273134
rect 78330 273218 78566 273454
rect 78330 272898 78566 273134
rect 109050 273218 109286 273454
rect 109050 272898 109286 273134
rect 139770 273218 140006 273454
rect 139770 272898 140006 273134
rect 170490 273218 170726 273454
rect 170490 272898 170726 273134
rect 201210 273218 201446 273454
rect 201210 272898 201446 273134
rect 231930 273218 232166 273454
rect 231930 272898 232166 273134
rect 262650 273218 262886 273454
rect 262650 272898 262886 273134
rect 293370 273218 293606 273454
rect 293370 272898 293606 273134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 32250 255218 32486 255454
rect 32250 254898 32486 255134
rect 62970 255218 63206 255454
rect 62970 254898 63206 255134
rect 93690 255218 93926 255454
rect 93690 254898 93926 255134
rect 124410 255218 124646 255454
rect 124410 254898 124646 255134
rect 155130 255218 155366 255454
rect 155130 254898 155366 255134
rect 185850 255218 186086 255454
rect 185850 254898 186086 255134
rect 216570 255218 216806 255454
rect 216570 254898 216806 255134
rect 247290 255218 247526 255454
rect 247290 254898 247526 255134
rect 278010 255218 278246 255454
rect 278010 254898 278246 255134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 47610 237218 47846 237454
rect 47610 236898 47846 237134
rect 78330 237218 78566 237454
rect 78330 236898 78566 237134
rect 109050 237218 109286 237454
rect 109050 236898 109286 237134
rect 139770 237218 140006 237454
rect 139770 236898 140006 237134
rect 170490 237218 170726 237454
rect 170490 236898 170726 237134
rect 201210 237218 201446 237454
rect 201210 236898 201446 237134
rect 231930 237218 232166 237454
rect 231930 236898 232166 237134
rect 262650 237218 262886 237454
rect 262650 236898 262886 237134
rect 293370 237218 293606 237454
rect 293370 236898 293606 237134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 32250 219218 32486 219454
rect 32250 218898 32486 219134
rect 62970 219218 63206 219454
rect 62970 218898 63206 219134
rect 93690 219218 93926 219454
rect 93690 218898 93926 219134
rect 124410 219218 124646 219454
rect 124410 218898 124646 219134
rect 155130 219218 155366 219454
rect 155130 218898 155366 219134
rect 185850 219218 186086 219454
rect 185850 218898 186086 219134
rect 216570 219218 216806 219454
rect 216570 218898 216806 219134
rect 247290 219218 247526 219454
rect 247290 218898 247526 219134
rect 278010 219218 278246 219454
rect 278010 218898 278246 219134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 47610 201218 47846 201454
rect 47610 200898 47846 201134
rect 78330 201218 78566 201454
rect 78330 200898 78566 201134
rect 109050 201218 109286 201454
rect 109050 200898 109286 201134
rect 139770 201218 140006 201454
rect 139770 200898 140006 201134
rect 170490 201218 170726 201454
rect 170490 200898 170726 201134
rect 201210 201218 201446 201454
rect 201210 200898 201446 201134
rect 231930 201218 232166 201454
rect 231930 200898 232166 201134
rect 262650 201218 262886 201454
rect 262650 200898 262886 201134
rect 293370 201218 293606 201454
rect 293370 200898 293606 201134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 32250 183218 32486 183454
rect 32250 182898 32486 183134
rect 62970 183218 63206 183454
rect 62970 182898 63206 183134
rect 93690 183218 93926 183454
rect 93690 182898 93926 183134
rect 124410 183218 124646 183454
rect 124410 182898 124646 183134
rect 155130 183218 155366 183454
rect 155130 182898 155366 183134
rect 185850 183218 186086 183454
rect 185850 182898 186086 183134
rect 216570 183218 216806 183454
rect 216570 182898 216806 183134
rect 247290 183218 247526 183454
rect 247290 182898 247526 183134
rect 278010 183218 278246 183454
rect 278010 182898 278246 183134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 47610 165218 47846 165454
rect 47610 164898 47846 165134
rect 78330 165218 78566 165454
rect 78330 164898 78566 165134
rect 109050 165218 109286 165454
rect 109050 164898 109286 165134
rect 139770 165218 140006 165454
rect 139770 164898 140006 165134
rect 170490 165218 170726 165454
rect 170490 164898 170726 165134
rect 201210 165218 201446 165454
rect 201210 164898 201446 165134
rect 231930 165218 232166 165454
rect 231930 164898 232166 165134
rect 262650 165218 262886 165454
rect 262650 164898 262886 165134
rect 293370 165218 293606 165454
rect 293370 164898 293606 165134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 32250 147218 32486 147454
rect 32250 146898 32486 147134
rect 62970 147218 63206 147454
rect 62970 146898 63206 147134
rect 93690 147218 93926 147454
rect 93690 146898 93926 147134
rect 124410 147218 124646 147454
rect 124410 146898 124646 147134
rect 155130 147218 155366 147454
rect 155130 146898 155366 147134
rect 185850 147218 186086 147454
rect 185850 146898 186086 147134
rect 216570 147218 216806 147454
rect 216570 146898 216806 147134
rect 247290 147218 247526 147454
rect 247290 146898 247526 147134
rect 278010 147218 278246 147454
rect 278010 146898 278246 147134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 47610 129218 47846 129454
rect 47610 128898 47846 129134
rect 78330 129218 78566 129454
rect 78330 128898 78566 129134
rect 109050 129218 109286 129454
rect 109050 128898 109286 129134
rect 139770 129218 140006 129454
rect 139770 128898 140006 129134
rect 170490 129218 170726 129454
rect 170490 128898 170726 129134
rect 201210 129218 201446 129454
rect 201210 128898 201446 129134
rect 231930 129218 232166 129454
rect 231930 128898 232166 129134
rect 262650 129218 262886 129454
rect 262650 128898 262886 129134
rect 293370 129218 293606 129454
rect 293370 128898 293606 129134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 32250 111218 32486 111454
rect 32250 110898 32486 111134
rect 62970 111218 63206 111454
rect 62970 110898 63206 111134
rect 93690 111218 93926 111454
rect 93690 110898 93926 111134
rect 124410 111218 124646 111454
rect 124410 110898 124646 111134
rect 155130 111218 155366 111454
rect 155130 110898 155366 111134
rect 185850 111218 186086 111454
rect 185850 110898 186086 111134
rect 216570 111218 216806 111454
rect 216570 110898 216806 111134
rect 247290 111218 247526 111454
rect 247290 110898 247526 111134
rect 278010 111218 278246 111454
rect 278010 110898 278246 111134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 47610 93218 47846 93454
rect 47610 92898 47846 93134
rect 78330 93218 78566 93454
rect 78330 92898 78566 93134
rect 109050 93218 109286 93454
rect 109050 92898 109286 93134
rect 139770 93218 140006 93454
rect 139770 92898 140006 93134
rect 170490 93218 170726 93454
rect 170490 92898 170726 93134
rect 201210 93218 201446 93454
rect 201210 92898 201446 93134
rect 231930 93218 232166 93454
rect 231930 92898 232166 93134
rect 262650 93218 262886 93454
rect 262650 92898 262886 93134
rect 293370 93218 293606 93454
rect 293370 92898 293606 93134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 32250 75218 32486 75454
rect 32250 74898 32486 75134
rect 62970 75218 63206 75454
rect 62970 74898 63206 75134
rect 93690 75218 93926 75454
rect 93690 74898 93926 75134
rect 124410 75218 124646 75454
rect 124410 74898 124646 75134
rect 155130 75218 155366 75454
rect 155130 74898 155366 75134
rect 185850 75218 186086 75454
rect 185850 74898 186086 75134
rect 216570 75218 216806 75454
rect 216570 74898 216806 75134
rect 247290 75218 247526 75454
rect 247290 74898 247526 75134
rect 278010 75218 278246 75454
rect 278010 74898 278246 75134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 47610 57218 47846 57454
rect 47610 56898 47846 57134
rect 78330 57218 78566 57454
rect 78330 56898 78566 57134
rect 109050 57218 109286 57454
rect 109050 56898 109286 57134
rect 139770 57218 140006 57454
rect 139770 56898 140006 57134
rect 170490 57218 170726 57454
rect 170490 56898 170726 57134
rect 201210 57218 201446 57454
rect 201210 56898 201446 57134
rect 231930 57218 232166 57454
rect 231930 56898 232166 57134
rect 262650 57218 262886 57454
rect 262650 56898 262886 57134
rect 293370 57218 293606 57454
rect 293370 56898 293606 57134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 32250 39218 32486 39454
rect 32250 38898 32486 39134
rect 62970 39218 63206 39454
rect 62970 38898 63206 39134
rect 93690 39218 93926 39454
rect 93690 38898 93926 39134
rect 124410 39218 124646 39454
rect 124410 38898 124646 39134
rect 155130 39218 155366 39454
rect 155130 38898 155366 39134
rect 185850 39218 186086 39454
rect 185850 38898 186086 39134
rect 216570 39218 216806 39454
rect 216570 38898 216806 39134
rect 247290 39218 247526 39454
rect 247290 38898 247526 39134
rect 278010 39218 278246 39454
rect 278010 38898 278246 39134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 394837 687218 395073 687454
rect 395157 687218 395393 687454
rect 395477 687218 395713 687454
rect 395797 687218 396033 687454
rect 396117 687218 396353 687454
rect 396437 687218 396673 687454
rect 396757 687218 396993 687454
rect 397077 687218 397313 687454
rect 397397 687218 397633 687454
rect 397717 687218 397953 687454
rect 394837 686898 395073 687134
rect 395157 686898 395393 687134
rect 395477 686898 395713 687134
rect 395797 686898 396033 687134
rect 396117 686898 396353 687134
rect 396437 686898 396673 687134
rect 396757 686898 396993 687134
rect 397077 686898 397313 687134
rect 397397 686898 397633 687134
rect 397717 686898 397953 687134
rect 461488 687218 461724 687454
rect 461808 687218 462044 687454
rect 462128 687218 462364 687454
rect 461488 686898 461724 687134
rect 461808 686898 462044 687134
rect 462128 686898 462364 687134
rect 538187 687218 538423 687454
rect 538507 687218 538743 687454
rect 538827 687218 539063 687454
rect 539147 687218 539383 687454
rect 539467 687218 539703 687454
rect 539787 687218 540023 687454
rect 540107 687218 540343 687454
rect 540427 687218 540663 687454
rect 540747 687218 540983 687454
rect 541067 687218 541303 687454
rect 541387 687218 541623 687454
rect 541707 687218 541943 687454
rect 542027 687218 542263 687454
rect 542347 687218 542583 687454
rect 542667 687218 542903 687454
rect 542987 687218 543223 687454
rect 543307 687218 543543 687454
rect 543627 687218 543863 687454
rect 543947 687218 544183 687454
rect 544267 687218 544503 687454
rect 544587 687218 544823 687454
rect 544907 687218 545143 687454
rect 545227 687218 545463 687454
rect 545547 687218 545783 687454
rect 545867 687218 546103 687454
rect 546187 687218 546423 687454
rect 546507 687218 546743 687454
rect 538187 686898 538423 687134
rect 538507 686898 538743 687134
rect 538827 686898 539063 687134
rect 539147 686898 539383 687134
rect 539467 686898 539703 687134
rect 539787 686898 540023 687134
rect 540107 686898 540343 687134
rect 540427 686898 540663 687134
rect 540747 686898 540983 687134
rect 541067 686898 541303 687134
rect 541387 686898 541623 687134
rect 541707 686898 541943 687134
rect 542027 686898 542263 687134
rect 542347 686898 542583 687134
rect 542667 686898 542903 687134
rect 542987 686898 543223 687134
rect 543307 686898 543543 687134
rect 543627 686898 543863 687134
rect 543947 686898 544183 687134
rect 544267 686898 544503 687134
rect 544587 686898 544823 687134
rect 544907 686898 545143 687134
rect 545227 686898 545463 687134
rect 545547 686898 545783 687134
rect 545867 686898 546103 687134
rect 546187 686898 546423 687134
rect 546507 686898 546743 687134
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 400049 669218 400285 669454
rect 400369 669218 400605 669454
rect 400689 669218 400925 669454
rect 401009 669218 401245 669454
rect 401329 669218 401565 669454
rect 401649 669218 401885 669454
rect 401969 669218 402205 669454
rect 402289 669218 402525 669454
rect 402609 669218 402845 669454
rect 402929 669218 403165 669454
rect 400049 668898 400285 669134
rect 400369 668898 400605 669134
rect 400689 668898 400925 669134
rect 401009 668898 401245 669134
rect 401329 668898 401565 669134
rect 401649 668898 401885 669134
rect 401969 668898 402205 669134
rect 402289 668898 402525 669134
rect 402609 668898 402845 669134
rect 402929 668898 403165 669134
rect 549345 669218 549581 669454
rect 549665 669218 549901 669454
rect 549985 669218 550221 669454
rect 550305 669218 550541 669454
rect 550625 669218 550861 669454
rect 550945 669218 551181 669454
rect 551265 669218 551501 669454
rect 551585 669218 551821 669454
rect 551905 669218 552141 669454
rect 552225 669218 552461 669454
rect 552545 669218 552781 669454
rect 552865 669218 553101 669454
rect 553185 669218 553421 669454
rect 553505 669218 553741 669454
rect 553825 669218 554061 669454
rect 554145 669218 554381 669454
rect 554465 669218 554701 669454
rect 554785 669218 555021 669454
rect 555105 669218 555341 669454
rect 555425 669218 555661 669454
rect 549345 668898 549581 669134
rect 549665 668898 549901 669134
rect 549985 668898 550221 669134
rect 550305 668898 550541 669134
rect 550625 668898 550861 669134
rect 550945 668898 551181 669134
rect 551265 668898 551501 669134
rect 551585 668898 551821 669134
rect 551905 668898 552141 669134
rect 552225 668898 552461 669134
rect 552545 668898 552781 669134
rect 552865 668898 553101 669134
rect 553185 668898 553421 669134
rect 553505 668898 553741 669134
rect 553825 668898 554061 669134
rect 554145 668898 554381 669134
rect 554465 668898 554701 669134
rect 554785 668898 555021 669134
rect 555105 668898 555341 669134
rect 555425 668898 555661 669134
rect 394837 651218 395073 651454
rect 395157 651218 395393 651454
rect 395477 651218 395713 651454
rect 395797 651218 396033 651454
rect 396117 651218 396353 651454
rect 396437 651218 396673 651454
rect 396757 651218 396993 651454
rect 397077 651218 397313 651454
rect 397397 651218 397633 651454
rect 397717 651218 397953 651454
rect 394837 650898 395073 651134
rect 395157 650898 395393 651134
rect 395477 650898 395713 651134
rect 395797 650898 396033 651134
rect 396117 650898 396353 651134
rect 396437 650898 396673 651134
rect 396757 650898 396993 651134
rect 397077 650898 397313 651134
rect 397397 650898 397633 651134
rect 397717 650898 397953 651134
rect 459802 651218 460038 651454
rect 460122 651218 460358 651454
rect 460442 651218 460678 651454
rect 459802 650898 460038 651134
rect 460122 650898 460358 651134
rect 460442 650898 460678 651134
rect 538187 651218 538423 651454
rect 538507 651218 538743 651454
rect 538827 651218 539063 651454
rect 539147 651218 539383 651454
rect 539467 651218 539703 651454
rect 539787 651218 540023 651454
rect 540107 651218 540343 651454
rect 540427 651218 540663 651454
rect 540747 651218 540983 651454
rect 541067 651218 541303 651454
rect 541387 651218 541623 651454
rect 541707 651218 541943 651454
rect 542027 651218 542263 651454
rect 542347 651218 542583 651454
rect 542667 651218 542903 651454
rect 542987 651218 543223 651454
rect 543307 651218 543543 651454
rect 543627 651218 543863 651454
rect 543947 651218 544183 651454
rect 544267 651218 544503 651454
rect 544587 651218 544823 651454
rect 544907 651218 545143 651454
rect 545227 651218 545463 651454
rect 545547 651218 545783 651454
rect 545867 651218 546103 651454
rect 546187 651218 546423 651454
rect 546507 651218 546743 651454
rect 538187 650898 538423 651134
rect 538507 650898 538743 651134
rect 538827 650898 539063 651134
rect 539147 650898 539383 651134
rect 539467 650898 539703 651134
rect 539787 650898 540023 651134
rect 540107 650898 540343 651134
rect 540427 650898 540663 651134
rect 540747 650898 540983 651134
rect 541067 650898 541303 651134
rect 541387 650898 541623 651134
rect 541707 650898 541943 651134
rect 542027 650898 542263 651134
rect 542347 650898 542583 651134
rect 542667 650898 542903 651134
rect 542987 650898 543223 651134
rect 543307 650898 543543 651134
rect 543627 650898 543863 651134
rect 543947 650898 544183 651134
rect 544267 650898 544503 651134
rect 544587 650898 544823 651134
rect 544907 650898 545143 651134
rect 545227 650898 545463 651134
rect 545547 650898 545783 651134
rect 545867 650898 546103 651134
rect 546187 650898 546423 651134
rect 546507 650898 546743 651134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 400049 633218 400285 633454
rect 400369 633218 400605 633454
rect 400689 633218 400925 633454
rect 401009 633218 401245 633454
rect 401329 633218 401565 633454
rect 401649 633218 401885 633454
rect 401969 633218 402205 633454
rect 402289 633218 402525 633454
rect 402609 633218 402845 633454
rect 402929 633218 403165 633454
rect 400049 632898 400285 633134
rect 400369 632898 400605 633134
rect 400689 632898 400925 633134
rect 401009 632898 401245 633134
rect 401329 632898 401565 633134
rect 401649 632898 401885 633134
rect 401969 632898 402205 633134
rect 402289 632898 402525 633134
rect 402609 632898 402845 633134
rect 402929 632898 403165 633134
rect 424725 633218 424961 633454
rect 424725 632898 424961 633134
rect 427394 633218 427630 633454
rect 427394 632898 427630 633134
rect 430063 633218 430299 633454
rect 430063 632898 430299 633134
rect 436754 633218 436990 633454
rect 437074 633218 437310 633454
rect 436754 632898 436990 633134
rect 437074 632898 437310 633134
rect 549345 633218 549581 633454
rect 549665 633218 549901 633454
rect 549985 633218 550221 633454
rect 550305 633218 550541 633454
rect 550625 633218 550861 633454
rect 550945 633218 551181 633454
rect 551265 633218 551501 633454
rect 551585 633218 551821 633454
rect 551905 633218 552141 633454
rect 552225 633218 552461 633454
rect 552545 633218 552781 633454
rect 552865 633218 553101 633454
rect 553185 633218 553421 633454
rect 553505 633218 553741 633454
rect 553825 633218 554061 633454
rect 554145 633218 554381 633454
rect 554465 633218 554701 633454
rect 554785 633218 555021 633454
rect 555105 633218 555341 633454
rect 555425 633218 555661 633454
rect 549345 632898 549581 633134
rect 549665 632898 549901 633134
rect 549985 632898 550221 633134
rect 550305 632898 550541 633134
rect 550625 632898 550861 633134
rect 550945 632898 551181 633134
rect 551265 632898 551501 633134
rect 551585 632898 551821 633134
rect 551905 632898 552141 633134
rect 552225 632898 552461 633134
rect 552545 632898 552781 633134
rect 552865 632898 553101 633134
rect 553185 632898 553421 633134
rect 553505 632898 553741 633134
rect 553825 632898 554061 633134
rect 554145 632898 554381 633134
rect 554465 632898 554701 633134
rect 554785 632898 555021 633134
rect 555105 632898 555341 633134
rect 555425 632898 555661 633134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 404916 561218 405152 561454
rect 404916 560898 405152 561134
rect 414847 561218 415083 561454
rect 414847 560898 415083 561134
rect 399951 543218 400187 543454
rect 399951 542898 400187 543134
rect 409881 543218 410117 543454
rect 409881 542898 410117 543134
rect 419812 543218 420048 543454
rect 419812 542898 420048 543134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
<< metal5 >>
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 394837 687454
rect 395073 687218 395157 687454
rect 395393 687218 395477 687454
rect 395713 687218 395797 687454
rect 396033 687218 396117 687454
rect 396353 687218 396437 687454
rect 396673 687218 396757 687454
rect 396993 687218 397077 687454
rect 397313 687218 397397 687454
rect 397633 687218 397717 687454
rect 397953 687218 461488 687454
rect 461724 687218 461808 687454
rect 462044 687218 462128 687454
rect 462364 687218 538187 687454
rect 538423 687218 538507 687454
rect 538743 687218 538827 687454
rect 539063 687218 539147 687454
rect 539383 687218 539467 687454
rect 539703 687218 539787 687454
rect 540023 687218 540107 687454
rect 540343 687218 540427 687454
rect 540663 687218 540747 687454
rect 540983 687218 541067 687454
rect 541303 687218 541387 687454
rect 541623 687218 541707 687454
rect 541943 687218 542027 687454
rect 542263 687218 542347 687454
rect 542583 687218 542667 687454
rect 542903 687218 542987 687454
rect 543223 687218 543307 687454
rect 543543 687218 543627 687454
rect 543863 687218 543947 687454
rect 544183 687218 544267 687454
rect 544503 687218 544587 687454
rect 544823 687218 544907 687454
rect 545143 687218 545227 687454
rect 545463 687218 545547 687454
rect 545783 687218 545867 687454
rect 546103 687218 546187 687454
rect 546423 687218 546507 687454
rect 546743 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 394837 687134
rect 395073 686898 395157 687134
rect 395393 686898 395477 687134
rect 395713 686898 395797 687134
rect 396033 686898 396117 687134
rect 396353 686898 396437 687134
rect 396673 686898 396757 687134
rect 396993 686898 397077 687134
rect 397313 686898 397397 687134
rect 397633 686898 397717 687134
rect 397953 686898 461488 687134
rect 461724 686898 461808 687134
rect 462044 686898 462128 687134
rect 462364 686898 538187 687134
rect 538423 686898 538507 687134
rect 538743 686898 538827 687134
rect 539063 686898 539147 687134
rect 539383 686898 539467 687134
rect 539703 686898 539787 687134
rect 540023 686898 540107 687134
rect 540343 686898 540427 687134
rect 540663 686898 540747 687134
rect 540983 686898 541067 687134
rect 541303 686898 541387 687134
rect 541623 686898 541707 687134
rect 541943 686898 542027 687134
rect 542263 686898 542347 687134
rect 542583 686898 542667 687134
rect 542903 686898 542987 687134
rect 543223 686898 543307 687134
rect 543543 686898 543627 687134
rect 543863 686898 543947 687134
rect 544183 686898 544267 687134
rect 544503 686898 544587 687134
rect 544823 686898 544907 687134
rect 545143 686898 545227 687134
rect 545463 686898 545547 687134
rect 545783 686898 545867 687134
rect 546103 686898 546187 687134
rect 546423 686898 546507 687134
rect 546743 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 53643 669454
rect 53879 669218 53963 669454
rect 54199 669218 54283 669454
rect 54519 669218 54603 669454
rect 54839 669218 54923 669454
rect 55159 669218 55243 669454
rect 55479 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 400049 669454
rect 400285 669218 400369 669454
rect 400605 669218 400689 669454
rect 400925 669218 401009 669454
rect 401245 669218 401329 669454
rect 401565 669218 401649 669454
rect 401885 669218 401969 669454
rect 402205 669218 402289 669454
rect 402525 669218 402609 669454
rect 402845 669218 402929 669454
rect 403165 669218 549345 669454
rect 549581 669218 549665 669454
rect 549901 669218 549985 669454
rect 550221 669218 550305 669454
rect 550541 669218 550625 669454
rect 550861 669218 550945 669454
rect 551181 669218 551265 669454
rect 551501 669218 551585 669454
rect 551821 669218 551905 669454
rect 552141 669218 552225 669454
rect 552461 669218 552545 669454
rect 552781 669218 552865 669454
rect 553101 669218 553185 669454
rect 553421 669218 553505 669454
rect 553741 669218 553825 669454
rect 554061 669218 554145 669454
rect 554381 669218 554465 669454
rect 554701 669218 554785 669454
rect 555021 669218 555105 669454
rect 555341 669218 555425 669454
rect 555661 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 53643 669134
rect 53879 668898 53963 669134
rect 54199 668898 54283 669134
rect 54519 668898 54603 669134
rect 54839 668898 54923 669134
rect 55159 668898 55243 669134
rect 55479 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 400049 669134
rect 400285 668898 400369 669134
rect 400605 668898 400689 669134
rect 400925 668898 401009 669134
rect 401245 668898 401329 669134
rect 401565 668898 401649 669134
rect 401885 668898 401969 669134
rect 402205 668898 402289 669134
rect 402525 668898 402609 669134
rect 402845 668898 402929 669134
rect 403165 668898 549345 669134
rect 549581 668898 549665 669134
rect 549901 668898 549985 669134
rect 550221 668898 550305 669134
rect 550541 668898 550625 669134
rect 550861 668898 550945 669134
rect 551181 668898 551265 669134
rect 551501 668898 551585 669134
rect 551821 668898 551905 669134
rect 552141 668898 552225 669134
rect 552461 668898 552545 669134
rect 552781 668898 552865 669134
rect 553101 668898 553185 669134
rect 553421 668898 553505 669134
rect 553741 668898 553825 669134
rect 554061 668898 554145 669134
rect 554381 668898 554465 669134
rect 554701 668898 554785 669134
rect 555021 668898 555105 669134
rect 555341 668898 555425 669134
rect 555661 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 394837 651454
rect 395073 651218 395157 651454
rect 395393 651218 395477 651454
rect 395713 651218 395797 651454
rect 396033 651218 396117 651454
rect 396353 651218 396437 651454
rect 396673 651218 396757 651454
rect 396993 651218 397077 651454
rect 397313 651218 397397 651454
rect 397633 651218 397717 651454
rect 397953 651218 459802 651454
rect 460038 651218 460122 651454
rect 460358 651218 460442 651454
rect 460678 651218 538187 651454
rect 538423 651218 538507 651454
rect 538743 651218 538827 651454
rect 539063 651218 539147 651454
rect 539383 651218 539467 651454
rect 539703 651218 539787 651454
rect 540023 651218 540107 651454
rect 540343 651218 540427 651454
rect 540663 651218 540747 651454
rect 540983 651218 541067 651454
rect 541303 651218 541387 651454
rect 541623 651218 541707 651454
rect 541943 651218 542027 651454
rect 542263 651218 542347 651454
rect 542583 651218 542667 651454
rect 542903 651218 542987 651454
rect 543223 651218 543307 651454
rect 543543 651218 543627 651454
rect 543863 651218 543947 651454
rect 544183 651218 544267 651454
rect 544503 651218 544587 651454
rect 544823 651218 544907 651454
rect 545143 651218 545227 651454
rect 545463 651218 545547 651454
rect 545783 651218 545867 651454
rect 546103 651218 546187 651454
rect 546423 651218 546507 651454
rect 546743 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 394837 651134
rect 395073 650898 395157 651134
rect 395393 650898 395477 651134
rect 395713 650898 395797 651134
rect 396033 650898 396117 651134
rect 396353 650898 396437 651134
rect 396673 650898 396757 651134
rect 396993 650898 397077 651134
rect 397313 650898 397397 651134
rect 397633 650898 397717 651134
rect 397953 650898 459802 651134
rect 460038 650898 460122 651134
rect 460358 650898 460442 651134
rect 460678 650898 538187 651134
rect 538423 650898 538507 651134
rect 538743 650898 538827 651134
rect 539063 650898 539147 651134
rect 539383 650898 539467 651134
rect 539703 650898 539787 651134
rect 540023 650898 540107 651134
rect 540343 650898 540427 651134
rect 540663 650898 540747 651134
rect 540983 650898 541067 651134
rect 541303 650898 541387 651134
rect 541623 650898 541707 651134
rect 541943 650898 542027 651134
rect 542263 650898 542347 651134
rect 542583 650898 542667 651134
rect 542903 650898 542987 651134
rect 543223 650898 543307 651134
rect 543543 650898 543627 651134
rect 543863 650898 543947 651134
rect 544183 650898 544267 651134
rect 544503 650898 544587 651134
rect 544823 650898 544907 651134
rect 545143 650898 545227 651134
rect 545463 650898 545547 651134
rect 545783 650898 545867 651134
rect 546103 650898 546187 651134
rect 546423 650898 546507 651134
rect 546743 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 36959 633454
rect 37195 633218 37279 633454
rect 37515 633218 37599 633454
rect 37835 633218 37919 633454
rect 38155 633218 38239 633454
rect 38475 633218 38559 633454
rect 38795 633218 38879 633454
rect 39115 633218 39199 633454
rect 39435 633218 39519 633454
rect 39755 633218 39839 633454
rect 40075 633218 40159 633454
rect 40395 633218 40479 633454
rect 40715 633218 40799 633454
rect 41035 633218 41119 633454
rect 41355 633218 41439 633454
rect 41675 633218 41759 633454
rect 41995 633218 42079 633454
rect 42315 633218 42399 633454
rect 42635 633218 42719 633454
rect 42955 633218 43039 633454
rect 43275 633218 43359 633454
rect 43595 633218 43679 633454
rect 43915 633218 43999 633454
rect 44235 633218 261535 633454
rect 261771 633218 261855 633454
rect 262091 633218 262175 633454
rect 262411 633218 262495 633454
rect 262731 633218 262815 633454
rect 263051 633218 263135 633454
rect 263371 633218 263455 633454
rect 263691 633218 263775 633454
rect 264011 633218 264095 633454
rect 264331 633218 264415 633454
rect 264651 633218 264735 633454
rect 264971 633218 265055 633454
rect 265291 633218 265375 633454
rect 265611 633218 265695 633454
rect 265931 633218 266015 633454
rect 266251 633218 266335 633454
rect 266571 633218 266655 633454
rect 266891 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 400049 633454
rect 400285 633218 400369 633454
rect 400605 633218 400689 633454
rect 400925 633218 401009 633454
rect 401245 633218 401329 633454
rect 401565 633218 401649 633454
rect 401885 633218 401969 633454
rect 402205 633218 402289 633454
rect 402525 633218 402609 633454
rect 402845 633218 402929 633454
rect 403165 633218 424725 633454
rect 424961 633218 427394 633454
rect 427630 633218 430063 633454
rect 430299 633218 436754 633454
rect 436990 633218 437074 633454
rect 437310 633218 549345 633454
rect 549581 633218 549665 633454
rect 549901 633218 549985 633454
rect 550221 633218 550305 633454
rect 550541 633218 550625 633454
rect 550861 633218 550945 633454
rect 551181 633218 551265 633454
rect 551501 633218 551585 633454
rect 551821 633218 551905 633454
rect 552141 633218 552225 633454
rect 552461 633218 552545 633454
rect 552781 633218 552865 633454
rect 553101 633218 553185 633454
rect 553421 633218 553505 633454
rect 553741 633218 553825 633454
rect 554061 633218 554145 633454
rect 554381 633218 554465 633454
rect 554701 633218 554785 633454
rect 555021 633218 555105 633454
rect 555341 633218 555425 633454
rect 555661 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 36959 633134
rect 37195 632898 37279 633134
rect 37515 632898 37599 633134
rect 37835 632898 37919 633134
rect 38155 632898 38239 633134
rect 38475 632898 38559 633134
rect 38795 632898 38879 633134
rect 39115 632898 39199 633134
rect 39435 632898 39519 633134
rect 39755 632898 39839 633134
rect 40075 632898 40159 633134
rect 40395 632898 40479 633134
rect 40715 632898 40799 633134
rect 41035 632898 41119 633134
rect 41355 632898 41439 633134
rect 41675 632898 41759 633134
rect 41995 632898 42079 633134
rect 42315 632898 42399 633134
rect 42635 632898 42719 633134
rect 42955 632898 43039 633134
rect 43275 632898 43359 633134
rect 43595 632898 43679 633134
rect 43915 632898 43999 633134
rect 44235 632898 261535 633134
rect 261771 632898 261855 633134
rect 262091 632898 262175 633134
rect 262411 632898 262495 633134
rect 262731 632898 262815 633134
rect 263051 632898 263135 633134
rect 263371 632898 263455 633134
rect 263691 632898 263775 633134
rect 264011 632898 264095 633134
rect 264331 632898 264415 633134
rect 264651 632898 264735 633134
rect 264971 632898 265055 633134
rect 265291 632898 265375 633134
rect 265611 632898 265695 633134
rect 265931 632898 266015 633134
rect 266251 632898 266335 633134
rect 266571 632898 266655 633134
rect 266891 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 400049 633134
rect 400285 632898 400369 633134
rect 400605 632898 400689 633134
rect 400925 632898 401009 633134
rect 401245 632898 401329 633134
rect 401565 632898 401649 633134
rect 401885 632898 401969 633134
rect 402205 632898 402289 633134
rect 402525 632898 402609 633134
rect 402845 632898 402929 633134
rect 403165 632898 424725 633134
rect 424961 632898 427394 633134
rect 427630 632898 430063 633134
rect 430299 632898 436754 633134
rect 436990 632898 437074 633134
rect 437310 632898 549345 633134
rect 549581 632898 549665 633134
rect 549901 632898 549985 633134
rect 550221 632898 550305 633134
rect 550541 632898 550625 633134
rect 550861 632898 550945 633134
rect 551181 632898 551265 633134
rect 551501 632898 551585 633134
rect 551821 632898 551905 633134
rect 552141 632898 552225 633134
rect 552461 632898 552545 633134
rect 552781 632898 552865 633134
rect 553101 632898 553185 633134
rect 553421 632898 553505 633134
rect 553741 632898 553825 633134
rect 554061 632898 554145 633134
rect 554381 632898 554465 633134
rect 554701 632898 554785 633134
rect 555021 632898 555105 633134
rect 555341 632898 555425 633134
rect 555661 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 47470 615454
rect 47706 615218 47790 615454
rect 48026 615218 48110 615454
rect 48346 615218 48430 615454
rect 48666 615218 48750 615454
rect 48986 615218 49070 615454
rect 49306 615218 49390 615454
rect 49626 615218 49710 615454
rect 49946 615218 50030 615454
rect 50266 615218 50350 615454
rect 50586 615218 50670 615454
rect 50906 615218 50990 615454
rect 51226 615218 51310 615454
rect 51546 615218 51630 615454
rect 51866 615218 51950 615454
rect 52186 615218 52270 615454
rect 52506 615218 52590 615454
rect 52826 615218 52910 615454
rect 53146 615218 253323 615454
rect 253559 615218 253643 615454
rect 253879 615218 253963 615454
rect 254199 615218 254283 615454
rect 254519 615218 254603 615454
rect 254839 615218 254923 615454
rect 255159 615218 255243 615454
rect 255479 615218 255563 615454
rect 255799 615218 255883 615454
rect 256119 615218 256203 615454
rect 256439 615218 256523 615454
rect 256759 615218 256843 615454
rect 257079 615218 257163 615454
rect 257399 615218 257483 615454
rect 257719 615218 257803 615454
rect 258039 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 47470 615134
rect 47706 614898 47790 615134
rect 48026 614898 48110 615134
rect 48346 614898 48430 615134
rect 48666 614898 48750 615134
rect 48986 614898 49070 615134
rect 49306 614898 49390 615134
rect 49626 614898 49710 615134
rect 49946 614898 50030 615134
rect 50266 614898 50350 615134
rect 50586 614898 50670 615134
rect 50906 614898 50990 615134
rect 51226 614898 51310 615134
rect 51546 614898 51630 615134
rect 51866 614898 51950 615134
rect 52186 614898 52270 615134
rect 52506 614898 52590 615134
rect 52826 614898 52910 615134
rect 53146 614898 253323 615134
rect 253559 614898 253643 615134
rect 253879 614898 253963 615134
rect 254199 614898 254283 615134
rect 254519 614898 254603 615134
rect 254839 614898 254923 615134
rect 255159 614898 255243 615134
rect 255479 614898 255563 615134
rect 255799 614898 255883 615134
rect 256119 614898 256203 615134
rect 256439 614898 256523 615134
rect 256759 614898 256843 615134
rect 257079 614898 257163 615134
rect 257399 614898 257483 615134
rect 257719 614898 257803 615134
rect 258039 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 36959 597454
rect 37195 597218 37279 597454
rect 37515 597218 37599 597454
rect 37835 597218 37919 597454
rect 38155 597218 38239 597454
rect 38475 597218 38559 597454
rect 38795 597218 38879 597454
rect 39115 597218 39199 597454
rect 39435 597218 39519 597454
rect 39755 597218 39839 597454
rect 40075 597218 40159 597454
rect 40395 597218 40479 597454
rect 40715 597218 40799 597454
rect 41035 597218 41119 597454
rect 41355 597218 41439 597454
rect 41675 597218 41759 597454
rect 41995 597218 42079 597454
rect 42315 597218 42399 597454
rect 42635 597218 42719 597454
rect 42955 597218 43039 597454
rect 43275 597218 43359 597454
rect 43595 597218 43679 597454
rect 43915 597218 43999 597454
rect 44235 597218 167626 597454
rect 167862 597218 171918 597454
rect 172154 597218 176210 597454
rect 176446 597218 180502 597454
rect 180738 597218 184794 597454
rect 185030 597218 189366 597454
rect 189602 597218 193658 597454
rect 193894 597218 197950 597454
rect 198186 597218 202242 597454
rect 202478 597218 206534 597454
rect 206770 597218 211138 597454
rect 211374 597218 215430 597454
rect 215666 597218 219722 597454
rect 219958 597218 224014 597454
rect 224250 597218 228306 597454
rect 228542 597218 232826 597454
rect 233062 597218 237118 597454
rect 237354 597218 241410 597454
rect 241646 597218 245702 597454
rect 245938 597218 249994 597454
rect 250230 597218 261535 597454
rect 261771 597218 261855 597454
rect 262091 597218 262175 597454
rect 262411 597218 262495 597454
rect 262731 597218 262815 597454
rect 263051 597218 263135 597454
rect 263371 597218 263455 597454
rect 263691 597218 263775 597454
rect 264011 597218 264095 597454
rect 264331 597218 264415 597454
rect 264651 597218 264735 597454
rect 264971 597218 265055 597454
rect 265291 597218 265375 597454
rect 265611 597218 265695 597454
rect 265931 597218 266015 597454
rect 266251 597218 266335 597454
rect 266571 597218 266655 597454
rect 266891 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 36959 597134
rect 37195 596898 37279 597134
rect 37515 596898 37599 597134
rect 37835 596898 37919 597134
rect 38155 596898 38239 597134
rect 38475 596898 38559 597134
rect 38795 596898 38879 597134
rect 39115 596898 39199 597134
rect 39435 596898 39519 597134
rect 39755 596898 39839 597134
rect 40075 596898 40159 597134
rect 40395 596898 40479 597134
rect 40715 596898 40799 597134
rect 41035 596898 41119 597134
rect 41355 596898 41439 597134
rect 41675 596898 41759 597134
rect 41995 596898 42079 597134
rect 42315 596898 42399 597134
rect 42635 596898 42719 597134
rect 42955 596898 43039 597134
rect 43275 596898 43359 597134
rect 43595 596898 43679 597134
rect 43915 596898 43999 597134
rect 44235 596898 167626 597134
rect 167862 596898 171918 597134
rect 172154 596898 176210 597134
rect 176446 596898 180502 597134
rect 180738 596898 184794 597134
rect 185030 596898 189366 597134
rect 189602 596898 193658 597134
rect 193894 596898 197950 597134
rect 198186 596898 202242 597134
rect 202478 596898 206534 597134
rect 206770 596898 211138 597134
rect 211374 596898 215430 597134
rect 215666 596898 219722 597134
rect 219958 596898 224014 597134
rect 224250 596898 228306 597134
rect 228542 596898 232826 597134
rect 233062 596898 237118 597134
rect 237354 596898 241410 597134
rect 241646 596898 245702 597134
rect 245938 596898 249994 597134
rect 250230 596898 261535 597134
rect 261771 596898 261855 597134
rect 262091 596898 262175 597134
rect 262411 596898 262495 597134
rect 262731 596898 262815 597134
rect 263051 596898 263135 597134
rect 263371 596898 263455 597134
rect 263691 596898 263775 597134
rect 264011 596898 264095 597134
rect 264331 596898 264415 597134
rect 264651 596898 264735 597134
rect 264971 596898 265055 597134
rect 265291 596898 265375 597134
rect 265611 596898 265695 597134
rect 265931 596898 266015 597134
rect 266251 596898 266335 597134
rect 266571 596898 266655 597134
rect 266891 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 47470 579454
rect 47706 579218 47790 579454
rect 48026 579218 48110 579454
rect 48346 579218 48430 579454
rect 48666 579218 48750 579454
rect 48986 579218 49070 579454
rect 49306 579218 49390 579454
rect 49626 579218 49710 579454
rect 49946 579218 50030 579454
rect 50266 579218 50350 579454
rect 50586 579218 50670 579454
rect 50906 579218 50990 579454
rect 51226 579218 51310 579454
rect 51546 579218 51630 579454
rect 51866 579218 51950 579454
rect 52186 579218 52270 579454
rect 52506 579218 52590 579454
rect 52826 579218 52910 579454
rect 53146 579218 253323 579454
rect 253559 579218 253643 579454
rect 253879 579218 253963 579454
rect 254199 579218 254283 579454
rect 254519 579218 254603 579454
rect 254839 579218 254923 579454
rect 255159 579218 255243 579454
rect 255479 579218 255563 579454
rect 255799 579218 255883 579454
rect 256119 579218 256203 579454
rect 256439 579218 256523 579454
rect 256759 579218 256843 579454
rect 257079 579218 257163 579454
rect 257399 579218 257483 579454
rect 257719 579218 257803 579454
rect 258039 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 47470 579134
rect 47706 578898 47790 579134
rect 48026 578898 48110 579134
rect 48346 578898 48430 579134
rect 48666 578898 48750 579134
rect 48986 578898 49070 579134
rect 49306 578898 49390 579134
rect 49626 578898 49710 579134
rect 49946 578898 50030 579134
rect 50266 578898 50350 579134
rect 50586 578898 50670 579134
rect 50906 578898 50990 579134
rect 51226 578898 51310 579134
rect 51546 578898 51630 579134
rect 51866 578898 51950 579134
rect 52186 578898 52270 579134
rect 52506 578898 52590 579134
rect 52826 578898 52910 579134
rect 53146 578898 253323 579134
rect 253559 578898 253643 579134
rect 253879 578898 253963 579134
rect 254199 578898 254283 579134
rect 254519 578898 254603 579134
rect 254839 578898 254923 579134
rect 255159 578898 255243 579134
rect 255479 578898 255563 579134
rect 255799 578898 255883 579134
rect 256119 578898 256203 579134
rect 256439 578898 256523 579134
rect 256759 578898 256843 579134
rect 257079 578898 257163 579134
rect 257399 578898 257483 579134
rect 257719 578898 257803 579134
rect 258039 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 404916 561454
rect 405152 561218 414847 561454
rect 415083 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 404916 561134
rect 405152 560898 414847 561134
rect 415083 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 399951 543454
rect 400187 543218 409881 543454
rect 410117 543218 419812 543454
rect 420048 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 399951 543134
rect 400187 542898 409881 543134
rect 410117 542898 419812 543134
rect 420048 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 32250 291454
rect 32486 291218 62970 291454
rect 63206 291218 93690 291454
rect 93926 291218 124410 291454
rect 124646 291218 155130 291454
rect 155366 291218 185850 291454
rect 186086 291218 216570 291454
rect 216806 291218 247290 291454
rect 247526 291218 278010 291454
rect 278246 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 32250 291134
rect 32486 290898 62970 291134
rect 63206 290898 93690 291134
rect 93926 290898 124410 291134
rect 124646 290898 155130 291134
rect 155366 290898 185850 291134
rect 186086 290898 216570 291134
rect 216806 290898 247290 291134
rect 247526 290898 278010 291134
rect 278246 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 47610 273454
rect 47846 273218 78330 273454
rect 78566 273218 109050 273454
rect 109286 273218 139770 273454
rect 140006 273218 170490 273454
rect 170726 273218 201210 273454
rect 201446 273218 231930 273454
rect 232166 273218 262650 273454
rect 262886 273218 293370 273454
rect 293606 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 47610 273134
rect 47846 272898 78330 273134
rect 78566 272898 109050 273134
rect 109286 272898 139770 273134
rect 140006 272898 170490 273134
rect 170726 272898 201210 273134
rect 201446 272898 231930 273134
rect 232166 272898 262650 273134
rect 262886 272898 293370 273134
rect 293606 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 32250 255454
rect 32486 255218 62970 255454
rect 63206 255218 93690 255454
rect 93926 255218 124410 255454
rect 124646 255218 155130 255454
rect 155366 255218 185850 255454
rect 186086 255218 216570 255454
rect 216806 255218 247290 255454
rect 247526 255218 278010 255454
rect 278246 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 32250 255134
rect 32486 254898 62970 255134
rect 63206 254898 93690 255134
rect 93926 254898 124410 255134
rect 124646 254898 155130 255134
rect 155366 254898 185850 255134
rect 186086 254898 216570 255134
rect 216806 254898 247290 255134
rect 247526 254898 278010 255134
rect 278246 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 47610 237454
rect 47846 237218 78330 237454
rect 78566 237218 109050 237454
rect 109286 237218 139770 237454
rect 140006 237218 170490 237454
rect 170726 237218 201210 237454
rect 201446 237218 231930 237454
rect 232166 237218 262650 237454
rect 262886 237218 293370 237454
rect 293606 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 47610 237134
rect 47846 236898 78330 237134
rect 78566 236898 109050 237134
rect 109286 236898 139770 237134
rect 140006 236898 170490 237134
rect 170726 236898 201210 237134
rect 201446 236898 231930 237134
rect 232166 236898 262650 237134
rect 262886 236898 293370 237134
rect 293606 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 32250 219454
rect 32486 219218 62970 219454
rect 63206 219218 93690 219454
rect 93926 219218 124410 219454
rect 124646 219218 155130 219454
rect 155366 219218 185850 219454
rect 186086 219218 216570 219454
rect 216806 219218 247290 219454
rect 247526 219218 278010 219454
rect 278246 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 32250 219134
rect 32486 218898 62970 219134
rect 63206 218898 93690 219134
rect 93926 218898 124410 219134
rect 124646 218898 155130 219134
rect 155366 218898 185850 219134
rect 186086 218898 216570 219134
rect 216806 218898 247290 219134
rect 247526 218898 278010 219134
rect 278246 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 47610 201454
rect 47846 201218 78330 201454
rect 78566 201218 109050 201454
rect 109286 201218 139770 201454
rect 140006 201218 170490 201454
rect 170726 201218 201210 201454
rect 201446 201218 231930 201454
rect 232166 201218 262650 201454
rect 262886 201218 293370 201454
rect 293606 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 47610 201134
rect 47846 200898 78330 201134
rect 78566 200898 109050 201134
rect 109286 200898 139770 201134
rect 140006 200898 170490 201134
rect 170726 200898 201210 201134
rect 201446 200898 231930 201134
rect 232166 200898 262650 201134
rect 262886 200898 293370 201134
rect 293606 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 32250 183454
rect 32486 183218 62970 183454
rect 63206 183218 93690 183454
rect 93926 183218 124410 183454
rect 124646 183218 155130 183454
rect 155366 183218 185850 183454
rect 186086 183218 216570 183454
rect 216806 183218 247290 183454
rect 247526 183218 278010 183454
rect 278246 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 32250 183134
rect 32486 182898 62970 183134
rect 63206 182898 93690 183134
rect 93926 182898 124410 183134
rect 124646 182898 155130 183134
rect 155366 182898 185850 183134
rect 186086 182898 216570 183134
rect 216806 182898 247290 183134
rect 247526 182898 278010 183134
rect 278246 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 47610 165454
rect 47846 165218 78330 165454
rect 78566 165218 109050 165454
rect 109286 165218 139770 165454
rect 140006 165218 170490 165454
rect 170726 165218 201210 165454
rect 201446 165218 231930 165454
rect 232166 165218 262650 165454
rect 262886 165218 293370 165454
rect 293606 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 47610 165134
rect 47846 164898 78330 165134
rect 78566 164898 109050 165134
rect 109286 164898 139770 165134
rect 140006 164898 170490 165134
rect 170726 164898 201210 165134
rect 201446 164898 231930 165134
rect 232166 164898 262650 165134
rect 262886 164898 293370 165134
rect 293606 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 32250 147454
rect 32486 147218 62970 147454
rect 63206 147218 93690 147454
rect 93926 147218 124410 147454
rect 124646 147218 155130 147454
rect 155366 147218 185850 147454
rect 186086 147218 216570 147454
rect 216806 147218 247290 147454
rect 247526 147218 278010 147454
rect 278246 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 32250 147134
rect 32486 146898 62970 147134
rect 63206 146898 93690 147134
rect 93926 146898 124410 147134
rect 124646 146898 155130 147134
rect 155366 146898 185850 147134
rect 186086 146898 216570 147134
rect 216806 146898 247290 147134
rect 247526 146898 278010 147134
rect 278246 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 47610 129454
rect 47846 129218 78330 129454
rect 78566 129218 109050 129454
rect 109286 129218 139770 129454
rect 140006 129218 170490 129454
rect 170726 129218 201210 129454
rect 201446 129218 231930 129454
rect 232166 129218 262650 129454
rect 262886 129218 293370 129454
rect 293606 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 47610 129134
rect 47846 128898 78330 129134
rect 78566 128898 109050 129134
rect 109286 128898 139770 129134
rect 140006 128898 170490 129134
rect 170726 128898 201210 129134
rect 201446 128898 231930 129134
rect 232166 128898 262650 129134
rect 262886 128898 293370 129134
rect 293606 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 32250 111454
rect 32486 111218 62970 111454
rect 63206 111218 93690 111454
rect 93926 111218 124410 111454
rect 124646 111218 155130 111454
rect 155366 111218 185850 111454
rect 186086 111218 216570 111454
rect 216806 111218 247290 111454
rect 247526 111218 278010 111454
rect 278246 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 32250 111134
rect 32486 110898 62970 111134
rect 63206 110898 93690 111134
rect 93926 110898 124410 111134
rect 124646 110898 155130 111134
rect 155366 110898 185850 111134
rect 186086 110898 216570 111134
rect 216806 110898 247290 111134
rect 247526 110898 278010 111134
rect 278246 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 47610 93454
rect 47846 93218 78330 93454
rect 78566 93218 109050 93454
rect 109286 93218 139770 93454
rect 140006 93218 170490 93454
rect 170726 93218 201210 93454
rect 201446 93218 231930 93454
rect 232166 93218 262650 93454
rect 262886 93218 293370 93454
rect 293606 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 47610 93134
rect 47846 92898 78330 93134
rect 78566 92898 109050 93134
rect 109286 92898 139770 93134
rect 140006 92898 170490 93134
rect 170726 92898 201210 93134
rect 201446 92898 231930 93134
rect 232166 92898 262650 93134
rect 262886 92898 293370 93134
rect 293606 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 32250 75454
rect 32486 75218 62970 75454
rect 63206 75218 93690 75454
rect 93926 75218 124410 75454
rect 124646 75218 155130 75454
rect 155366 75218 185850 75454
rect 186086 75218 216570 75454
rect 216806 75218 247290 75454
rect 247526 75218 278010 75454
rect 278246 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 32250 75134
rect 32486 74898 62970 75134
rect 63206 74898 93690 75134
rect 93926 74898 124410 75134
rect 124646 74898 155130 75134
rect 155366 74898 185850 75134
rect 186086 74898 216570 75134
rect 216806 74898 247290 75134
rect 247526 74898 278010 75134
rect 278246 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 47610 57454
rect 47846 57218 78330 57454
rect 78566 57218 109050 57454
rect 109286 57218 139770 57454
rect 140006 57218 170490 57454
rect 170726 57218 201210 57454
rect 201446 57218 231930 57454
rect 232166 57218 262650 57454
rect 262886 57218 293370 57454
rect 293606 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 47610 57134
rect 47846 56898 78330 57134
rect 78566 56898 109050 57134
rect 109286 56898 139770 57134
rect 140006 56898 170490 57134
rect 170726 56898 201210 57134
rect 201446 56898 231930 57134
rect 232166 56898 262650 57134
rect 262886 56898 293370 57134
rect 293606 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 32250 39454
rect 32486 39218 62970 39454
rect 63206 39218 93690 39454
rect 93926 39218 124410 39454
rect 124646 39218 155130 39454
rect 155366 39218 185850 39454
rect 186086 39218 216570 39454
rect 216806 39218 247290 39454
rect 247526 39218 278010 39454
rect 278246 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 32250 39134
rect 32486 38898 62970 39134
rect 63206 38898 93690 39134
rect 93926 38898 124410 39134
rect 124646 38898 155130 39134
rect 155366 38898 185850 39134
rect 186086 38898 216570 39134
rect 216806 38898 247290 39134
rect 247526 38898 278010 39134
rect 278246 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
use LVDT  temp3
timestamp 1637989401
transform 1 0 58022 0 1 575250
box -26022 -21250 209012 98114
use temp_digital  temp2
timestamp 1637989401
transform 1 0 394000 0 1 535600
box 0 0 32000 32000
use analog_macro  temp1
timestamp 1637989401
transform 1 0 401554 0 1 620054
box -7554 -8854 157400 79208
use user_proj_example  mprj
timestamp 1637989401
transform 1 0 28000 0 1 34000
box 289 0 274238 276712
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 32000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 533600 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 312712 38414 552000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 312712 74414 552000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 312712 110414 552000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 312712 146414 552000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 312712 182414 552000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 312712 218414 552000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 312712 254414 552000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 569600 398414 609200 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 609200 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 609200 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 609200 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 609200 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 675364 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 675364 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 675364 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 675364 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 675364 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 675364 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 675364 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 312712 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 701262 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 701262 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 701262 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 701262 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 701262 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 55794 -1894 56414 32000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 91794 -1894 92414 32000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 127794 -1894 128414 32000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 163794 -1894 164414 32000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 199794 -1894 200414 32000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 235794 -1894 236414 32000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 271794 -1894 272414 32000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 415794 -1894 416414 533600 6 vssd1
port 532 nsew ground input
rlabel metal4 s 55794 312712 56414 552000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 91794 312712 92414 552000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 127794 312712 128414 552000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 163794 312712 164414 552000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 199794 312712 200414 552000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 235794 312712 236414 552000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 415794 569600 416414 609200 6 vssd1
port 532 nsew ground input
rlabel metal4 s 451794 -1894 452414 609200 6 vssd1
port 532 nsew ground input
rlabel metal4 s 487794 -1894 488414 609200 6 vssd1
port 532 nsew ground input
rlabel metal4 s 523794 -1894 524414 609200 6 vssd1
port 532 nsew ground input
rlabel metal4 s 559794 -1894 560414 609200 6 vssd1
port 532 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 532 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 55794 675364 56414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 91794 675364 92414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 127794 675364 128414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 163794 675364 164414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 199794 675364 200414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 235794 675364 236414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 271794 312712 272414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 415794 701262 416414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 451794 701262 452414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 487794 701262 488414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 523794 701262 524414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 559794 701262 560414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 532 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 533 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 534 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 535 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 536 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 537 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 538 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 539 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 540 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 541 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 542 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 543 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 544 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 545 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 546 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 547 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 548 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 549 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 550 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 551 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 552 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 553 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 554 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 555 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 556 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 557 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 558 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 559 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 560 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 561 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 562 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 563 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 564 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 565 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 566 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 567 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 568 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 569 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 570 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 571 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 572 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 573 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 574 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 575 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 576 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 577 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 578 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 579 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 580 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 581 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 582 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 583 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 584 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 585 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 586 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 587 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 588 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 589 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 590 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 591 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 592 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 593 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 594 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 595 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 596 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 597 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 598 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 599 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 600 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 601 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 602 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 603 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 604 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 605 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 606 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 607 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 608 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 609 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 610 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 611 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 612 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 613 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 614 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 615 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 616 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 617 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 618 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 619 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 620 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 621 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 622 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 623 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 624 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 625 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 626 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 627 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 628 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 629 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 630 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 631 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 632 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 633 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 634 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 635 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 636 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 637 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 638 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
